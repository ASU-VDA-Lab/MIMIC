module fake_ariane_3121_n_1873 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1873);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1873;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g177 ( 
.A(n_20),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_9),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_127),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_99),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_44),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_67),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_33),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_66),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_115),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_20),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_14),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_59),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_45),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_74),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_34),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_61),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_19),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_53),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_25),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_0),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_55),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_96),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_47),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_95),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_154),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_23),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_65),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_16),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_151),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_129),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_98),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_15),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_110),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_49),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_31),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_163),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_42),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_137),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_42),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_79),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_103),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_40),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_82),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_30),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_94),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_14),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_105),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_72),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_44),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_153),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_43),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_81),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_50),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_125),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_24),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_70),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_84),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_18),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_111),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_33),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_113),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_52),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_156),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_166),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_60),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_58),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_162),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_63),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_25),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_65),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_34),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_31),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_52),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_58),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_30),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_75),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_55),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_71),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_4),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_116),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_48),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_10),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_56),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_119),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_29),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_59),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_91),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_0),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_175),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_62),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_57),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_43),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_54),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_26),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_35),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_49),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_60),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_21),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_139),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_22),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_170),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_117),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_123),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_131),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_152),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_124),
.Y(n_318)
);

BUFx2_ASAP7_75t_SL g319 ( 
.A(n_77),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_120),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_63),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_1),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_122),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_87),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_106),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_27),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_12),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_145),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_40),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_28),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_126),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_53),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_10),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_147),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_101),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_157),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_24),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_108),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_69),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_11),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_57),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_28),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_136),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_12),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_9),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_56),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_107),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_90),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_143),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_118),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_304),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_185),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_272),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_2),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_178),
.B(n_3),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_186),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_329),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_213),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_188),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_245),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_211),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_201),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_225),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_301),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_258),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_344),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_329),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_349),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_285),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_190),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_181),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_201),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_192),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_193),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_187),
.B(n_3),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_285),
.B(n_4),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_229),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_236),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_187),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_196),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_178),
.B(n_5),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_196),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_197),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_199),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_288),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_248),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_268),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_203),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_290),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_197),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_198),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_198),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_206),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_206),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_210),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_210),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_308),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_228),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_326),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_228),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_234),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_250),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_191),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_234),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_237),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_250),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_305),
.B(n_5),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_237),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_201),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_288),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_250),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_205),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_209),
.B(n_7),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_238),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_212),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_311),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_214),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_218),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_238),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_221),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_281),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_334),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_239),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_239),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_334),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_256),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_230),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_202),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_256),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_240),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_371),
.B(n_434),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_362),
.Y(n_453)
);

AND2x6_ASAP7_75t_L g454 ( 
.A(n_392),
.B(n_202),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_260),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_362),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_372),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_392),
.B(n_260),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_394),
.B(n_261),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_394),
.B(n_240),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_395),
.B(n_261),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_385),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_354),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_403),
.B(n_267),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_403),
.B(n_243),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_404),
.B(n_243),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_404),
.B(n_267),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_405),
.B(n_406),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_359),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_364),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_406),
.B(n_270),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_408),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_365),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_409),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_387),
.B(n_246),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_411),
.A2(n_274),
.B(n_270),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_363),
.B(n_376),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_379),
.B(n_274),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_369),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_413),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_414),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_417),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_418),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_383),
.B(n_317),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_246),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_378),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_360),
.B(n_201),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_427),
.B(n_317),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_427),
.B(n_307),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_440),
.B(n_318),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_432),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_436),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_439),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_402),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_489),
.A2(n_387),
.B1(n_420),
.B2(n_393),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_486),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_493),
.B(n_384),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_443),
.B(n_396),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_495),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_439),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_401),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_423),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_455),
.B(n_425),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_416),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_366),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_455),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_493),
.B(n_428),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_461),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_485),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_485),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_481),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_448),
.A2(n_320),
.B(n_318),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_485),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_497),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_497),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_458),
.Y(n_546)
);

INVx4_ASAP7_75t_SL g547 ( 
.A(n_444),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_455),
.B(n_430),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_479),
.B(n_431),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_497),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_484),
.B(n_366),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_503),
.B(n_433),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_320),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_503),
.B(n_361),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_484),
.B(n_331),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_497),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_510),
.B(n_356),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_484),
.B(n_397),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_481),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_497),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_498),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_429),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_491),
.B(n_438),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_491),
.B(n_435),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_498),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_446),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_498),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_489),
.B(n_472),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_467),
.B(n_386),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_498),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_446),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_489),
.A2(n_426),
.B1(n_257),
.B2(n_259),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_470),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_467),
.B(n_353),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_467),
.B(n_217),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_498),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_489),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_498),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_459),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_331),
.Y(n_587)
);

AND3x2_ASAP7_75t_L g588 ( 
.A(n_470),
.B(n_183),
.C(n_177),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_498),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_489),
.B(n_307),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_502),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_459),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_459),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_502),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_467),
.B(n_373),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_502),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_489),
.A2(n_253),
.B1(n_343),
.B2(n_342),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_490),
.B(n_264),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_467),
.B(n_224),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_490),
.A2(n_472),
.B1(n_507),
.B2(n_464),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_506),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_447),
.B(n_415),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_463),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_447),
.B(n_419),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_480),
.B(n_249),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_505),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_463),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_480),
.B(n_352),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_505),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_488),
.B(n_339),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_505),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_339),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_505),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_492),
.B(n_377),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_490),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_492),
.B(n_179),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_505),
.Y(n_625)
);

INVx4_ASAP7_75t_SL g626 ( 
.A(n_444),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_463),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_494),
.B(n_424),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_490),
.A2(n_283),
.B1(n_282),
.B2(n_298),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_451),
.A2(n_251),
.B1(n_286),
.B2(n_284),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_494),
.B(n_180),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_463),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_475),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_505),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_513),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_513),
.Y(n_636)
);

BUFx4f_ASAP7_75t_L g637 ( 
.A(n_513),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_496),
.B(n_182),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_513),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_496),
.B(n_281),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_499),
.B(n_184),
.Y(n_642)
);

BUFx4f_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_513),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_475),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_516),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_461),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_449),
.B(n_177),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_499),
.B(n_281),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_449),
.B(n_183),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_475),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_475),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_501),
.B(n_281),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_501),
.B(n_514),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_514),
.B(n_189),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_475),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_516),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_506),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_448),
.Y(n_660)
);

NOR2x1p5_ASAP7_75t_L g661 ( 
.A(n_460),
.B(n_195),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_515),
.B(n_232),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_515),
.B(n_235),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_461),
.Y(n_666)
);

INVx11_ASAP7_75t_L g667 ( 
.A(n_444),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_461),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_516),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_517),
.B(n_456),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_584),
.A2(n_460),
.B1(n_482),
.B2(n_477),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_584),
.A2(n_462),
.B(n_477),
.C(n_468),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_538),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_559),
.B(n_516),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_660),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_526),
.B(n_456),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_602),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_608),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_525),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_590),
.A2(n_462),
.B1(n_508),
.B2(n_482),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_660),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_566),
.B(n_507),
.C(n_452),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_527),
.B(n_483),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_590),
.A2(n_572),
.B1(n_549),
.B2(n_600),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_483),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_609),
.B(n_500),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_611),
.B(n_500),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_660),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_555),
.B(n_450),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_530),
.B(n_500),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_655),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_567),
.B(n_450),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_550),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_548),
.B(n_511),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_612),
.B(n_511),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_616),
.B(n_511),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_550),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_559),
.B(n_512),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_559),
.A2(n_512),
.B1(n_472),
.B2(n_476),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_531),
.B(n_449),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_608),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_629),
.A2(n_520),
.B(n_528),
.C(n_468),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_535),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_559),
.A2(n_512),
.B1(n_472),
.B2(n_504),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_538),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_528),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_559),
.B(n_452),
.Y(n_707)
);

BUFx4_ASAP7_75t_L g708 ( 
.A(n_525),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_521),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_522),
.B(n_453),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_539),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_570),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_559),
.A2(n_490),
.B1(n_454),
.B2(n_444),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_578),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_572),
.B(n_464),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_559),
.A2(n_444),
.B1(n_454),
.B2(n_471),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_539),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_578),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_532),
.B(n_553),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_575),
.B(n_453),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_532),
.B(n_509),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_581),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_590),
.A2(n_509),
.B1(n_464),
.B2(n_504),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_535),
.B(n_457),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_572),
.B(n_476),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_546),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_546),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_601),
.A2(n_444),
.B1(n_454),
.B2(n_508),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_573),
.B(n_457),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_586),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_572),
.B(n_476),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_586),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_666),
.A2(n_469),
.B(n_465),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_661),
.B(n_465),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_661),
.B(n_469),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_555),
.B(n_473),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_592),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_580),
.B(n_473),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_SL g739 ( 
.A1(n_659),
.A2(n_410),
.B1(n_389),
.B2(n_390),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_623),
.A2(n_471),
.B(n_442),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_555),
.B(n_461),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_652),
.B(n_461),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_652),
.B(n_466),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_563),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_518),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_605),
.B(n_504),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_535),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_590),
.A2(n_509),
.B1(n_454),
.B2(n_444),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_590),
.A2(n_300),
.B1(n_271),
.B2(n_275),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_572),
.B(n_355),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_SL g751 ( 
.A(n_659),
.B(n_370),
.C(n_367),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_534),
.B(n_474),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_592),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_593),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_554),
.A2(n_302),
.B1(n_263),
.B2(n_278),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_648),
.B(n_375),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_568),
.B(n_474),
.Y(n_757)
);

BUFx5_ASAP7_75t_L g758 ( 
.A(n_652),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_541),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_533),
.B(n_466),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_579),
.A2(n_454),
.B1(n_444),
.B2(n_247),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_593),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_533),
.B(n_466),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_557),
.B(n_466),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_594),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_657),
.B(n_466),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_553),
.B(n_380),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_563),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_666),
.A2(n_474),
.B(n_466),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_601),
.A2(n_195),
.B(n_207),
.C(n_298),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_657),
.B(n_474),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_657),
.B(n_474),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_562),
.B(n_398),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_557),
.B(n_466),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_280),
.C(n_279),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_557),
.B(n_474),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_558),
.A2(n_454),
.B1(n_444),
.B2(n_216),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_618),
.A2(n_207),
.B(n_297),
.C(n_293),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_594),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_598),
.B(n_474),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_604),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_604),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_535),
.B(n_454),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_557),
.B(n_441),
.Y(n_784)
);

BUFx8_ASAP7_75t_L g785 ( 
.A(n_562),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_610),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_576),
.A2(n_454),
.B1(n_276),
.B2(n_319),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_557),
.B(n_441),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_602),
.B(n_400),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_557),
.B(n_442),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_615),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_615),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_627),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_627),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_601),
.B(n_264),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_294),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_632),
.B(n_277),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_633),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_663),
.B(n_295),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_645),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_653),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_535),
.B(n_445),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_653),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_582),
.B(n_445),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_668),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_557),
.B(n_607),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_582),
.B(n_277),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_602),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_648),
.B(n_651),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_648),
.B(n_454),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_668),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_582),
.B(n_277),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_208),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_536),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_582),
.B(n_277),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_628),
.B(n_412),
.Y(n_817)
);

O2A1O1Ixp5_ASAP7_75t_L g818 ( 
.A1(n_637),
.A2(n_662),
.B(n_643),
.C(n_591),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_602),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_582),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_624),
.A2(n_303),
.B1(n_306),
.B2(n_348),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_647),
.B(n_277),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_651),
.B(n_208),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_651),
.B(n_220),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_620),
.A2(n_283),
.B1(n_220),
.B2(n_226),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_651),
.B(n_226),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_631),
.B(n_638),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_642),
.B(n_227),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_665),
.B(n_309),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_561),
.A2(n_319),
.B1(n_350),
.B2(n_314),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_519),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_536),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_647),
.B(n_351),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_656),
.B(n_227),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_640),
.B(n_310),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_623),
.B(n_253),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_827),
.A2(n_643),
.B(n_637),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_692),
.A2(n_569),
.B(n_536),
.C(n_658),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_715),
.B(n_649),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_729),
.A2(n_643),
.B(n_637),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_796),
.A2(n_542),
.B(n_523),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_750),
.B(n_654),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_796),
.A2(n_542),
.B(n_523),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_715),
.B(n_547),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_685),
.A2(n_662),
.B(n_529),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_703),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_745),
.B(n_630),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_701),
.B(n_551),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_677),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_709),
.B(n_551),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_692),
.B(n_647),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_678),
.B(n_551),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_740),
.A2(n_529),
.B(n_519),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_670),
.B(n_552),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_797),
.A2(n_540),
.B(n_537),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_677),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_759),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_690),
.A2(n_662),
.B(n_540),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_703),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_694),
.A2(n_543),
.B(n_537),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_725),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_693),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_738),
.A2(n_544),
.B(n_543),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_810),
.A2(n_595),
.B1(n_551),
.B2(n_664),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_684),
.A2(n_591),
.B1(n_664),
.B2(n_595),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_756),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_686),
.B(n_687),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_676),
.B(n_552),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_725),
.B(n_647),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_680),
.A2(n_565),
.B1(n_595),
.B2(n_664),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_719),
.B(n_588),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_710),
.A2(n_569),
.B(n_658),
.C(n_552),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_710),
.A2(n_646),
.B(n_658),
.C(n_569),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_697),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_673),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_731),
.B(n_647),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_683),
.A2(n_545),
.B(n_544),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_721),
.B(n_255),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_767),
.B(n_255),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_756),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_785),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_679),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_773),
.B(n_266),
.Y(n_883)
);

O2A1O1Ixp5_ASAP7_75t_L g884 ( 
.A1(n_780),
.A2(n_565),
.B(n_664),
.C(n_595),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_760),
.A2(n_556),
.B(n_545),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_785),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_680),
.A2(n_266),
.B(n_282),
.C(n_291),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_712),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_672),
.A2(n_560),
.B(n_556),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_700),
.B(n_583),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_746),
.B(n_583),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_807),
.A2(n_591),
.B(n_565),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_768),
.B(n_293),
.C(n_291),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_731),
.B(n_547),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_789),
.B(n_565),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_763),
.A2(n_564),
.B(n_560),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_672),
.A2(n_571),
.B(n_564),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_706),
.B(n_591),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_733),
.A2(n_669),
.B(n_650),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_702),
.B(n_583),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_751),
.B(n_596),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_770),
.A2(n_343),
.B(n_342),
.C(n_327),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_702),
.B(n_596),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_723),
.B(n_596),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_824),
.B(n_621),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_757),
.A2(n_621),
.B(n_646),
.C(n_635),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_770),
.A2(n_327),
.B(n_330),
.C(n_599),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_809),
.B(n_819),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_758),
.B(n_621),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_826),
.B(n_671),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_695),
.B(n_635),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_703),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_689),
.A2(n_599),
.B(n_574),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_750),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_699),
.A2(n_635),
.B1(n_646),
.B2(n_636),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_736),
.A2(n_589),
.B(n_644),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_780),
.A2(n_606),
.B(n_644),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_758),
.B(n_636),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_736),
.A2(n_589),
.B(n_641),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_720),
.A2(n_585),
.B(n_641),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_744),
.B(n_587),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_696),
.B(n_636),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_714),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_708),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_757),
.A2(n_735),
.B1(n_734),
.B2(n_797),
.Y(n_925)
);

BUFx2_ASAP7_75t_SL g926 ( 
.A(n_758),
.Y(n_926)
);

AO21x1_ASAP7_75t_L g927 ( 
.A1(n_752),
.A2(n_606),
.B(n_639),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_L g928 ( 
.A1(n_752),
.A2(n_574),
.B(n_639),
.C(n_634),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_718),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_707),
.A2(n_571),
.B(n_634),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_775),
.B(n_585),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_674),
.A2(n_614),
.B(n_625),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_828),
.B(n_597),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_834),
.B(n_597),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_703),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_764),
.A2(n_617),
.B(n_613),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_817),
.B(n_603),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_769),
.A2(n_625),
.B(n_619),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_830),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_741),
.A2(n_743),
.B(n_742),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_755),
.A2(n_330),
.B(n_617),
.C(n_614),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_835),
.B(n_603),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_814),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_741),
.A2(n_613),
.B(n_619),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_800),
.A2(n_335),
.B(n_312),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_747),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_704),
.A2(n_667),
.B1(n_321),
.B2(n_347),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_742),
.A2(n_292),
.B(n_200),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_722),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_691),
.B(n_547),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_823),
.B(n_587),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_743),
.A2(n_296),
.B(n_204),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_766),
.A2(n_299),
.B(n_215),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_675),
.B(n_667),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_758),
.B(n_547),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_681),
.B(n_587),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_766),
.A2(n_289),
.B(n_219),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_698),
.A2(n_322),
.B(n_333),
.C(n_346),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_747),
.Y(n_960)
);

INVx11_ASAP7_75t_L g961 ( 
.A(n_798),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_800),
.A2(n_338),
.B(n_341),
.C(n_201),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_771),
.A2(n_273),
.B(n_222),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_688),
.B(n_587),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_771),
.A2(n_287),
.B(n_223),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_835),
.B(n_587),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_829),
.A2(n_313),
.B(n_231),
.C(n_233),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_829),
.A2(n_323),
.B(n_241),
.C(n_242),
.Y(n_968)
);

OAI21xp33_ASAP7_75t_L g969 ( 
.A1(n_821),
.A2(n_194),
.B(n_244),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_749),
.B(n_252),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_705),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_772),
.A2(n_328),
.B(n_262),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_737),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_774),
.A2(n_587),
.B(n_336),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_682),
.A2(n_787),
.B(n_801),
.C(n_802),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_732),
.B(n_587),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_811),
.A2(n_325),
.B1(n_265),
.B2(n_345),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_777),
.Y(n_978)
);

O2A1O1Ixp5_ASAP7_75t_L g979 ( 
.A1(n_818),
.A2(n_626),
.B(n_8),
.C(n_11),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_772),
.A2(n_795),
.B(n_753),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_748),
.B(n_626),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_747),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_732),
.A2(n_324),
.B(n_269),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_836),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_815),
.B(n_254),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_754),
.A2(n_340),
.B(n_337),
.C(n_315),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_753),
.B(n_782),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_762),
.A2(n_7),
.B(n_8),
.C(n_13),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_758),
.B(n_626),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_747),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_778),
.B(n_626),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_832),
.B(n_13),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_820),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_765),
.B(n_16),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_781),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_786),
.A2(n_17),
.B(n_18),
.C(n_21),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_782),
.A2(n_351),
.B(n_23),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_792),
.B(n_794),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_791),
.A2(n_351),
.B(n_26),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_799),
.A2(n_351),
.B(n_27),
.C(n_29),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_791),
.A2(n_351),
.B(n_32),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_795),
.B(n_22),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_776),
.A2(n_85),
.B(n_172),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_730),
.B(n_32),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_779),
.B(n_35),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_793),
.B(n_36),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_803),
.A2(n_36),
.B(n_37),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_804),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_803),
.A2(n_37),
.B(n_38),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_820),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_758),
.B(n_38),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_820),
.B(n_39),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_825),
.B(n_39),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_820),
.B(n_761),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_825),
.B(n_41),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_713),
.B(n_41),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_711),
.B(n_46),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_717),
.B(n_48),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_831),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_867),
.A2(n_724),
.B(n_805),
.Y(n_1020)
);

INVx6_ASAP7_75t_L g1021 ( 
.A(n_861),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_837),
.A2(n_805),
.B(n_783),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_837),
.A2(n_806),
.B(n_812),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_862),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_847),
.A2(n_728),
.B(n_716),
.C(n_713),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_967),
.B(n_784),
.C(n_788),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_887),
.A2(n_728),
.B(n_716),
.C(n_790),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_944),
.B(n_727),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_858),
.A2(n_822),
.B(n_816),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_881),
.B(n_726),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_910),
.A2(n_833),
.B1(n_822),
.B2(n_816),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_943),
.A2(n_833),
.B(n_813),
.C(n_808),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_866),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_970),
.A2(n_813),
.B(n_808),
.C(n_798),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_844),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_882),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_SL g1037 ( 
.A(n_924),
.B(n_50),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_SL g1038 ( 
.A1(n_1011),
.A2(n_51),
.B(n_54),
.C(n_62),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_962),
.A2(n_1015),
.B(n_1013),
.C(n_968),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_SL g1040 ( 
.A1(n_934),
.A2(n_51),
.B1(n_64),
.B2(n_798),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_844),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_925),
.A2(n_798),
.B(n_64),
.C(n_78),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_886),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_940),
.A2(n_76),
.B1(n_80),
.B2(n_83),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1019),
.A2(n_86),
.B1(n_89),
.B2(n_97),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1016),
.A2(n_100),
.B1(n_102),
.B2(n_112),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_857),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_861),
.B(n_880),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_858),
.A2(n_128),
.B(n_133),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_966),
.B(n_134),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_942),
.A2(n_140),
.B(n_146),
.C(n_148),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_883),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_840),
.A2(n_158),
.B(n_159),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_871),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_840),
.A2(n_160),
.B(n_167),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_994),
.A2(n_174),
.B(n_946),
.C(n_902),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_879),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_938),
.B(n_984),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_850),
.B(n_839),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_914),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_854),
.A2(n_868),
.B(n_845),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_874),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_888),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_878),
.B(n_848),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_842),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_923),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_905),
.A2(n_852),
.B1(n_890),
.B2(n_978),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_993),
.B(n_846),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_971),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_894),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_992),
.A2(n_1006),
.B(n_907),
.C(n_855),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_839),
.B(n_842),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_894),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_842),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_893),
.B(n_1012),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_869),
.B(n_876),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_901),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_993),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_908),
.B(n_849),
.Y(n_1079)
);

CKINVDCx16_ASAP7_75t_R g1080 ( 
.A(n_921),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_845),
.A2(n_860),
.B(n_877),
.Y(n_1081)
);

AOI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_948),
.A2(n_904),
.B(n_895),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1012),
.B(n_929),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_950),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_973),
.B(n_995),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_993),
.Y(n_1086)
);

BUFx4f_ASAP7_75t_L g1087 ( 
.A(n_951),
.Y(n_1087)
);

AND2x2_ASAP7_75t_SL g1088 ( 
.A(n_900),
.B(n_903),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_1000),
.A2(n_996),
.B(n_988),
.C(n_959),
.Y(n_1089)
);

BUFx4f_ASAP7_75t_SL g1090 ( 
.A(n_846),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_849),
.B(n_856),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_838),
.A2(n_873),
.B(n_872),
.C(n_851),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_993),
.B(n_856),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_991),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_898),
.B(n_846),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_969),
.B(n_1009),
.C(n_1007),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_SL g1097 ( 
.A(n_951),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_926),
.A2(n_865),
.B1(n_891),
.B2(n_935),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_859),
.B(n_912),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_933),
.A2(n_998),
.B1(n_952),
.B2(n_870),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_860),
.A2(n_877),
.B(n_922),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_985),
.B(n_1008),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_911),
.A2(n_885),
.B(n_920),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_987),
.B(n_936),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_936),
.B(n_947),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_859),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_991),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1004),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_981),
.B(n_1007),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_961),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1009),
.B(n_991),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_859),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1005),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_L g1114 ( 
.A(n_986),
.B(n_975),
.C(n_983),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_947),
.B(n_982),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_841),
.A2(n_843),
.B(n_939),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_912),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_1017),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_885),
.A2(n_920),
.B(n_939),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_912),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_990),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_906),
.A2(n_1002),
.B(n_1018),
.C(n_915),
.Y(n_1122)
);

BUFx8_ASAP7_75t_L g1123 ( 
.A(n_990),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_941),
.A2(n_1001),
.B(n_999),
.C(n_997),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_976),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_960),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_941),
.A2(n_1001),
.B(n_999),
.C(n_997),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_909),
.A2(n_918),
.B(n_932),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_932),
.A2(n_863),
.B(n_853),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_931),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_864),
.A2(n_983),
.B(n_979),
.C(n_928),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_957),
.B(n_964),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_960),
.B(n_1010),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1010),
.B(n_977),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_889),
.B(n_897),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1014),
.B(n_955),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_892),
.A2(n_917),
.B(n_927),
.C(n_930),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_R g1138 ( 
.A(n_955),
.B(n_956),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_899),
.A2(n_963),
.B(n_965),
.C(n_972),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_974),
.A2(n_937),
.B1(n_930),
.B2(n_980),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_913),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_916),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_963),
.B(n_965),
.Y(n_1143)
);

AND2x2_ASAP7_75t_SL g1144 ( 
.A(n_989),
.B(n_884),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_949),
.B(n_953),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1003),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_954),
.B(n_958),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_972),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_916),
.B(n_919),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_919),
.B(n_945),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_896),
.B(n_745),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_875),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_943),
.B(n_680),
.Y(n_1153)
);

INVx8_ASAP7_75t_L g1154 ( 
.A(n_844),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_844),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_861),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_847),
.A2(n_910),
.B1(n_745),
.B2(n_810),
.Y(n_1157)
);

BUFx12f_ASAP7_75t_L g1158 ( 
.A(n_924),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_847),
.B(n_745),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_L g1160 ( 
.A1(n_892),
.A2(n_917),
.B(n_927),
.C(n_851),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_866),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_928),
.A2(n_941),
.B(n_672),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_861),
.B(n_709),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_867),
.A2(n_729),
.B(n_694),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_847),
.B(n_745),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_875),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1168)
);

BUFx4_ASAP7_75t_SL g1169 ( 
.A(n_1043),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1153),
.A2(n_1103),
.B(n_1101),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1159),
.B(n_1165),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1157),
.B(n_1135),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1085),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1059),
.A2(n_1052),
.B1(n_1058),
.B2(n_1057),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1137),
.A2(n_1025),
.B(n_1160),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1088),
.B(n_1064),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1023),
.A2(n_1029),
.B(n_1146),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1088),
.B(n_1058),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1146),
.A2(n_1061),
.B(n_1128),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1124),
.A2(n_1127),
.A3(n_1100),
.B(n_1150),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1154),
.Y(n_1182)
);

BUFx12f_ASAP7_75t_L g1183 ( 
.A(n_1158),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_1096),
.A2(n_1114),
.B1(n_1113),
.B2(n_1108),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1022),
.A2(n_1149),
.B(n_1162),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1057),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1039),
.A2(n_1071),
.B(n_1056),
.C(n_1089),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_L g1188 ( 
.A(n_1099),
.B(n_1078),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1150),
.A2(n_1032),
.A3(n_1132),
.B(n_1034),
.Y(n_1189)
);

O2A1O1Ixp5_ASAP7_75t_L g1190 ( 
.A1(n_1149),
.A2(n_1137),
.B(n_1160),
.C(n_1145),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1164),
.A2(n_1122),
.B(n_1067),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1123),
.Y(n_1192)
);

AO21x1_ASAP7_75t_L g1193 ( 
.A1(n_1096),
.A2(n_1082),
.B(n_1139),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1151),
.A2(n_1147),
.B(n_1092),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1132),
.A2(n_1031),
.A3(n_1136),
.B(n_1130),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1111),
.A2(n_1109),
.B1(n_1118),
.B2(n_1075),
.Y(n_1196)
);

AO21x1_ASAP7_75t_L g1197 ( 
.A1(n_1050),
.A2(n_1136),
.B(n_1095),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1141),
.A2(n_1142),
.B(n_1131),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1141),
.A2(n_1142),
.B(n_1144),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1080),
.A2(n_1059),
.B1(n_1027),
.B2(n_1040),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1036),
.B(n_1048),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1154),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1083),
.B(n_1102),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1144),
.A2(n_1140),
.B(n_1055),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1024),
.B(n_1062),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1094),
.A2(n_1107),
.B1(n_1087),
.B2(n_1046),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1063),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1051),
.A2(n_1166),
.A3(n_1069),
.B(n_1152),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1033),
.B(n_1072),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1049),
.A2(n_1053),
.B(n_1140),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1020),
.A2(n_1143),
.B(n_1050),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1026),
.A2(n_1118),
.B(n_1042),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1038),
.A2(n_1163),
.B(n_1079),
.C(n_1076),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1156),
.B(n_1099),
.Y(n_1215)
);

BUFx10_ASAP7_75t_L g1216 ( 
.A(n_1048),
.Y(n_1216)
);

NAND2x1_ASAP7_75t_L g1217 ( 
.A(n_1078),
.B(n_1112),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1154),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1161),
.B(n_1054),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1104),
.A2(n_1105),
.B(n_1115),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_1110),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1066),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1097),
.A2(n_1134),
.B(n_1078),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1065),
.B(n_1074),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1028),
.A2(n_1079),
.A3(n_1045),
.B(n_1076),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1097),
.A2(n_1078),
.B(n_1077),
.Y(n_1226)
);

CKINVDCx8_ASAP7_75t_R g1227 ( 
.A(n_1030),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1026),
.A2(n_1091),
.B(n_1093),
.C(n_1125),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1068),
.A2(n_1133),
.B(n_1046),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1155),
.B(n_1041),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1035),
.B(n_1041),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1091),
.A2(n_1044),
.B(n_1117),
.Y(n_1232)
);

AOI31xp67_ASAP7_75t_L g1233 ( 
.A1(n_1148),
.A2(n_1138),
.A3(n_1117),
.B(n_1106),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1086),
.A2(n_1112),
.B(n_1106),
.Y(n_1234)
);

AOI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1086),
.A2(n_1126),
.B(n_1030),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1028),
.A2(n_1156),
.A3(n_1138),
.B(n_1030),
.Y(n_1236)
);

INVx3_ASAP7_75t_SL g1237 ( 
.A(n_1021),
.Y(n_1237)
);

AOI221xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1106),
.A2(n_1112),
.B1(n_1035),
.B2(n_1041),
.C(n_1037),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1106),
.A2(n_1112),
.A3(n_1060),
.B(n_1121),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1087),
.A2(n_1120),
.B(n_1155),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1035),
.A2(n_1041),
.B(n_1090),
.Y(n_1241)
);

AO21x1_ASAP7_75t_L g1242 ( 
.A1(n_1021),
.A2(n_1153),
.B(n_1096),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_1052),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1084),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1025),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1058),
.B(n_719),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1159),
.A2(n_1015),
.B1(n_1013),
.B2(n_1165),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1081),
.A2(n_1119),
.B(n_1137),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1058),
.B(n_719),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1084),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1025),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1025),
.A2(n_1153),
.B(n_1100),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1052),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1085),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1081),
.A2(n_1101),
.B(n_1103),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1081),
.A2(n_1101),
.B(n_1103),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1059),
.B(n_709),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1159),
.B(n_1165),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1154),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1153),
.A2(n_847),
.B(n_1039),
.C(n_1071),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1158),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1036),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1025),
.Y(n_1273)
);

OAI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1159),
.A2(n_1015),
.B1(n_1013),
.B2(n_1165),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1154),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1084),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1123),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1153),
.A2(n_847),
.B(n_1039),
.C(n_1071),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1123),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1157),
.B(n_1135),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1085),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1154),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1153),
.A2(n_1096),
.B(n_1100),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1159),
.B(n_1165),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1124),
.A2(n_927),
.A3(n_917),
.B(n_892),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1153),
.A2(n_847),
.B(n_1039),
.C(n_1071),
.Y(n_1288)
);

NOR2x1_ASAP7_75t_L g1289 ( 
.A(n_1120),
.B(n_1047),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1058),
.B(n_719),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1085),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1025),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_L g1294 ( 
.A(n_1153),
.B(n_847),
.C(n_970),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1153),
.A2(n_1159),
.B(n_1165),
.C(n_1157),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1084),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_1135),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1124),
.A2(n_927),
.A3(n_917),
.B(n_892),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1059),
.B(n_709),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1157),
.B(n_1135),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1153),
.A2(n_847),
.B1(n_1165),
.B2(n_1159),
.C(n_1157),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1081),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1153),
.A2(n_1098),
.B(n_1129),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1123),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1057),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1085),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1059),
.B(n_709),
.Y(n_1310)
);

AO32x2_ASAP7_75t_L g1311 ( 
.A1(n_1157),
.A2(n_1100),
.A3(n_1098),
.B1(n_1067),
.B2(n_1031),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1057),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1159),
.B(n_1165),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1036),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1153),
.A2(n_910),
.B1(n_1157),
.B2(n_1135),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1124),
.A2(n_927),
.A3(n_917),
.B(n_892),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1217),
.B(n_1231),
.Y(n_1317)
);

OAI22x1_ASAP7_75t_L g1318 ( 
.A1(n_1294),
.A2(n_1174),
.B1(n_1286),
.B2(n_1313),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1205),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1205),
.Y(n_1320)
);

BUFx2_ASAP7_75t_R g1321 ( 
.A(n_1278),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1303),
.A2(n_1274),
.B1(n_1247),
.B2(n_1200),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1303),
.A2(n_1200),
.B1(n_1281),
.B2(n_1302),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1237),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1271),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1308),
.A2(n_1312),
.B1(n_1313),
.B2(n_1171),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1186),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1267),
.A2(n_1171),
.B1(n_1286),
.B2(n_1288),
.Y(n_1328)
);

BUFx4_ASAP7_75t_R g1329 ( 
.A(n_1216),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1247),
.A2(n_1274),
.B1(n_1315),
.B2(n_1302),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1183),
.Y(n_1331)
);

INVx3_ASAP7_75t_SL g1332 ( 
.A(n_1243),
.Y(n_1332)
);

CKINVDCx9p33_ASAP7_75t_R g1333 ( 
.A(n_1172),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1315),
.A2(n_1281),
.B1(n_1172),
.B2(n_1285),
.Y(n_1334)
);

INVx5_ASAP7_75t_L g1335 ( 
.A(n_1218),
.Y(n_1335)
);

CKINVDCx6p67_ASAP7_75t_R g1336 ( 
.A(n_1280),
.Y(n_1336)
);

CKINVDCx6p67_ASAP7_75t_R g1337 ( 
.A(n_1306),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1246),
.A2(n_1251),
.B1(n_1290),
.B2(n_1184),
.Y(n_1338)
);

CKINVDCx6p67_ASAP7_75t_R g1339 ( 
.A(n_1237),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1203),
.B(n_1296),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1179),
.A2(n_1293),
.B1(n_1245),
.B2(n_1273),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1207),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1203),
.B(n_1296),
.Y(n_1343)
);

INVx6_ASAP7_75t_L g1344 ( 
.A(n_1218),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1221),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1222),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1270),
.A2(n_1279),
.B(n_1213),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1221),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1173),
.B(n_1259),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1184),
.A2(n_1293),
.B1(n_1273),
.B2(n_1255),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1283),
.B(n_1291),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1184),
.A2(n_1255),
.B1(n_1245),
.B2(n_1179),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1169),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1201),
.A2(n_1310),
.B1(n_1301),
.B2(n_1266),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1196),
.A2(n_1213),
.B1(n_1176),
.B2(n_1309),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1244),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1268),
.Y(n_1357)
);

BUFx2_ASAP7_75t_SL g1358 ( 
.A(n_1192),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1210),
.B(n_1219),
.Y(n_1359)
);

BUFx8_ASAP7_75t_SL g1360 ( 
.A(n_1258),
.Y(n_1360)
);

INVx5_ASAP7_75t_L g1361 ( 
.A(n_1268),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1196),
.A2(n_1206),
.B1(n_1298),
.B2(n_1232),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1168),
.B(n_1209),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1196),
.A2(n_1206),
.B1(n_1298),
.B2(n_1232),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1216),
.Y(n_1365)
);

BUFx4_ASAP7_75t_R g1366 ( 
.A(n_1257),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1272),
.Y(n_1367)
);

INVx3_ASAP7_75t_SL g1368 ( 
.A(n_1250),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1289),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1314),
.B(n_1176),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1175),
.A2(n_1253),
.B1(n_1297),
.B2(n_1277),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1238),
.A2(n_1230),
.B1(n_1197),
.B2(n_1187),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1307),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1227),
.Y(n_1374)
);

INVx6_ASAP7_75t_L g1375 ( 
.A(n_1268),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1250),
.A2(n_1256),
.B1(n_1175),
.B2(n_1169),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1275),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1193),
.A2(n_1242),
.B1(n_1191),
.B2(n_1305),
.Y(n_1378)
);

CKINVDCx11_ASAP7_75t_R g1379 ( 
.A(n_1275),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1230),
.A2(n_1224),
.B1(n_1215),
.B2(n_1256),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1275),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1191),
.A2(n_1167),
.B(n_1292),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1182),
.B(n_1202),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1188),
.Y(n_1384)
);

BUFx2_ASAP7_75t_SL g1385 ( 
.A(n_1182),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1208),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1226),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1167),
.A2(n_1300),
.B1(n_1292),
.B2(n_1305),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1254),
.A2(n_1300),
.B1(n_1264),
.B2(n_1263),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1223),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1202),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1254),
.A2(n_1269),
.B1(n_1263),
.B2(n_1264),
.Y(n_1392)
);

OAI22x1_ASAP7_75t_L g1393 ( 
.A1(n_1235),
.A2(n_1284),
.B1(n_1311),
.B2(n_1214),
.Y(n_1393)
);

BUFx4f_ASAP7_75t_SL g1394 ( 
.A(n_1284),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1233),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1269),
.A2(n_1204),
.B1(n_1194),
.B2(n_1311),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1214),
.A2(n_1204),
.B(n_1199),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1241),
.B(n_1236),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1311),
.A2(n_1194),
.B1(n_1212),
.B2(n_1225),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1239),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1248),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1181),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1311),
.A2(n_1199),
.B1(n_1198),
.B2(n_1240),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1241),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1239),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1240),
.A2(n_1198),
.B1(n_1170),
.B2(n_1220),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1228),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1225),
.A2(n_1211),
.B1(n_1229),
.B2(n_1189),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1185),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1220),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1170),
.A2(n_1228),
.B1(n_1248),
.B2(n_1234),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1189),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1234),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1189),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1225),
.A2(n_1181),
.B1(n_1195),
.B2(n_1190),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1262),
.A2(n_1265),
.B1(n_1195),
.B2(n_1181),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1265),
.A2(n_1195),
.B1(n_1190),
.B2(n_1261),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1287),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1299),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1299),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1316),
.A2(n_1177),
.B1(n_1304),
.B2(n_1295),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1316),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1180),
.A2(n_1276),
.B1(n_1249),
.B2(n_1252),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1316),
.A2(n_1178),
.B1(n_1260),
.B2(n_1282),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1201),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1153),
.B2(n_1274),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1200),
.B2(n_1281),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1271),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1294),
.A2(n_739),
.B1(n_355),
.B2(n_370),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1153),
.B2(n_1274),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1153),
.B2(n_1274),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1237),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1153),
.B2(n_1274),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1153),
.B2(n_1274),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1205),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1219),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1237),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1294),
.A2(n_1303),
.B1(n_1165),
.B2(n_1159),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1323),
.A2(n_1347),
.B1(n_1328),
.B2(n_1427),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1370),
.B(n_1340),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1333),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1323),
.A2(n_1322),
.B1(n_1418),
.B2(n_1407),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1322),
.A2(n_1330),
.B(n_1426),
.C(n_1430),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1409),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1319),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1409),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1410),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1343),
.B(n_1320),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1419),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1421),
.A2(n_1382),
.B(n_1392),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1411),
.A2(n_1388),
.B(n_1406),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1350),
.B(n_1338),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1422),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1402),
.B(n_1352),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1420),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1358),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1413),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

INVx5_ASAP7_75t_L g1459 ( 
.A(n_1409),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1405),
.B(n_1398),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1352),
.B(n_1412),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1414),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1388),
.A2(n_1406),
.B(n_1417),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1417),
.A2(n_1416),
.B(n_1378),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1409),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1427),
.A2(n_1438),
.B1(n_1330),
.B2(n_1433),
.C(n_1431),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1435),
.Y(n_1467)
);

OR2x6_ASAP7_75t_L g1468 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1429),
.A2(n_1338),
.B1(n_1433),
.B2(n_1430),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1400),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1333),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1342),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1416),
.A2(n_1378),
.B(n_1386),
.Y(n_1473)
);

AOI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1393),
.A2(n_1318),
.B(n_1369),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1346),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1401),
.B(n_1372),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1359),
.B(n_1334),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1415),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1401),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1334),
.B(n_1399),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1426),
.A2(n_1434),
.B1(n_1431),
.B2(n_1362),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1415),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1434),
.A2(n_1371),
.B(n_1317),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1355),
.B(n_1324),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1355),
.B(n_1341),
.Y(n_1485)
);

INVx8_ASAP7_75t_L g1486 ( 
.A(n_1384),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1341),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1371),
.A2(n_1317),
.B(n_1391),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1403),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1403),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1396),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1396),
.A2(n_1349),
.B(n_1351),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1356),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1354),
.A2(n_1326),
.B1(n_1389),
.B2(n_1364),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1408),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1424),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1436),
.B(n_1425),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1367),
.A2(n_1380),
.B(n_1437),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1329),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1423),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1366),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1404),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1391),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1324),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1383),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1390),
.A2(n_1387),
.B1(n_1425),
.B2(n_1376),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1329),
.A2(n_1373),
.B(n_1385),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1432),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1381),
.A2(n_1374),
.B1(n_1332),
.B2(n_1337),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1365),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1363),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1363),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1432),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1437),
.Y(n_1515)
);

BUFx2_ASAP7_75t_SL g1516 ( 
.A(n_1335),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1344),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1368),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1339),
.A2(n_1368),
.B1(n_1332),
.B2(n_1394),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1377),
.B(n_1336),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1344),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1345),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1394),
.A2(n_1375),
.B(n_1344),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1472),
.Y(n_1524)
);

INVx5_ASAP7_75t_L g1525 ( 
.A(n_1468),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_SL g1526 ( 
.A1(n_1439),
.A2(n_1348),
.B(n_1353),
.C(n_1360),
.Y(n_1526)
);

O2A1O1Ixp33_ASAP7_75t_SL g1527 ( 
.A1(n_1443),
.A2(n_1379),
.B(n_1321),
.C(n_1327),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1466),
.A2(n_1335),
.B(n_1361),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1494),
.A2(n_1331),
.B(n_1357),
.C(n_1375),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1481),
.A2(n_1335),
.B(n_1361),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1450),
.A2(n_1451),
.B(n_1463),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_L g1532 ( 
.A(n_1518),
.B(n_1335),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1475),
.B(n_1325),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_R g1534 ( 
.A(n_1441),
.B(n_1471),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1496),
.B(n_1361),
.C(n_1428),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1445),
.B(n_1357),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1442),
.A2(n_1469),
.B1(n_1480),
.B2(n_1485),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1450),
.A2(n_1451),
.B(n_1463),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1491),
.B(n_1489),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1468),
.A2(n_1441),
.B(n_1471),
.Y(n_1540)
);

A2O1A1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1485),
.A2(n_1480),
.B(n_1490),
.C(n_1452),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1490),
.A2(n_1452),
.B(n_1487),
.C(n_1483),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1477),
.B(n_1496),
.Y(n_1543)
);

O2A1O1Ixp33_ASAP7_75t_SL g1544 ( 
.A1(n_1499),
.A2(n_1519),
.B(n_1456),
.C(n_1515),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1467),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

AO21x2_ASAP7_75t_L g1547 ( 
.A1(n_1478),
.A2(n_1482),
.B(n_1500),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1520),
.B(n_1522),
.Y(n_1548)
);

AND2x6_ASAP7_75t_L g1549 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1493),
.Y(n_1550)
);

NAND2xp33_ASAP7_75t_R g1551 ( 
.A(n_1523),
.B(n_1468),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1510),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1497),
.B(n_1505),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1492),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1484),
.A2(n_1495),
.B1(n_1501),
.B2(n_1502),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1509),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1484),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1440),
.B(n_1448),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_SL g1559 ( 
.A(n_1516),
.B(n_1511),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1487),
.A2(n_1476),
.B(n_1468),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1510),
.A2(n_1468),
.B1(n_1507),
.B2(n_1511),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1482),
.A2(n_1500),
.B(n_1495),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1476),
.A2(n_1474),
.B(n_1464),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1484),
.B(n_1503),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1484),
.B(n_1503),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_SL g1566 ( 
.A(n_1498),
.B(n_1521),
.C(n_1517),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1511),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1523),
.A2(n_1508),
.B(n_1457),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1464),
.B(n_1454),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1512),
.A2(n_1513),
.B1(n_1514),
.B2(n_1518),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1486),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1454),
.B(n_1461),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1493),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1486),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1461),
.B(n_1447),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1460),
.B(n_1473),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1447),
.B(n_1444),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1474),
.A2(n_1483),
.B(n_1488),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1473),
.A2(n_1488),
.B(n_1479),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1459),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1517),
.B(n_1521),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1455),
.A2(n_1458),
.B1(n_1462),
.B2(n_1449),
.C(n_1453),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1558),
.B(n_1458),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1531),
.B(n_1446),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1550),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1573),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1538),
.B(n_1569),
.Y(n_1589)
);

NAND2x1_ASAP7_75t_L g1590 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1575),
.B(n_1460),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1540),
.B(n_1518),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1554),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1524),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1546),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1575),
.B(n_1462),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1545),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1534),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1577),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1549),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1459),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1539),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1539),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1449),
.Y(n_1605)
);

NOR2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1535),
.B(n_1457),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1538),
.B(n_1569),
.Y(n_1607)
);

INVx5_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1577),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_1525),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1579),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1544),
.B(n_1504),
.Y(n_1612)
);

INVx8_ASAP7_75t_L g1613 ( 
.A(n_1525),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1572),
.B(n_1465),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1549),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1572),
.B(n_1465),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1556),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1553),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1589),
.B(n_1543),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1589),
.B(n_1557),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1607),
.B(n_1547),
.Y(n_1623)
);

INVx5_ASAP7_75t_SL g1624 ( 
.A(n_1602),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_L g1625 ( 
.A1(n_1595),
.A2(n_1541),
.B(n_1537),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1583),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1599),
.B(n_1552),
.Y(n_1627)
);

OAI31xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1595),
.A2(n_1566),
.A3(n_1534),
.B(n_1560),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1601),
.Y(n_1629)
);

OAI31xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1612),
.A2(n_1563),
.A3(n_1570),
.B(n_1528),
.Y(n_1630)
);

OAI31xp33_ASAP7_75t_L g1631 ( 
.A1(n_1606),
.A2(n_1541),
.A3(n_1527),
.B(n_1529),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1601),
.Y(n_1632)
);

INVx5_ASAP7_75t_SL g1633 ( 
.A(n_1602),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1599),
.A2(n_1561),
.B1(n_1542),
.B2(n_1555),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1583),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1607),
.B(n_1576),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1576),
.Y(n_1637)
);

AO21x2_ASAP7_75t_L g1638 ( 
.A1(n_1611),
.A2(n_1578),
.B(n_1542),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1615),
.B(n_1576),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1611),
.Y(n_1641)
);

INVx5_ASAP7_75t_L g1642 ( 
.A(n_1613),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1583),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1605),
.A2(n_1527),
.B1(n_1526),
.B2(n_1562),
.C(n_1547),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1587),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1588),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1584),
.B(n_1562),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1586),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1602),
.Y(n_1649)
);

OAI33xp33_ASAP7_75t_L g1650 ( 
.A1(n_1605),
.A2(n_1533),
.A3(n_1536),
.B1(n_1504),
.B2(n_1453),
.B3(n_1470),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1525),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1585),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1591),
.A2(n_1525),
.B1(n_1567),
.B2(n_1518),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1585),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1526),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1585),
.Y(n_1656)
);

AOI211xp5_ASAP7_75t_L g1657 ( 
.A1(n_1592),
.A2(n_1530),
.B(n_1548),
.C(n_1559),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1590),
.A2(n_1551),
.B1(n_1457),
.B2(n_1581),
.C(n_1525),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1619),
.B(n_1594),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1600),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1629),
.B(n_1608),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1630),
.B(n_1592),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1619),
.B(n_1594),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1652),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1620),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1629),
.B(n_1606),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1651),
.B(n_1590),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1645),
.B(n_1598),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1621),
.B(n_1600),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1645),
.Y(n_1671)
);

AND2x2_ASAP7_75t_SL g1672 ( 
.A(n_1628),
.B(n_1610),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1625),
.A2(n_1565),
.B1(n_1564),
.B2(n_1608),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1646),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1623),
.B(n_1597),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1646),
.B(n_1598),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1623),
.B(n_1597),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1622),
.B(n_1609),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1622),
.B(n_1609),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1627),
.B(n_1603),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1622),
.B(n_1614),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1627),
.B(n_1603),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1614),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1639),
.Y(n_1685)
);

AND2x4_ASAP7_75t_SL g1686 ( 
.A(n_1637),
.B(n_1602),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1629),
.B(n_1616),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1652),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1652),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1639),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1639),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1618),
.B(n_1596),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1652),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1659),
.B(n_1647),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1662),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1662),
.B(n_1630),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1688),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1688),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1688),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1665),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1666),
.B(n_1633),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1665),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1694),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1633),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1694),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1686),
.B(n_1633),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1671),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1694),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1680),
.B(n_1655),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1671),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1674),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1672),
.B(n_1642),
.Y(n_1716)
);

OR2x6_ASAP7_75t_L g1717 ( 
.A(n_1668),
.B(n_1625),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1659),
.B(n_1626),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1669),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1663),
.B(n_1626),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1686),
.B(n_1633),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1672),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1690),
.A2(n_1634),
.B1(n_1655),
.B2(n_1658),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1672),
.B(n_1628),
.Y(n_1724)
);

INVx3_ASAP7_75t_SL g1725 ( 
.A(n_1672),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1669),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1686),
.B(n_1633),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1663),
.B(n_1635),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1694),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1644),
.C(n_1631),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1690),
.A2(n_1650),
.B1(n_1644),
.B2(n_1634),
.C(n_1643),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1676),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1680),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1682),
.B(n_1617),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1668),
.B(n_1661),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1676),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1686),
.B(n_1633),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1697),
.A2(n_1638),
.B1(n_1631),
.B2(n_1650),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1701),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1696),
.B(n_1682),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1712),
.B(n_1693),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1567),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1733),
.B(n_1693),
.Y(n_1743)
);

NOR2x1_ASAP7_75t_L g1744 ( 
.A(n_1722),
.B(n_1661),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1730),
.A2(n_1638),
.B1(n_1657),
.B2(n_1673),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1725),
.B(n_1683),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1701),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1731),
.B(n_1693),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1725),
.B(n_1683),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1725),
.B(n_1661),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1734),
.B(n_1660),
.Y(n_1751)
);

AND2x2_ASAP7_75t_SL g1752 ( 
.A(n_1702),
.B(n_1661),
.Y(n_1752)
);

A2O1A1Ixp33_ASAP7_75t_SL g1753 ( 
.A1(n_1702),
.A2(n_1657),
.B(n_1688),
.C(n_1664),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1718),
.B(n_1675),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1723),
.B(n_1692),
.C(n_1658),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1718),
.B(n_1675),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1675),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1703),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1703),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1698),
.A2(n_1691),
.B(n_1685),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1717),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1719),
.B(n_1726),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1717),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1706),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1698),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1706),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1707),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1723),
.B(n_1571),
.Y(n_1769)
);

OAI332xp33_ASAP7_75t_L g1770 ( 
.A1(n_1695),
.A2(n_1677),
.A3(n_1684),
.B1(n_1691),
.B2(n_1685),
.B3(n_1648),
.C1(n_1632),
.C2(n_1593),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1709),
.B(n_1687),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1716),
.B(n_1649),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1720),
.B(n_1677),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1709),
.B(n_1687),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1738),
.A2(n_1748),
.B1(n_1753),
.B2(n_1756),
.C(n_1745),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1769),
.A2(n_1717),
.B1(n_1742),
.B2(n_1638),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1740),
.A2(n_1717),
.B1(n_1716),
.B2(n_1673),
.Y(n_1777)
);

AOI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1753),
.A2(n_1695),
.B1(n_1736),
.B2(n_1732),
.C(n_1719),
.Y(n_1778)
);

AOI21xp33_ASAP7_75t_L g1779 ( 
.A1(n_1739),
.A2(n_1717),
.B(n_1726),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1770),
.A2(n_1705),
.B(n_1716),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1763),
.A2(n_1732),
.B1(n_1736),
.B2(n_1704),
.C(n_1729),
.Y(n_1781)
);

NAND3x1_ASAP7_75t_L g1782 ( 
.A(n_1744),
.B(n_1705),
.C(n_1721),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1741),
.B(n_1660),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1739),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1768),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1743),
.B(n_1728),
.Y(n_1786)
);

NAND4xp75_ASAP7_75t_L g1787 ( 
.A(n_1750),
.B(n_1752),
.C(n_1746),
.D(n_1749),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1752),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1750),
.A2(n_1727),
.B(n_1721),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1746),
.A2(n_1737),
.B(n_1727),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1768),
.Y(n_1791)
);

NOR2xp67_ASAP7_75t_L g1792 ( 
.A(n_1749),
.B(n_1737),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1754),
.B(n_1660),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1762),
.A2(n_1638),
.B1(n_1735),
.B2(n_1661),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1754),
.B(n_1687),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1764),
.A2(n_1636),
.B(n_1728),
.C(n_1635),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1755),
.A2(n_1735),
.B1(n_1668),
.B2(n_1643),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1755),
.B(n_1670),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1747),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1766),
.A2(n_1638),
.B1(n_1636),
.B2(n_1640),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1775),
.A2(n_1735),
.B(n_1761),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1776),
.A2(n_1766),
.B1(n_1761),
.B2(n_1758),
.C(n_1773),
.Y(n_1802)
);

NAND3xp33_ASAP7_75t_SL g1803 ( 
.A(n_1788),
.B(n_1758),
.C(n_1757),
.Y(n_1803)
);

OAI22x1_ASAP7_75t_L g1804 ( 
.A1(n_1800),
.A2(n_1772),
.B1(n_1759),
.B2(n_1767),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1787),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1795),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1778),
.B(n_1760),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1782),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1792),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1757),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1794),
.A2(n_1761),
.B1(n_1771),
.B2(n_1774),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1784),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1785),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1799),
.B(n_1765),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1798),
.B(n_1773),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1779),
.A2(n_1774),
.B(n_1771),
.C(n_1751),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1791),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1781),
.B(n_1707),
.Y(n_1818)
);

AOI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1779),
.A2(n_1710),
.B(n_1713),
.C(n_1715),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_R g1820 ( 
.A(n_1793),
.B(n_1571),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1810),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1805),
.B(n_1797),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1809),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1814),
.Y(n_1824)
);

XOR2xp5_ASAP7_75t_L g1825 ( 
.A(n_1803),
.B(n_1777),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1806),
.B(n_1783),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1807),
.A2(n_1777),
.B1(n_1780),
.B2(n_1796),
.C(n_1789),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1801),
.A2(n_1807),
.B1(n_1802),
.B2(n_1818),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1811),
.A2(n_1790),
.B1(n_1700),
.B2(n_1729),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1804),
.A2(n_1699),
.B1(n_1700),
.B2(n_1711),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1815),
.B(n_1710),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1814),
.Y(n_1832)
);

NOR2xp67_ASAP7_75t_SL g1833 ( 
.A(n_1821),
.B(n_1808),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1824),
.B(n_1816),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_L g1835 ( 
.A1(n_1827),
.A2(n_1819),
.B(n_1818),
.C(n_1820),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1832),
.B(n_1812),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1823),
.B(n_1813),
.Y(n_1837)
);

OAI211xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1828),
.A2(n_1817),
.B(n_1715),
.C(n_1714),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1825),
.B(n_1831),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1826),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1822),
.B(n_1713),
.Y(n_1841)
);

XOR2x2_ASAP7_75t_L g1842 ( 
.A(n_1839),
.B(n_1829),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1833),
.B(n_1830),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1838),
.A2(n_1704),
.B1(n_1711),
.B2(n_1708),
.C(n_1699),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1835),
.B(n_1735),
.C(n_1708),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_L g1846 ( 
.A(n_1841),
.B(n_1574),
.Y(n_1846)
);

AOI222xp33_ASAP7_75t_L g1847 ( 
.A1(n_1843),
.A2(n_1834),
.B1(n_1837),
.B2(n_1836),
.C1(n_1840),
.C2(n_1714),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1842),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1845),
.A2(n_1735),
.B1(n_1668),
.B2(n_1677),
.C(n_1664),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1844),
.A2(n_1654),
.B1(n_1689),
.B2(n_1664),
.C(n_1639),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1846),
.A2(n_1668),
.B1(n_1689),
.B2(n_1684),
.C(n_1654),
.Y(n_1851)
);

NAND3xp33_ASAP7_75t_L g1852 ( 
.A(n_1843),
.B(n_1668),
.C(n_1632),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1848),
.B(n_1689),
.Y(n_1853)
);

NOR3xp33_ASAP7_75t_L g1854 ( 
.A(n_1849),
.B(n_1641),
.C(n_1574),
.Y(n_1854)
);

NAND4xp75_ASAP7_75t_L g1855 ( 
.A(n_1850),
.B(n_1640),
.C(n_1637),
.D(n_1632),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1852),
.B(n_1684),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1847),
.Y(n_1857)
);

AND4x1_ASAP7_75t_L g1858 ( 
.A(n_1857),
.B(n_1851),
.C(n_1670),
.D(n_1681),
.Y(n_1858)
);

NOR3xp33_ASAP7_75t_SL g1859 ( 
.A(n_1853),
.B(n_1653),
.C(n_1551),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1856),
.B(n_1854),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1858),
.B(n_1855),
.Y(n_1861)
);

OA22x2_ASAP7_75t_L g1862 ( 
.A1(n_1861),
.A2(n_1860),
.B1(n_1859),
.B2(n_1617),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1862),
.Y(n_1863)
);

AO22x2_ASAP7_75t_L g1864 ( 
.A1(n_1862),
.A2(n_1648),
.B1(n_1670),
.B2(n_1681),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1863),
.A2(n_1648),
.B1(n_1679),
.B2(n_1678),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1864),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1866),
.A2(n_1641),
.B1(n_1656),
.B2(n_1636),
.C(n_1679),
.Y(n_1867)
);

OAI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1865),
.A2(n_1668),
.B1(n_1656),
.B2(n_1486),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1486),
.B(n_1679),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1869),
.A2(n_1867),
.B(n_1640),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1870),
.A2(n_1486),
.B1(n_1656),
.B2(n_1678),
.Y(n_1871)
);

OAI221xp5_ASAP7_75t_R g1872 ( 
.A1(n_1871),
.A2(n_1633),
.B1(n_1624),
.B2(n_1649),
.C(n_1681),
.Y(n_1872)
);

AOI211xp5_ASAP7_75t_L g1873 ( 
.A1(n_1872),
.A2(n_1532),
.B(n_1518),
.C(n_1653),
.Y(n_1873)
);


endmodule