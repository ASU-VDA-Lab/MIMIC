module fake_jpeg_4903_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_23),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_42),
.B(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_60),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_57),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_39),
.C(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_33),
.B1(n_44),
.B2(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_7),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_26),
.B1(n_29),
.B2(n_19),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_37),
.B1(n_33),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_67),
.A2(n_71),
.B1(n_68),
.B2(n_98),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_33),
.B1(n_40),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_110)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_70),
.B(n_73),
.Y(n_133)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_75),
.B(n_78),
.Y(n_140)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_85),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_57),
.B1(n_28),
.B2(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_106),
.B1(n_96),
.B2(n_83),
.Y(n_113)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_29),
.B1(n_34),
.B2(n_38),
.Y(n_86)
);

NAND2x1_ASAP7_75t_SL g142 ( 
.A(n_87),
.B(n_6),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_32),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_48),
.B(n_22),
.Y(n_95)
);

NAND5xp2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_22),
.C(n_17),
.D(n_2),
.E(n_3),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_100),
.Y(n_125)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_59),
.B(n_31),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_45),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_47),
.A2(n_31),
.B1(n_25),
.B2(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_113),
.B1(n_116),
.B2(n_132),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_111),
.A2(n_145),
.B(n_141),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_22),
.B1(n_17),
.B2(n_2),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_134),
.B1(n_71),
.B2(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_17),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g126 ( 
.A(n_95),
.Y(n_126)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_17),
.Y(n_127)
);

XNOR2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_67),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_81),
.A2(n_5),
.B1(n_11),
.B2(n_9),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_141),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_75),
.C(n_73),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_92),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_144),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_3),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_76),
.B1(n_74),
.B2(n_79),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_4),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_80),
.A2(n_11),
.B(n_13),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_149),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g209 ( 
.A(n_147),
.B(n_157),
.C(n_165),
.Y(n_209)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_92),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_155),
.B(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_153),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_91),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_171),
.Y(n_197)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_128),
.B1(n_134),
.B2(n_115),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_159),
.Y(n_210)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_70),
.A3(n_103),
.B1(n_108),
.B2(n_64),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_120),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_77),
.C(n_88),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_181),
.C(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_167),
.B(n_174),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_105),
.B1(n_85),
.B2(n_97),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_169),
.B1(n_115),
.B2(n_114),
.Y(n_191)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_72),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_131),
.B(n_145),
.Y(n_183)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_179),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_74),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_79),
.C(n_112),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_142),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_214),
.B(n_177),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_186),
.B1(n_188),
.B2(n_200),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_136),
.B1(n_120),
.B2(n_112),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_125),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_201),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_118),
.C(n_130),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_130),
.C(n_111),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_142),
.B1(n_111),
.B2(n_128),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_198),
.A2(n_205),
.B1(n_185),
.B2(n_209),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_117),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_137),
.B1(n_114),
.B2(n_117),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_207),
.B1(n_212),
.B2(n_214),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_150),
.B1(n_180),
.B2(n_156),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_178),
.B1(n_153),
.B2(n_159),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_139),
.B1(n_147),
.B2(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_149),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_147),
.A2(n_180),
.B1(n_170),
.B2(n_156),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_150),
.B(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_214),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_155),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_219),
.B(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_203),
.B(n_177),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_227),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_230),
.B(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_229),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_169),
.C(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_237),
.C(n_186),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_198),
.B1(n_196),
.B2(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_184),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_185),
.C(n_193),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_223),
.Y(n_261)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_188),
.B(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_256),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_255),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_247),
.B1(n_239),
.B2(n_240),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_233),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_258),
.C(n_232),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_189),
.B(n_212),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_203),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_200),
.B1(n_183),
.B2(n_184),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_187),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_273),
.C(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_241),
.B1(n_257),
.B2(n_230),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_276),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_258),
.C(n_224),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_237),
.C(n_226),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_217),
.Y(n_276)
);

INVxp33_ASAP7_75t_SL g277 ( 
.A(n_248),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_228),
.B1(n_236),
.B2(n_220),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_255),
.B(n_251),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_286),
.B(n_289),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_246),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_288),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_247),
.C(n_252),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_241),
.B(n_243),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_270),
.A2(n_215),
.B1(n_222),
.B2(n_247),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_259),
.B1(n_266),
.B2(n_249),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_266),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_279),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_269),
.C(n_273),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_296),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_274),
.C(n_275),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_259),
.B1(n_250),
.B2(n_272),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_303),
.B(n_254),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_304),
.A2(n_282),
.B1(n_244),
.B2(n_293),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_249),
.B(n_280),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_298),
.B(n_292),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_247),
.C(n_281),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

OA21x2_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_283),
.B(n_275),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_302),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_316),
.C(n_317),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_256),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_301),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_218),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_260),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_321),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_315),
.B1(n_318),
.B2(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_308),
.Y(n_326)
);


endmodule