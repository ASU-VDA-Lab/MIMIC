module real_aes_6446_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g236 ( .A1(n_0), .A2(n_237), .B(n_238), .C(n_242), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_1), .B(n_178), .Y(n_243) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_92), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g459 ( .A(n_2), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_3), .B(n_150), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_4), .A2(n_136), .B(n_141), .C(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_5), .A2(n_131), .B(n_542), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_6), .A2(n_131), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_7), .B(n_178), .Y(n_548) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_8), .A2(n_166), .B(n_182), .Y(n_181) );
AND2x6_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_10), .A2(n_136), .B(n_141), .C(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g486 ( .A(n_11), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_12), .B(n_42), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_13), .B(n_241), .Y(n_506) );
INVx1_ASAP7_75t_L g160 ( .A(n_14), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_15), .B(n_150), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_16), .A2(n_151), .B(n_494), .C(n_496), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_17), .B(n_178), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_18), .A2(n_467), .B1(n_745), .B2(n_751), .C1(n_754), .C2(n_755), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_19), .B(n_215), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_20), .A2(n_141), .B(n_192), .C(n_211), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_21), .A2(n_190), .B(n_240), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_22), .B(n_241), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_23), .B(n_241), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_24), .Y(n_533) );
INVx1_ASAP7_75t_L g525 ( .A(n_25), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_26), .A2(n_141), .B(n_185), .C(n_192), .Y(n_184) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_28), .Y(n_502) );
INVx1_ASAP7_75t_L g582 ( .A(n_29), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_30), .A2(n_104), .B1(n_113), .B2(n_761), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_31), .A2(n_131), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g134 ( .A(n_32), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_33), .A2(n_139), .B(n_154), .C(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_34), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_35), .A2(n_240), .B(n_545), .C(n_547), .Y(n_544) );
INVxp67_ASAP7_75t_L g583 ( .A(n_36), .Y(n_583) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_37), .A2(n_47), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_37), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_38), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_39), .A2(n_141), .B(n_192), .C(n_524), .Y(n_523) );
CKINVDCx14_ASAP7_75t_R g543 ( .A(n_40), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_41), .A2(n_46), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_41), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_43), .A2(n_242), .B(n_484), .C(n_485), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_44), .B(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_45), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_46), .Y(n_749) );
INVx1_ASAP7_75t_L g123 ( .A(n_47), .Y(n_123) );
OAI321xp33_ASAP7_75t_L g119 ( .A1(n_48), .A2(n_120), .A3(n_454), .B1(n_460), .B2(n_461), .C(n_463), .Y(n_119) );
INVx1_ASAP7_75t_L g460 ( .A(n_48), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_49), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_50), .B(n_131), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_51), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_52), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_53), .A2(n_139), .B(n_144), .C(n_154), .Y(n_138) );
INVx1_ASAP7_75t_L g239 ( .A(n_54), .Y(n_239) );
INVx1_ASAP7_75t_L g145 ( .A(n_55), .Y(n_145) );
INVx1_ASAP7_75t_L g514 ( .A(n_56), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_57), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_58), .B(n_131), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_59), .Y(n_218) );
CKINVDCx14_ASAP7_75t_R g482 ( .A(n_60), .Y(n_482) );
INVx1_ASAP7_75t_L g137 ( .A(n_61), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_62), .B(n_131), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_63), .B(n_178), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_64), .A2(n_172), .B(n_174), .C(n_176), .Y(n_171) );
INVx1_ASAP7_75t_L g159 ( .A(n_65), .Y(n_159) );
INVx1_ASAP7_75t_SL g546 ( .A(n_66), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_67), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_68), .B(n_150), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_69), .B(n_178), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_70), .B(n_151), .Y(n_253) );
INVx1_ASAP7_75t_L g536 ( .A(n_71), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_72), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_73), .B(n_147), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_74), .A2(n_141), .B(n_154), .C(n_224), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_75), .Y(n_170) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_77), .A2(n_131), .B(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_78), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_79), .A2(n_131), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_80), .A2(n_209), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g492 ( .A(n_81), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_82), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_83), .B(n_146), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_84), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_84), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_85), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_86), .A2(n_131), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g495 ( .A(n_87), .Y(n_495) );
INVx2_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
INVx1_ASAP7_75t_L g505 ( .A(n_89), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_90), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_91), .B(n_241), .Y(n_254) );
OR2x2_ASAP7_75t_L g456 ( .A(n_92), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g473 ( .A(n_92), .Y(n_473) );
OR2x2_ASAP7_75t_L g744 ( .A(n_92), .B(n_458), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_93), .A2(n_141), .B(n_154), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_94), .B(n_131), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_95), .Y(n_201) );
INVxp67_ASAP7_75t_L g175 ( .A(n_96), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_97), .B(n_166), .Y(n_487) );
INVx2_ASAP7_75t_L g517 ( .A(n_98), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g225 ( .A(n_100), .Y(n_225) );
INVx1_ASAP7_75t_L g249 ( .A(n_101), .Y(n_249) );
AND2x2_ASAP7_75t_L g161 ( .A(n_102), .B(n_156), .Y(n_161) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g761 ( .A(n_106), .Y(n_761) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g458 ( .A(n_107), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_465), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g760 ( .A(n_117), .Y(n_760) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_120), .B(n_462), .Y(n_461) );
XOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_124), .A2(n_469), .B1(n_474), .B2(n_741), .Y(n_468) );
INVx4_ASAP7_75t_L g758 ( .A(n_124), .Y(n_758) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR5x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_327), .C(n_405), .D(n_429), .E(n_446), .Y(n_125) );
OAI211xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_193), .B(n_244), .C(n_304), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
AND2x2_ASAP7_75t_L g258 ( .A(n_128), .B(n_164), .Y(n_258) );
INVx5_ASAP7_75t_SL g286 ( .A(n_128), .Y(n_286) );
AND2x2_ASAP7_75t_L g322 ( .A(n_128), .B(n_307), .Y(n_322) );
OR2x2_ASAP7_75t_L g361 ( .A(n_128), .B(n_163), .Y(n_361) );
OR2x2_ASAP7_75t_L g392 ( .A(n_128), .B(n_283), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_128), .B(n_296), .Y(n_428) );
AND2x2_ASAP7_75t_L g440 ( .A(n_128), .B(n_283), .Y(n_440) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_161), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_138), .B(n_156), .Y(n_129) );
BUFx2_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g250 ( .A(n_132), .B(n_136), .Y(n_250) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
INVx1_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
INVx1_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
INVx1_ASAP7_75t_L g187 ( .A(n_135), .Y(n_187) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_135), .Y(n_241) );
INVx4_ASAP7_75t_SL g155 ( .A(n_136), .Y(n_155) );
BUFx3_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_140), .A2(n_155), .B(n_170), .C(n_171), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_140), .A2(n_155), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_140), .A2(n_155), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_140), .A2(n_155), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_140), .A2(n_155), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_140), .A2(n_155), .B(n_543), .C(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_SL g578 ( .A1(n_140), .A2(n_155), .B(n_579), .C(n_580), .Y(n_578) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_142), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_149), .C(n_152), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_146), .A2(n_152), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_146), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_146), .A2(n_507), .B(n_536), .C(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_150), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g237 ( .A(n_150), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_150), .A2(n_214), .B(n_525), .C(n_526), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_150), .A2(n_173), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_151), .B(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g242 ( .A(n_153), .Y(n_242) );
INVx1_ASAP7_75t_L g496 ( .A(n_153), .Y(n_496) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_156), .A2(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g216 ( .A(n_156), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_156), .Y(n_219) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_156), .A2(n_480), .B(n_487), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_156), .A2(n_250), .B(n_522), .C(n_523), .Y(n_521) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g167 ( .A(n_157), .B(n_158), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g439 ( .A(n_162), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g302 ( .A(n_163), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_164), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_164), .Y(n_295) );
INVx3_ASAP7_75t_L g310 ( .A(n_164), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_164), .B(n_180), .Y(n_334) );
OR2x2_ASAP7_75t_L g343 ( .A(n_164), .B(n_286), .Y(n_343) );
AND2x2_ASAP7_75t_L g347 ( .A(n_164), .B(n_307), .Y(n_347) );
AND2x2_ASAP7_75t_L g353 ( .A(n_164), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g390 ( .A(n_164), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_164), .B(n_247), .Y(n_404) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_177), .Y(n_164) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_165), .A2(n_490), .B(n_497), .Y(n_489) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_165), .A2(n_512), .B(n_518), .Y(n_511) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_165), .A2(n_541), .B(n_548), .Y(n_540) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g179 ( .A(n_166), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_166), .A2(n_183), .B(n_184), .Y(n_182) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g257 ( .A(n_167), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_172), .A2(n_225), .B(n_226), .C(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_173), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_173), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g214 ( .A(n_176), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_176), .B(n_581), .Y(n_580) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_178), .A2(n_233), .B(n_243), .Y(n_232) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_179), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_179), .A2(n_222), .B(n_230), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_179), .B(n_231), .Y(n_230) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_179), .A2(n_248), .B(n_255), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_179), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_179), .B(n_528), .Y(n_527) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_179), .A2(n_532), .B(n_538), .Y(n_531) );
OR2x2_ASAP7_75t_L g296 ( .A(n_180), .B(n_247), .Y(n_296) );
AND2x2_ASAP7_75t_L g307 ( .A(n_180), .B(n_283), .Y(n_307) );
AND2x2_ASAP7_75t_L g319 ( .A(n_180), .B(n_310), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_180), .B(n_247), .Y(n_342) );
INVx1_ASAP7_75t_SL g354 ( .A(n_180), .Y(n_354) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g246 ( .A(n_181), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_181), .B(n_286), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_188), .B(n_189), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_189), .A2(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_205), .Y(n_194) );
AND2x2_ASAP7_75t_L g267 ( .A(n_195), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_195), .B(n_220), .Y(n_271) );
AND2x2_ASAP7_75t_L g274 ( .A(n_195), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_195), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g299 ( .A(n_195), .B(n_290), .Y(n_299) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_195), .Y(n_318) );
AND2x2_ASAP7_75t_L g339 ( .A(n_195), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g349 ( .A(n_195), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g395 ( .A(n_195), .B(n_278), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_195), .B(n_301), .Y(n_422) );
INVx5_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
AND2x2_ASAP7_75t_L g358 ( .A(n_196), .B(n_290), .Y(n_358) );
AND2x2_ASAP7_75t_L g442 ( .A(n_196), .B(n_310), .Y(n_442) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_203), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_205), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_205), .Y(n_431) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_220), .Y(n_205) );
AND2x2_ASAP7_75t_L g261 ( .A(n_206), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g270 ( .A(n_206), .B(n_268), .Y(n_270) );
INVx5_ASAP7_75t_L g278 ( .A(n_206), .Y(n_278) );
AND2x2_ASAP7_75t_L g301 ( .A(n_206), .B(n_232), .Y(n_301) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_206), .Y(n_338) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AOI21xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_210), .B(n_215), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_216), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_219), .A2(n_501), .B(n_508), .Y(n_500) );
INVx1_ASAP7_75t_L g379 ( .A(n_220), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_220), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g412 ( .A(n_220), .B(n_278), .Y(n_412) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_220), .A2(n_335), .B(n_442), .C(n_443), .Y(n_441) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_232), .Y(n_220) );
BUFx2_ASAP7_75t_L g262 ( .A(n_221), .Y(n_262) );
INVx2_ASAP7_75t_L g266 ( .A(n_221), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g547 ( .A(n_228), .Y(n_547) );
INVx2_ASAP7_75t_L g268 ( .A(n_232), .Y(n_268) );
AND2x2_ASAP7_75t_L g275 ( .A(n_232), .B(n_266), .Y(n_275) );
AND2x2_ASAP7_75t_L g366 ( .A(n_232), .B(n_278), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_240), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g484 ( .A(n_241), .Y(n_484) );
INVx2_ASAP7_75t_L g507 ( .A(n_242), .Y(n_507) );
AOI211x1_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_259), .B(n_272), .C(n_297), .Y(n_244) );
INVx1_ASAP7_75t_L g363 ( .A(n_245), .Y(n_363) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_258), .Y(n_245) );
INVx5_ASAP7_75t_SL g283 ( .A(n_247), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_247), .B(n_353), .Y(n_352) );
AOI311xp33_ASAP7_75t_L g371 ( .A1(n_247), .A2(n_372), .A3(n_374), .B(n_375), .C(n_381), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_247), .A2(n_319), .B(n_407), .C(n_410), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_251), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_250), .A2(n_502), .B(n_503), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_250), .A2(n_533), .B(n_534), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g575 ( .A(n_257), .Y(n_575) );
INVxp67_ASAP7_75t_L g326 ( .A(n_258), .Y(n_326) );
NAND4xp25_ASAP7_75t_SL g259 ( .A(n_260), .B(n_263), .C(n_269), .D(n_271), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_260), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g317 ( .A(n_261), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_264), .B(n_270), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_264), .B(n_277), .Y(n_397) );
BUFx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_265), .B(n_278), .Y(n_415) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
INVxp67_ASAP7_75t_L g325 ( .A(n_267), .Y(n_325) );
AND2x4_ASAP7_75t_L g277 ( .A(n_268), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g351 ( .A(n_268), .B(n_290), .Y(n_351) );
INVx1_ASAP7_75t_L g378 ( .A(n_268), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_268), .B(n_365), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_269), .B(n_339), .Y(n_359) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_270), .B(n_292), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_270), .B(n_339), .Y(n_438) );
INVx1_ASAP7_75t_L g449 ( .A(n_271), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B(n_279), .C(n_287), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g291 ( .A(n_275), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_275), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g311 ( .A(n_276), .Y(n_311) );
AND2x2_ASAP7_75t_L g288 ( .A(n_277), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_277), .B(n_339), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_277), .B(n_358), .Y(n_382) );
OR2x2_ASAP7_75t_L g298 ( .A(n_278), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g330 ( .A(n_278), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_278), .B(n_290), .Y(n_345) );
AND2x2_ASAP7_75t_L g402 ( .A(n_278), .B(n_358), .Y(n_402) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_278), .Y(n_409) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_280), .A2(n_292), .B1(n_414), .B2(n_416), .C(n_419), .Y(n_413) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_286), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_283), .B(n_353), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_283), .B(n_310), .Y(n_418) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g403 ( .A(n_285), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g417 ( .A(n_285), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_286), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_307), .Y(n_314) );
AND2x2_ASAP7_75t_L g384 ( .A(n_286), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_286), .B(n_333), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_286), .B(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_291), .B(n_293), .Y(n_287) );
INVx2_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g340 ( .A(n_290), .Y(n_340) );
OR2x2_ASAP7_75t_L g344 ( .A(n_292), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g447 ( .A(n_292), .B(n_415), .Y(n_447) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AOI21xp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_300), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_L g451 ( .A(n_298), .Y(n_451) );
INVx2_ASAP7_75t_SL g365 ( .A(n_299), .Y(n_365) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_302), .A2(n_383), .B(n_447), .C(n_448), .Y(n_446) );
OAI322xp33_ASAP7_75t_SL g315 ( .A1(n_303), .A2(n_316), .A3(n_319), .B1(n_320), .B2(n_321), .C1(n_323), .C2(n_326), .Y(n_315) );
INVx2_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_311), .B1(n_312), .B2(n_314), .C(n_315), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp33_ASAP7_75t_SL g381 ( .A1(n_306), .A2(n_382), .B1(n_383), .B2(n_386), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_307), .B(n_310), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_307), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g380 ( .A(n_309), .B(n_342), .Y(n_380) );
INVx1_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_314), .A2(n_424), .B(n_426), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_316), .A2(n_349), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp67_ASAP7_75t_SL g377 ( .A(n_318), .B(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_318), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g434 ( .A(n_319), .Y(n_434) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_328), .B(n_355), .C(n_371), .D(n_387), .Y(n_327) );
AOI211xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B(n_336), .C(n_348), .Y(n_328) );
INVx1_ASAP7_75t_L g420 ( .A(n_329), .Y(n_420) );
AND2x2_ASAP7_75t_L g368 ( .A(n_330), .B(n_351), .Y(n_368) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_335), .B(n_370), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B1(n_344), .B2(n_346), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_338), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_339), .A2(n_378), .B(n_401), .C(n_403), .Y(n_400) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
INVx1_ASAP7_75t_L g445 ( .A(n_343), .Y(n_445) );
NAND2xp33_ASAP7_75t_SL g435 ( .A(n_344), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B(n_360), .C(n_362), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_367), .B2(n_369), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_365), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_370), .B(n_391), .Y(n_453) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_379), .B(n_380), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B1(n_396), .B2(n_398), .C(n_400), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_403), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
NAND3xp33_ASAP7_75t_SL g405 ( .A(n_406), .B(n_413), .C(n_423), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_432), .C(n_441), .Y(n_429) );
INVx1_ASAP7_75t_L g450 ( .A(n_430), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B1(n_437), .B2(n_439), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_451), .B2(n_452), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g462 ( .A(n_456), .Y(n_462) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_457), .B(n_473), .Y(n_753) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g472 ( .A(n_458), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g464 ( .A(n_462), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_463), .B(n_466), .C(n_759), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI22x1_ASAP7_75t_SL g756 ( .A1(n_469), .A2(n_741), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g757 ( .A(n_474), .Y(n_757) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_671), .Y(n_474) );
NAND5xp2_ASAP7_75t_L g475 ( .A(n_476), .B(n_586), .C(n_618), .D(n_635), .E(n_658), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_519), .B1(n_549), .B2(n_553), .C(n_557), .Y(n_476) );
INVx1_ASAP7_75t_L g698 ( .A(n_477), .Y(n_698) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_498), .Y(n_477) );
AND3x2_ASAP7_75t_L g673 ( .A(n_478), .B(n_500), .C(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_479), .B(n_555), .Y(n_554) );
BUFx3_ASAP7_75t_L g564 ( .A(n_479), .Y(n_564) );
AND2x2_ASAP7_75t_L g568 ( .A(n_479), .B(n_510), .Y(n_568) );
INVx2_ASAP7_75t_L g595 ( .A(n_479), .Y(n_595) );
OR2x2_ASAP7_75t_L g606 ( .A(n_479), .B(n_511), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_479), .B(n_499), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_479), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g685 ( .A(n_479), .B(n_511), .Y(n_685) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_488), .Y(n_567) );
AND2x2_ASAP7_75t_L g626 ( .A(n_488), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_488), .B(n_499), .Y(n_645) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g556 ( .A(n_489), .B(n_499), .Y(n_556) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
AND2x2_ASAP7_75t_L g612 ( .A(n_489), .B(n_511), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_489), .B(n_498), .C(n_595), .Y(n_637) );
AND2x2_ASAP7_75t_L g702 ( .A(n_489), .B(n_500), .Y(n_702) );
AND2x2_ASAP7_75t_L g736 ( .A(n_489), .B(n_499), .Y(n_736) );
INVxp67_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_499), .B(n_595), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_499), .B(n_626), .Y(n_634) );
AND2x2_ASAP7_75t_L g684 ( .A(n_499), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g712 ( .A(n_499), .Y(n_712) );
INVx4_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g619 ( .A(n_500), .B(n_612), .Y(n_619) );
BUFx3_ASAP7_75t_L g651 ( .A(n_500), .Y(n_651) );
INVx2_ASAP7_75t_L g627 ( .A(n_510), .Y(n_627) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_511), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_519), .A2(n_687), .B1(n_689), .B2(n_690), .Y(n_686) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
AND2x2_ASAP7_75t_L g549 ( .A(n_520), .B(n_550), .Y(n_549) );
INVx3_ASAP7_75t_SL g560 ( .A(n_520), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_520), .B(n_590), .Y(n_622) );
OR2x2_ASAP7_75t_L g641 ( .A(n_520), .B(n_530), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_520), .B(n_598), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_520), .B(n_591), .Y(n_649) );
AND2x2_ASAP7_75t_L g661 ( .A(n_520), .B(n_540), .Y(n_661) );
AND2x2_ASAP7_75t_L g677 ( .A(n_520), .B(n_531), .Y(n_677) );
AND2x4_ASAP7_75t_L g680 ( .A(n_520), .B(n_551), .Y(n_680) );
OR2x2_ASAP7_75t_L g697 ( .A(n_520), .B(n_633), .Y(n_697) );
OR2x2_ASAP7_75t_L g728 ( .A(n_520), .B(n_573), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_520), .B(n_656), .Y(n_730) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .Y(n_520) );
AND2x2_ASAP7_75t_L g604 ( .A(n_529), .B(n_571), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_529), .B(n_591), .Y(n_723) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
AND2x2_ASAP7_75t_L g559 ( .A(n_530), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g590 ( .A(n_530), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_530), .B(n_573), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_530), .B(n_551), .Y(n_616) );
OR2x2_ASAP7_75t_L g633 ( .A(n_530), .B(n_591), .Y(n_633) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
AND2x2_ASAP7_75t_L g656 ( .A(n_531), .B(n_540), .Y(n_656) );
INVx2_ASAP7_75t_L g551 ( .A(n_540), .Y(n_551) );
INVx1_ASAP7_75t_L g668 ( .A(n_540), .Y(n_668) );
AND2x2_ASAP7_75t_L g718 ( .A(n_540), .B(n_560), .Y(n_718) );
AND2x2_ASAP7_75t_L g570 ( .A(n_550), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g602 ( .A(n_550), .B(n_560), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_550), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g589 ( .A(n_551), .B(n_560), .Y(n_589) );
OR2x2_ASAP7_75t_L g705 ( .A(n_552), .B(n_679), .Y(n_705) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_555), .B(n_685), .Y(n_691) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g647 ( .A1(n_556), .A2(n_648), .A3(n_650), .B1(n_652), .B2(n_653), .Y(n_647) );
OR2x2_ASAP7_75t_L g664 ( .A(n_556), .B(n_606), .Y(n_664) );
OAI21xp33_ASAP7_75t_SL g689 ( .A1(n_556), .A2(n_566), .B(n_594), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_566), .B2(n_569), .Y(n_557) );
INVxp33_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_559), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_560), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g615 ( .A(n_560), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g715 ( .A(n_560), .B(n_656), .Y(n_715) );
OR2x2_ASAP7_75t_L g739 ( .A(n_560), .B(n_633), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_561), .A2(n_621), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g599 ( .A(n_563), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_563), .B(n_568), .Y(n_617) );
AND2x2_ASAP7_75t_L g639 ( .A(n_564), .B(n_612), .Y(n_639) );
INVx1_ASAP7_75t_L g652 ( .A(n_564), .Y(n_652) );
OR2x2_ASAP7_75t_L g657 ( .A(n_564), .B(n_591), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_567), .B(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_568), .A2(n_588), .B1(n_593), .B2(n_597), .Y(n_587) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_571), .A2(n_630), .B1(n_637), .B2(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g714 ( .A(n_571), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_573), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g733 ( .A(n_573), .B(n_616), .Y(n_733) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_584), .Y(n_573) );
INVx1_ASAP7_75t_L g592 ( .A(n_574), .Y(n_592) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_577), .A2(n_585), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_599), .B1(n_600), .B2(n_605), .C(n_607), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_589), .B(n_591), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_589), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g608 ( .A(n_590), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g695 ( .A1(n_590), .A2(n_696), .B(n_697), .C(n_698), .Y(n_695) );
AND2x2_ASAP7_75t_L g700 ( .A(n_590), .B(n_680), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_SL g738 ( .A1(n_590), .A2(n_679), .B(n_739), .C(n_740), .Y(n_738) );
BUFx3_ASAP7_75t_L g630 ( .A(n_591), .Y(n_630) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_594), .B(n_651), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_594), .A2(n_714), .B(n_716), .C(n_722), .Y(n_713) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVxp67_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_598), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_602), .A2(n_619), .B(n_620), .C(n_628), .Y(n_618) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g703 ( .A(n_606), .Y(n_703) );
OR2x2_ASAP7_75t_L g720 ( .A(n_606), .B(n_650), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_614), .B2(n_617), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_609), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
OR2x2_ASAP7_75t_L g707 ( .A(n_611), .B(n_651), .Y(n_707) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g662 ( .A(n_612), .B(n_652), .Y(n_662) );
INVx1_ASAP7_75t_L g670 ( .A(n_613), .Y(n_670) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_616), .B(n_630), .Y(n_678) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_626), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g735 ( .A(n_627), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_634), .Y(n_628) );
INVx1_ASAP7_75t_L g665 ( .A(n_629), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_630), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_630), .B(n_661), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g681 ( .A(n_630), .B(n_656), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_630), .B(n_677), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_630), .A2(n_640), .B(n_680), .C(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_640), .B1(n_642), .B2(n_646), .C(n_647), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_644), .B(n_652), .Y(n_726) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_646), .A2(n_661), .B(n_663), .C(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_649), .B(n_656), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_650), .B(n_703), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g650 ( .A(n_651), .Y(n_650) );
INVxp33_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
AOI21xp33_ASAP7_75t_SL g666 ( .A1(n_655), .A2(n_667), .B(n_669), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_655), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_656), .B(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B1(n_663), .B2(n_665), .C(n_666), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_662), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g696 ( .A(n_668), .Y(n_696) );
NAND5xp2_ASAP7_75t_L g671 ( .A(n_672), .B(n_699), .C(n_713), .D(n_724), .E(n_737), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_682), .C(n_695), .Y(n_672) );
INVx2_ASAP7_75t_SL g719 ( .A(n_673), .Y(n_719) );
NAND4xp25_ASAP7_75t_SL g675 ( .A(n_676), .B(n_678), .C(n_679), .D(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_681), .A2(n_683), .B(n_686), .C(n_692), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_684), .A2(n_725), .B1(n_727), .B2(n_729), .C(n_731), .Y(n_724) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI221xp5_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_701), .B1(n_704), .B2(n_706), .C(n_708), .Y(n_699) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_707), .A2(n_730), .B1(n_732), .B2(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_745), .Y(n_754) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
endmodule