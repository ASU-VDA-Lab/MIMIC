module real_aes_6943_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g271 ( .A1(n_0), .A2(n_272), .B(n_273), .C(n_276), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_1), .B(n_213), .Y(n_277) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_3), .B(n_183), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_4), .A2(n_153), .B(n_156), .C(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_5), .A2(n_173), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_6), .A2(n_173), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_7), .B(n_213), .Y(n_527) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_8), .A2(n_140), .B(n_193), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_9), .A2(n_743), .B1(n_746), .B2(n_747), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_9), .Y(n_747) );
AND2x6_ASAP7_75t_L g153 ( .A(n_10), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_11), .A2(n_153), .B(n_156), .C(n_159), .Y(n_155) );
INVx1_ASAP7_75t_L g497 ( .A(n_12), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_13), .B(n_42), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_13), .B(n_42), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_14), .A2(n_46), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_14), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_15), .B(n_163), .Y(n_483) );
INVx1_ASAP7_75t_L g145 ( .A(n_16), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_17), .B(n_183), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_18), .A2(n_161), .B(n_505), .C(n_507), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_19), .B(n_213), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_20), .A2(n_105), .B1(n_118), .B2(n_756), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_21), .B(n_237), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_22), .A2(n_156), .B(n_200), .C(n_233), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_23), .A2(n_165), .B(n_275), .C(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_24), .B(n_163), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_25), .B(n_163), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_26), .Y(n_555) );
INVx1_ASAP7_75t_L g547 ( .A(n_27), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_28), .A2(n_156), .B(n_196), .C(n_200), .Y(n_195) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_29), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_30), .Y(n_479) );
INVx1_ASAP7_75t_L g538 ( .A(n_31), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_32), .A2(n_173), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g151 ( .A(n_33), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_34), .A2(n_175), .B(n_186), .C(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_35), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_36), .A2(n_275), .B(n_524), .C(n_526), .Y(n_523) );
INVxp67_ASAP7_75t_L g539 ( .A(n_37), .Y(n_539) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_38), .A2(n_79), .B1(n_454), .B2(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_38), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_39), .B(n_198), .Y(n_197) );
CKINVDCx14_ASAP7_75t_R g522 ( .A(n_40), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_41), .A2(n_156), .B(n_200), .C(n_546), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_43), .A2(n_276), .B(n_495), .C(n_496), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_44), .B(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_45), .Y(n_168) );
INVx1_ASAP7_75t_L g745 ( .A(n_46), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_47), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_48), .B(n_173), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_49), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_50), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_51), .A2(n_175), .B(n_177), .C(n_186), .Y(n_174) );
INVx1_ASAP7_75t_L g274 ( .A(n_52), .Y(n_274) );
INVx1_ASAP7_75t_L g178 ( .A(n_53), .Y(n_178) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_54), .A2(n_465), .B1(n_738), .B2(n_739), .C1(n_748), .C2(n_751), .Y(n_464) );
INVx1_ASAP7_75t_L g512 ( .A(n_55), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_56), .B(n_173), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_57), .A2(n_60), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_57), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_58), .Y(n_240) );
CKINVDCx14_ASAP7_75t_R g493 ( .A(n_59), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_60), .Y(n_128) );
INVx1_ASAP7_75t_L g154 ( .A(n_61), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_62), .B(n_173), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_63), .B(n_213), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_64), .A2(n_207), .B(n_209), .C(n_211), .Y(n_206) );
INVx1_ASAP7_75t_L g144 ( .A(n_65), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_66), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g525 ( .A(n_67), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_68), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_69), .B(n_183), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_70), .B(n_213), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_71), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g558 ( .A(n_72), .Y(n_558) );
CKINVDCx16_ASAP7_75t_R g270 ( .A(n_73), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_74), .B(n_180), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_75), .A2(n_156), .B(n_186), .C(n_247), .Y(n_246) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_76), .Y(n_205) );
INVx1_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_78), .A2(n_173), .B(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_79), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_80), .A2(n_173), .B(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_81), .A2(n_231), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g503 ( .A(n_82), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_83), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_84), .B(n_179), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_85), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_86), .A2(n_173), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g506 ( .A(n_87), .Y(n_506) );
INVx2_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
INVx1_ASAP7_75t_L g482 ( .A(n_89), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_90), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_91), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
OR2x2_ASAP7_75t_L g449 ( .A(n_92), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g468 ( .A(n_92), .B(n_451), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_93), .A2(n_156), .B(n_186), .C(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_94), .B(n_173), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_95), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_95), .Y(n_740) );
INVx1_ASAP7_75t_L g222 ( .A(n_96), .Y(n_222) );
INVxp67_ASAP7_75t_L g210 ( .A(n_97), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_98), .B(n_140), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_99), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g147 ( .A(n_100), .Y(n_147) );
INVx1_ASAP7_75t_L g248 ( .A(n_101), .Y(n_248) );
INVx2_ASAP7_75t_L g515 ( .A(n_102), .Y(n_515) );
AND2x2_ASAP7_75t_L g189 ( .A(n_103), .B(n_188), .Y(n_189) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g756 ( .A(n_107), .Y(n_756) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g451 ( .A(n_113), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g737 ( .A(n_114), .B(n_451), .Y(n_737) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_114), .B(n_450), .Y(n_753) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_463), .Y(n_118) );
BUFx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g755 ( .A(n_122), .Y(n_755) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI321xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_447), .A3(n_453), .B1(n_456), .B2(n_457), .C(n_460), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_125), .B(n_458), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_SL g465 ( .A1(n_130), .A2(n_466), .B1(n_469), .B2(n_735), .Y(n_465) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_131), .A2(n_470), .B1(n_749), .B2(n_750), .Y(n_748) );
OR3x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_345), .C(n_410), .Y(n_131) );
NAND4xp25_ASAP7_75t_SL g132 ( .A(n_133), .B(n_286), .C(n_312), .D(n_335), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_214), .B1(n_255), .B2(n_262), .C(n_278), .Y(n_133) );
CKINVDCx14_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_135), .A2(n_279), .B1(n_303), .B2(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_190), .Y(n_135) );
INVx1_ASAP7_75t_SL g339 ( .A(n_136), .Y(n_339) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_170), .Y(n_136) );
OR2x2_ASAP7_75t_L g260 ( .A(n_137), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g281 ( .A(n_137), .B(n_191), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_137), .B(n_201), .Y(n_294) );
AND2x2_ASAP7_75t_L g311 ( .A(n_137), .B(n_170), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_137), .B(n_258), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_137), .B(n_310), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_137), .B(n_190), .Y(n_432) );
AOI211xp5_ASAP7_75t_SL g443 ( .A1(n_137), .A2(n_349), .B(n_444), .C(n_445), .Y(n_443) );
INVx5_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_138), .B(n_191), .Y(n_315) );
AND2x2_ASAP7_75t_L g318 ( .A(n_138), .B(n_192), .Y(n_318) );
OR2x2_ASAP7_75t_L g363 ( .A(n_138), .B(n_191), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_138), .B(n_201), .Y(n_372) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_167), .Y(n_138) );
INVx3_ASAP7_75t_L g213 ( .A(n_139), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_139), .B(n_225), .Y(n_224) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_139), .A2(n_245), .B(n_253), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_139), .B(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_139), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_139), .B(n_550), .Y(n_549) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_139), .A2(n_554), .B(n_560), .Y(n_553) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_140), .A2(n_194), .B(n_195), .Y(n_193) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g188 ( .A(n_142), .B(n_143), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_155), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_148), .A2(n_479), .B(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_148), .A2(n_188), .B(n_544), .C(n_545), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_148), .A2(n_555), .B(n_556), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
AND2x4_ASAP7_75t_L g173 ( .A(n_149), .B(n_153), .Y(n_173) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx1_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx3_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx1_ASAP7_75t_L g198 ( .A(n_152), .Y(n_198) );
INVx4_ASAP7_75t_SL g187 ( .A(n_153), .Y(n_187) );
BUFx3_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVx5_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_157), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_164), .Y(n_159) );
INVx5_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_161), .B(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g275 ( .A(n_163), .Y(n_275) );
INVx2_ASAP7_75t_L g495 ( .A(n_163), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_164), .A2(n_197), .B(n_199), .Y(n_196) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx2_ASAP7_75t_L g532 ( .A(n_169), .Y(n_532) );
INVx5_ASAP7_75t_SL g261 ( .A(n_170), .Y(n_261) );
AND2x2_ASAP7_75t_L g280 ( .A(n_170), .B(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_170), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g366 ( .A(n_170), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g398 ( .A(n_170), .B(n_201), .Y(n_398) );
OR2x2_ASAP7_75t_L g404 ( .A(n_170), .B(n_294), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_170), .B(n_354), .Y(n_413) );
OR2x6_ASAP7_75t_L g170 ( .A(n_171), .B(n_189), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_188), .Y(n_171) );
BUFx2_ASAP7_75t_L g231 ( .A(n_173), .Y(n_231) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_176), .A2(n_187), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_176), .A2(n_187), .B(n_270), .C(n_271), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_176), .A2(n_187), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_176), .A2(n_187), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_176), .A2(n_187), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_176), .A2(n_187), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_176), .A2(n_187), .B(n_535), .C(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_182), .C(n_184), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_179), .A2(n_184), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp5_ASAP7_75t_L g481 ( .A1(n_179), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_179), .A2(n_484), .B(n_558), .C(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g208 ( .A(n_181), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_183), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g272 ( .A(n_183), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_183), .A2(n_208), .B1(n_538), .B2(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_183), .A2(n_236), .B(n_547), .C(n_548), .Y(n_546) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g276 ( .A(n_185), .Y(n_276) );
INVx1_ASAP7_75t_L g507 ( .A(n_185), .Y(n_507) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_188), .A2(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
INVx1_ASAP7_75t_L g241 ( .A(n_188), .Y(n_241) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_188), .A2(n_491), .B(n_498), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
AND2x2_ASAP7_75t_L g295 ( .A(n_191), .B(n_261), .Y(n_295) );
INVx1_ASAP7_75t_SL g308 ( .A(n_191), .Y(n_308) );
OR2x2_ASAP7_75t_L g343 ( .A(n_191), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g349 ( .A(n_191), .B(n_201), .Y(n_349) );
AND2x2_ASAP7_75t_L g407 ( .A(n_191), .B(n_258), .Y(n_407) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_192), .B(n_261), .Y(n_334) );
INVx3_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
OR2x2_ASAP7_75t_L g300 ( .A(n_201), .B(n_261), .Y(n_300) );
AND2x2_ASAP7_75t_L g310 ( .A(n_201), .B(n_308), .Y(n_310) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_201), .Y(n_358) );
AND2x2_ASAP7_75t_L g367 ( .A(n_201), .B(n_281), .Y(n_367) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_201) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_202), .A2(n_501), .B(n_508), .Y(n_500) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_202), .A2(n_510), .B(n_516), .Y(n_509) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_202), .A2(n_520), .B(n_527), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_207), .A2(n_248), .B(n_249), .C(n_250), .Y(n_247) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_208), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_208), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g236 ( .A(n_211), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_211), .B(n_537), .Y(n_536) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_213), .A2(n_268), .B(n_277), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_214), .A2(n_384), .B1(n_386), .B2(n_388), .C(n_391), .Y(n_383) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
AND2x2_ASAP7_75t_L g357 ( .A(n_216), .B(n_338), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_216), .B(n_416), .Y(n_420) );
OR2x2_ASAP7_75t_L g441 ( .A(n_216), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_216), .B(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx5_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
AND2x2_ASAP7_75t_L g365 ( .A(n_217), .B(n_228), .Y(n_365) );
AND2x2_ASAP7_75t_L g426 ( .A(n_217), .B(n_305), .Y(n_426) );
AND2x2_ASAP7_75t_L g439 ( .A(n_217), .B(n_258), .Y(n_439) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_242), .Y(n_226) );
AND2x4_ASAP7_75t_L g265 ( .A(n_227), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g284 ( .A(n_227), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
AND2x2_ASAP7_75t_L g360 ( .A(n_227), .B(n_338), .Y(n_360) );
AND2x2_ASAP7_75t_L g370 ( .A(n_227), .B(n_288), .Y(n_370) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_227), .Y(n_378) );
AND2x2_ASAP7_75t_L g390 ( .A(n_227), .B(n_267), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_227), .B(n_322), .Y(n_394) );
AND2x2_ASAP7_75t_L g431 ( .A(n_227), .B(n_426), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_227), .B(n_305), .Y(n_442) );
OR2x2_ASAP7_75t_L g444 ( .A(n_227), .B(n_380), .Y(n_444) );
INVx5_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g330 ( .A(n_228), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g340 ( .A(n_228), .B(n_285), .Y(n_340) );
AND2x2_ASAP7_75t_L g352 ( .A(n_228), .B(n_267), .Y(n_352) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_228), .Y(n_382) );
AND2x4_ASAP7_75t_L g416 ( .A(n_228), .B(n_266), .Y(n_416) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_239), .Y(n_228) );
AOI21xp5_ASAP7_75t_SL g229 ( .A1(n_230), .A2(n_232), .B(n_237), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .Y(n_233) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_238), .B(n_455), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_241), .A2(n_478), .B(n_485), .Y(n_477) );
BUFx2_ASAP7_75t_L g264 ( .A(n_242), .Y(n_264) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g305 ( .A(n_243), .Y(n_305) );
AND2x2_ASAP7_75t_L g338 ( .A(n_243), .B(n_267), .Y(n_338) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g285 ( .A(n_244), .B(n_267), .Y(n_285) );
BUFx2_ASAP7_75t_L g331 ( .A(n_244), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_252), .Y(n_245) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g526 ( .A(n_251), .Y(n_526) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_257), .B(n_339), .Y(n_418) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_258), .B(n_281), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_258), .B(n_261), .Y(n_320) );
AND2x2_ASAP7_75t_L g375 ( .A(n_258), .B(n_311), .Y(n_375) );
AOI221xp5_ASAP7_75t_SL g312 ( .A1(n_259), .A2(n_313), .B1(n_321), .B2(n_323), .C(n_327), .Y(n_312) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g307 ( .A(n_260), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g348 ( .A(n_260), .B(n_349), .Y(n_348) );
OAI321xp33_ASAP7_75t_L g355 ( .A1(n_260), .A2(n_314), .A3(n_356), .B1(n_358), .B2(n_359), .C(n_361), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_261), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_264), .B(n_416), .Y(n_434) );
AND2x2_ASAP7_75t_L g321 ( .A(n_265), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_265), .B(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
AND2x2_ASAP7_75t_L g304 ( .A(n_266), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_266), .B(n_379), .Y(n_409) );
INVx1_ASAP7_75t_L g446 ( .A(n_266), .Y(n_446) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_275), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g484 ( .A(n_276), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B(n_283), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_280), .A2(n_390), .B(n_439), .C(n_440), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_281), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_281), .B(n_319), .Y(n_385) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_285), .B(n_288), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_285), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_285), .B(n_370), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B1(n_301), .B2(n_306), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g302 ( .A(n_288), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g337 ( .A(n_288), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_288), .B(n_331), .Y(n_373) );
OR2x2_ASAP7_75t_L g380 ( .A(n_288), .B(n_305), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_288), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g430 ( .A(n_288), .B(n_416), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .B1(n_296), .B2(n_298), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g336 ( .A(n_291), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_294), .A2(n_309), .B1(n_377), .B2(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g424 ( .A(n_295), .Y(n_424) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_299), .A2(n_336), .B1(n_339), .B2(n_340), .C(n_341), .Y(n_335) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g314 ( .A(n_300), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_304), .B(n_370), .Y(n_402) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_305), .Y(n_322) );
INVx1_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
NAND2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_311), .B(n_354), .Y(n_353) );
NAND2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g397 ( .A(n_318), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_321), .A2(n_347), .B1(n_350), .B2(n_353), .C(n_355), .Y(n_346) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_325), .B(n_382), .Y(n_381) );
AOI21xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_329), .B(n_332), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_332), .Y(n_429) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OR2x2_ASAP7_75t_L g371 ( .A(n_334), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g392 ( .A(n_337), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_337), .B(n_397), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_340), .B(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g345 ( .A(n_346), .B(n_364), .C(n_383), .D(n_396), .Y(n_345) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g354 ( .A(n_349), .Y(n_354) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_363), .Y(n_387) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_368), .C(n_376), .Y(n_364) );
AOI211xp5_ASAP7_75t_L g435 ( .A1(n_366), .A2(n_408), .B(n_436), .C(n_443), .Y(n_435) );
INVx1_ASAP7_75t_SL g395 ( .A(n_367), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B1(n_373), .B2(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g399 ( .A(n_373), .Y(n_399) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_379), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_379), .B(n_390), .Y(n_423) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g400 ( .A(n_390), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_395), .Y(n_391) );
INVxp33_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI322xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .A3(n_400), .B1(n_401), .B2(n_403), .C1(n_405), .C2(n_408), .Y(n_396) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_411), .B(n_428), .C(n_435), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_417), .B2(n_419), .C(n_421), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g427 ( .A(n_416), .Y(n_427) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_431), .B2(n_432), .C(n_433), .Y(n_428) );
NAND2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g459 ( .A(n_449), .Y(n_459) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_449), .Y(n_462) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g456 ( .A(n_453), .Y(n_456) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_460), .B(n_464), .C(n_754), .Y(n_463) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g749 ( .A(n_467), .Y(n_749) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_690), .Y(n_470) );
NAND5xp2_ASAP7_75t_L g471 ( .A(n_472), .B(n_602), .C(n_640), .D(n_661), .E(n_678), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_574), .C(n_595), .Y(n_472) );
OAI221xp5_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_517), .B1(n_541), .B2(n_561), .C(n_565), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_487), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_476), .B(n_563), .Y(n_582) );
OR2x2_ASAP7_75t_L g609 ( .A(n_476), .B(n_500), .Y(n_609) );
AND2x2_ASAP7_75t_L g623 ( .A(n_476), .B(n_500), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_476), .B(n_490), .Y(n_637) );
AND2x2_ASAP7_75t_L g675 ( .A(n_476), .B(n_639), .Y(n_675) );
AND2x2_ASAP7_75t_L g704 ( .A(n_476), .B(n_614), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_476), .B(n_586), .Y(n_721) );
INVx4_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g601 ( .A(n_477), .B(n_499), .Y(n_601) );
BUFx3_ASAP7_75t_L g626 ( .A(n_477), .Y(n_626) );
AND2x2_ASAP7_75t_L g655 ( .A(n_477), .B(n_500), .Y(n_655) );
AND3x2_ASAP7_75t_L g668 ( .A(n_477), .B(n_669), .C(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g591 ( .A(n_487), .Y(n_591) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_499), .Y(n_487) );
AOI32xp33_ASAP7_75t_L g646 ( .A1(n_488), .A2(n_598), .A3(n_647), .B1(n_650), .B2(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g573 ( .A(n_489), .B(n_499), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_489), .B(n_601), .Y(n_644) );
AND2x2_ASAP7_75t_L g651 ( .A(n_489), .B(n_623), .Y(n_651) );
OR2x2_ASAP7_75t_L g657 ( .A(n_489), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_489), .B(n_612), .Y(n_682) );
OR2x2_ASAP7_75t_L g700 ( .A(n_489), .B(n_529), .Y(n_700) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g564 ( .A(n_490), .B(n_509), .Y(n_564) );
INVx2_ASAP7_75t_L g586 ( .A(n_490), .Y(n_586) );
OR2x2_ASAP7_75t_L g608 ( .A(n_490), .B(n_509), .Y(n_608) );
AND2x2_ASAP7_75t_L g613 ( .A(n_490), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_490), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g669 ( .A(n_490), .B(n_563), .Y(n_669) );
INVx1_ASAP7_75t_SL g720 ( .A(n_499), .Y(n_720) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
INVx1_ASAP7_75t_SL g563 ( .A(n_500), .Y(n_563) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_500), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_500), .B(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_500), .B(n_586), .C(n_704), .Y(n_715) );
INVx2_ASAP7_75t_L g614 ( .A(n_509), .Y(n_614) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_509), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx1_ASAP7_75t_L g650 ( .A(n_518), .Y(n_650) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g568 ( .A(n_519), .B(n_552), .Y(n_568) );
INVx2_ASAP7_75t_L g585 ( .A(n_519), .Y(n_585) );
AND2x2_ASAP7_75t_L g590 ( .A(n_519), .B(n_553), .Y(n_590) );
AND2x2_ASAP7_75t_L g605 ( .A(n_519), .B(n_542), .Y(n_605) );
AND2x2_ASAP7_75t_L g617 ( .A(n_519), .B(n_589), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_528), .B(n_633), .Y(n_632) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_528), .B(n_590), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_528), .B(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_528), .B(n_584), .Y(n_712) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g551 ( .A(n_529), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_529), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g594 ( .A(n_529), .B(n_542), .Y(n_594) );
AND2x2_ASAP7_75t_L g620 ( .A(n_529), .B(n_552), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_529), .B(n_660), .Y(n_659) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_533), .B(n_540), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_531), .A2(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g579 ( .A(n_533), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_540), .Y(n_580) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_551), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_542), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g584 ( .A(n_542), .B(n_585), .Y(n_584) );
INVx3_ASAP7_75t_SL g589 ( .A(n_542), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_542), .B(n_576), .Y(n_642) );
OR2x2_ASAP7_75t_L g652 ( .A(n_542), .B(n_578), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_542), .B(n_620), .Y(n_680) );
OR2x2_ASAP7_75t_L g710 ( .A(n_542), .B(n_552), .Y(n_710) );
AND2x2_ASAP7_75t_L g714 ( .A(n_542), .B(n_553), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_542), .B(n_590), .Y(n_727) );
AND2x2_ASAP7_75t_L g734 ( .A(n_542), .B(n_616), .Y(n_734) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_549), .Y(n_542) );
INVx1_ASAP7_75t_SL g677 ( .A(n_551), .Y(n_677) );
AND2x2_ASAP7_75t_L g616 ( .A(n_552), .B(n_578), .Y(n_616) );
AND2x2_ASAP7_75t_L g630 ( .A(n_552), .B(n_585), .Y(n_630) );
AND2x2_ASAP7_75t_L g633 ( .A(n_552), .B(n_589), .Y(n_633) );
INVx1_ASAP7_75t_L g660 ( .A(n_552), .Y(n_660) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g572 ( .A(n_553), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_562), .A2(n_608), .B(n_732), .C(n_733), .Y(n_731) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g638 ( .A(n_563), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_564), .B(n_581), .Y(n_596) );
AND2x2_ASAP7_75t_L g622 ( .A(n_564), .B(n_623), .Y(n_622) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_569), .B(n_573), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_567), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g593 ( .A(n_568), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_568), .B(n_589), .Y(n_634) );
AND2x2_ASAP7_75t_L g725 ( .A(n_568), .B(n_576), .Y(n_725) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g598 ( .A(n_572), .B(n_585), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_572), .B(n_583), .Y(n_599) );
OAI322xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_582), .A3(n_583), .B1(n_586), .B2(n_587), .C1(n_591), .C2(n_592), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_581), .Y(n_575) );
AND2x2_ASAP7_75t_L g686 ( .A(n_576), .B(n_598), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_576), .B(n_650), .Y(n_732) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g629 ( .A(n_578), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g695 ( .A(n_582), .B(n_608), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_583), .B(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_584), .B(n_616), .Y(n_673) );
AND2x2_ASAP7_75t_L g619 ( .A(n_585), .B(n_589), .Y(n_619) );
AND2x2_ASAP7_75t_L g627 ( .A(n_586), .B(n_628), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_586), .A2(n_665), .B(n_725), .C(n_726), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_587), .A2(n_600), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_589), .B(n_616), .Y(n_656) );
AND2x2_ASAP7_75t_L g662 ( .A(n_589), .B(n_630), .Y(n_662) );
AND2x2_ASAP7_75t_L g696 ( .A(n_589), .B(n_598), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_590), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g706 ( .A(n_590), .Y(n_706) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_594), .A2(n_622), .B1(n_624), .B2(n_629), .Y(n_621) );
OAI22xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B1(n_599), .B2(n_600), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_596), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_631) );
INVxp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_601), .A2(n_703), .B1(n_705), .B2(n_707), .C(n_711), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B(n_610), .C(n_631), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g672 ( .A(n_608), .B(n_625), .Y(n_672) );
INVx1_ASAP7_75t_L g723 ( .A(n_608), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_609), .A2(n_611), .B1(n_615), .B2(n_618), .C(n_621), .Y(n_610) );
INVx2_ASAP7_75t_SL g665 ( .A(n_609), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g730 ( .A(n_612), .Y(n_730) );
AND2x2_ASAP7_75t_L g654 ( .A(n_613), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g639 ( .A(n_614), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g701 ( .A(n_617), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_625), .B(n_727), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g625 ( .A(n_626), .Y(n_625) );
INVxp67_ASAP7_75t_L g670 ( .A(n_628), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_629), .A2(n_641), .B(n_643), .C(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g718 ( .A(n_632), .Y(n_718) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_636), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx2_ASAP7_75t_L g649 ( .A(n_639), .Y(n_649) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI222xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_652), .B1(n_653), .B2(n_656), .C1(n_657), .C2(n_659), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g685 ( .A(n_649), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_652), .B(n_706), .Y(n_705) );
NAND2xp33_ASAP7_75t_SL g683 ( .A(n_653), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g658 ( .A(n_655), .Y(n_658) );
AND2x2_ASAP7_75t_L g722 ( .A(n_655), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g688 ( .A(n_658), .B(n_685), .Y(n_688) );
INVx1_ASAP7_75t_L g717 ( .A(n_659), .Y(n_717) );
AOI211xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B(n_666), .C(n_671), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_665), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g716 ( .A1(n_668), .A2(n_696), .A3(n_701), .B1(n_717), .B2(n_718), .C1(n_719), .C2(n_722), .Y(n_716) );
AND2x2_ASAP7_75t_L g703 ( .A(n_669), .B(n_704), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_674), .B2(n_676), .Y(n_671) );
INVxp33_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B1(n_683), .B2(n_686), .C(n_687), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NAND5xp2_ASAP7_75t_L g690 ( .A(n_691), .B(n_702), .C(n_716), .D(n_724), .E(n_728), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B(n_697), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp33_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_704), .A2(n_729), .B(n_730), .C(n_731), .Y(n_728) );
AOI31xp33_ASAP7_75t_L g711 ( .A1(n_706), .A2(n_712), .A3(n_713), .B(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g729 ( .A(n_727), .Y(n_729) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g750 ( .A(n_736), .Y(n_750) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_743), .Y(n_746) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx3_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
endmodule