module fake_jpeg_24982_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_16),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_12),
.B1(n_10),
.B2(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_7),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_19),
.B1(n_15),
.B2(n_14),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_23),
.B1(n_0),
.B2(n_1),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_6),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_13),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_0),
.B(n_2),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_32),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_29),
.C(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_31),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_3),
.C(n_30),
.Y(n_39)
);


endmodule