module real_jpeg_4042_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_1),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_43),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_43),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_43),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_25),
.B1(n_102),
.B2(n_106),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_25),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_25),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_30),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_3),
.A2(n_335),
.B(n_337),
.C(n_343),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_3),
.B(n_85),
.C(n_164),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_3),
.B(n_141),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_3),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_3),
.B(n_89),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_4),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_4),
.A2(n_218),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_4),
.A2(n_218),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_4),
.A2(n_218),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_6),
.Y(n_166)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_6),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_6),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_8),
.Y(n_264)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_11),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_11),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_12),
.A2(n_32),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_12),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_12),
.A2(n_131),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_131),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_131),
.B1(n_164),
.B2(n_269),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_445),
.Y(n_19)
);

OAI221xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_58),
.B1(n_62),
.B2(n_440),
.C(n_443),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_21),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_21),
.B(n_58),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_22),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_23),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_47),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_28),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g337 ( 
.A1(n_25),
.A2(n_338),
.B(n_340),
.Y(n_337)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_26),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_27),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_28),
.Y(n_219)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_30),
.B(n_216),
.Y(n_247)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_31),
.B(n_117),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_32),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_111)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_34),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_34),
.Y(n_211)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_40),
.A2(n_60),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_40),
.B(n_247),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_47),
.B(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_58),
.A2(n_158),
.B(n_185),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_160),
.B1(n_185),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_58),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B(n_61),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_59),
.A2(n_71),
.B(n_226),
.Y(n_436)
);

A2O1A1O1Ixp25_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_240),
.B(n_429),
.C(n_432),
.D(n_439),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_220),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_186),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_65),
.B(n_186),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_157),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_142),
.B2(n_143),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_68),
.B(n_142),
.C(n_157),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_69),
.A2(n_70),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_70),
.B(n_75),
.C(n_108),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_70),
.B(n_223),
.C(n_238),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_71),
.B(n_215),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_72),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_107),
.B2(n_108),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_75),
.A2(n_76),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_75),
.A2(n_76),
.B1(n_249),
.B2(n_257),
.Y(n_248)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_76),
.B(n_246),
.C(n_249),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_76),
.B(n_234),
.C(n_237),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_99),
.B(n_100),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_77),
.A2(n_178),
.B(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_78),
.B(n_101),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_78),
.B(n_349),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_82),
.Y(n_350)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_83),
.Y(n_342)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_87),
.Y(n_180)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_89),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_89),
.B(n_349),
.Y(n_365)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_92),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_93),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_96),
.Y(n_374)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_100),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_99),
.A2(n_147),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_128),
.B(n_132),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_109),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_109),
.B(n_252),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_109),
.A2(n_141),
.B(n_209),
.Y(n_305)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_110),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_118),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_113),
.Y(n_336)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_114),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_118),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_124),
.Y(n_353)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_141),
.B(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_133),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_133),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_140),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_141),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_144),
.B(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_154),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_145),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_147),
.B(n_365),
.Y(n_409)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_155),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_159),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_177),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_160),
.A2(n_177),
.B1(n_185),
.B2(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_160),
.B(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_160),
.A2(n_185),
.B1(n_334),
.B2(n_412),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B(n_169),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_161),
.B(n_169),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_161),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_161),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_177),
.Y(n_317)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_184),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_184),
.B(n_348),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_193),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_187),
.A2(n_191),
.B1(n_192),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_187),
.Y(n_321)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_193),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_207),
.C(n_214),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_194),
.A2(n_195),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_196),
.B(n_206),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_197),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_199),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_268),
.B(n_270),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_201),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_205),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_207),
.B(n_214),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_208),
.B(n_251),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_209),
.Y(n_236)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_220),
.A2(n_430),
.B(n_431),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_239),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_221),
.B(n_239),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_231),
.B1(n_232),
.B2(n_237),
.Y(n_224)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_261),
.A3(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_260)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_421),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_310),
.C(n_324),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_297),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_283),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_244),
.B(n_283),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_258),
.C(n_273),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_245),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_258),
.A2(n_259),
.B1(n_273),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_280),
.B(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_272),
.Y(n_396)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_278),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_279),
.B(n_386),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_280),
.B(n_369),
.Y(n_399)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_286),
.C(n_291),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_290),
.B(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_297),
.A2(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_309),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_298),
.B(n_309),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_305),
.A2(n_307),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_305),
.B(n_436),
.C(n_437),
.Y(n_442)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_322),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_311),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_312),
.B(n_323),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_312),
.B(n_319),
.Y(n_428)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_316),
.CI(n_318),
.CON(n_312),
.SN(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_354),
.B(n_420),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_326),
.B(n_329),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.C(n_345),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_330),
.B(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_333),
.A2(n_345),
.B1(n_346),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_414),
.B(n_419),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_404),
.B(n_413),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_380),
.B(n_403),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_366),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_358),
.B(n_366),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_364),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_359),
.A2(n_360),
.B1(n_364),
.B2(n_383),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_375),
.Y(n_366)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_378),
.C(n_406),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_389),
.B(n_402),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_384),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_398),
.B(n_401),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_397),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_399),
.B(n_400),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_407),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_410),
.C(n_411),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_418),
.Y(n_419)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g421 ( 
.A1(n_422),
.A2(n_423),
.B(n_426),
.C(n_427),
.D(n_428),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_438),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_438),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_442),
.Y(n_444)
);


endmodule