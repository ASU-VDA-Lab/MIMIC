module fake_ariane_1974_n_1395 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_155, n_127, n_1395);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_155;
input n_127;

output n_1395;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

INVx2_ASAP7_75t_SL g356 ( 
.A(n_16),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_222),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_192),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_9),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_119),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_113),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_201),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_137),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_351),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_255),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_252),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_315),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_265),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_38),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_330),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_322),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_228),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_172),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_176),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_196),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_126),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_336),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_165),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_68),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_307),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_287),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_263),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_189),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_84),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_293),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_20),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_251),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_142),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_204),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_225),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_153),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_13),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_43),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_158),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_212),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_69),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_70),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_85),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_112),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_130),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_312),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_106),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_262),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_145),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_134),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_338),
.Y(n_411)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_297),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_29),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_257),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_304),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_195),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_285),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_268),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_168),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_327),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_29),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_340),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_131),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_69),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_260),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_279),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_199),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_281),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_230),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_169),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_15),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_180),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_104),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_98),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_95),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_46),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_19),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_125),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_152),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_220),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_242),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_346),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_53),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_184),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_217),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_105),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_348),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_250),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_300),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_84),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_303),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_140),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_47),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_59),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_58),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_88),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_191),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_354),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_232),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_209),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_229),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_167),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_73),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_298),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_299),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_256),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_236),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_91),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_332),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_101),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_53),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_352),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_58),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_243),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_221),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_88),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_355),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_22),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_87),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_301),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_302),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_33),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_277),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_162),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_82),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_306),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_118),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_46),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_144),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_127),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_49),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_237),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_213),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_289),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_188),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_278),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_231),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_291),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_309),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_325),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_120),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_305),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_35),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_87),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_271),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_334),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_65),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_179),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_38),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_154),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_311),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_219),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_143),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_224),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_333),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_163),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_324),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_280),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_335),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_31),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_216),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_339),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_227),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_82),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_249),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_5),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_347),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_68),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_296),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_183),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_170),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_206),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_60),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_178),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_115),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_107),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_239),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_254),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_27),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_282),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_40),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_382),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_367),
.B(n_0),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_369),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_0),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_382),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_382),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_1),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_397),
.B(n_1),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_402),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_418),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_494),
.B(n_2),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_443),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_523),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_435),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_382),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_382),
.B(n_2),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_402),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_444),
.B(n_3),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_523),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_444),
.B(n_3),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_523),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_523),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_366),
.Y(n_573)
);

BUFx8_ASAP7_75t_SL g574 ( 
.A(n_432),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_359),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_472),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_504),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_363),
.B(n_4),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_366),
.B(n_4),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_359),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_435),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_386),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_382),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_472),
.B(n_5),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_537),
.B(n_6),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_537),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_365),
.B(n_6),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_370),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_525),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_400),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_386),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_374),
.B(n_7),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_404),
.B(n_7),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_399),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_377),
.B(n_8),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_525),
.Y(n_596)
);

CKINVDCx11_ASAP7_75t_R g597 ( 
.A(n_508),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_399),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_408),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_439),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_378),
.B(n_8),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_381),
.B(n_9),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_408),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_404),
.B(n_10),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_467),
.B(n_10),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_467),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_525),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_383),
.B(n_11),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_387),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_389),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_422),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_425),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_361),
.Y(n_616)
);

BUFx8_ASAP7_75t_SL g617 ( 
.A(n_376),
.Y(n_617)
);

BUFx8_ASAP7_75t_L g618 ( 
.A(n_356),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_357),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_396),
.B(n_11),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_451),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_392),
.B(n_12),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_398),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_510),
.B(n_12),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_455),
.B(n_13),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_358),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_401),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_361),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_384),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_459),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_464),
.B(n_477),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_384),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_527),
.B(n_14),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_479),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_403),
.B(n_14),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_426),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_406),
.B(n_15),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_414),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_437),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_426),
.B(n_92),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_483),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_461),
.B(n_93),
.Y(n_642)
);

BUFx12f_ASAP7_75t_L g643 ( 
.A(n_438),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_407),
.B(n_16),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_548),
.A2(n_376),
.B1(n_466),
.B2(n_456),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

AO22x2_ASAP7_75t_L g647 ( 
.A1(n_559),
.A2(n_492),
.B1(n_505),
.B2(n_486),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_590),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_593),
.A2(n_457),
.B1(n_474),
.B2(n_454),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_605),
.A2(n_489),
.B1(n_529),
.B2(n_480),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_545),
.A2(n_540),
.B1(n_534),
.B2(n_415),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_545),
.A2(n_420),
.B1(n_423),
.B2(n_405),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_560),
.B(n_521),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_559),
.A2(n_578),
.B1(n_633),
.B2(n_624),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_594),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_629),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_596),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_601),
.A2(n_468),
.B1(n_491),
.B2(n_458),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_630),
.A2(n_496),
.B1(n_513),
.B2(n_461),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_587),
.A2(n_538),
.B1(n_513),
.B2(n_522),
.Y(n_662)
);

OA22x2_ASAP7_75t_L g663 ( 
.A1(n_588),
.A2(n_419),
.B1(n_429),
.B2(n_416),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_581),
.B(n_496),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_604),
.B(n_627),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_578),
.A2(n_497),
.B1(n_531),
.B2(n_522),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_606),
.A2(n_531),
.B1(n_433),
.B2(n_440),
.Y(n_668)
);

AOI22x1_ASAP7_75t_SL g669 ( 
.A1(n_617),
.A2(n_447),
.B1(n_450),
.B2(n_430),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_620),
.A2(n_470),
.B1(n_475),
.B2(n_465),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_556),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_546),
.B(n_360),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_617),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_609),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_556),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_556),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_620),
.A2(n_482),
.B1(n_484),
.B2(n_476),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_640),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_629),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_564),
.A2(n_503),
.B1(n_519),
.B2(n_493),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_555),
.B(n_362),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_613),
.B(n_520),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_638),
.A2(n_535),
.B1(n_533),
.B2(n_368),
.Y(n_684)
);

AO22x2_ASAP7_75t_L g685 ( 
.A1(n_554),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_558),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_568),
.A2(n_371),
.B1(n_372),
.B2(n_364),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_SL g689 ( 
.A1(n_639),
.A2(n_375),
.B1(n_379),
.B2(n_373),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_561),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_623),
.B(n_380),
.Y(n_691)
);

OA22x2_ASAP7_75t_L g692 ( 
.A1(n_588),
.A2(n_388),
.B1(n_390),
.B2(n_385),
.Y(n_692)
);

AO22x2_ASAP7_75t_L g693 ( 
.A1(n_554),
.A2(n_584),
.B1(n_570),
.B2(n_631),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_629),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_567),
.B(n_391),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_561),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_643),
.B(n_17),
.Y(n_697)
);

OA22x2_ASAP7_75t_L g698 ( 
.A1(n_631),
.A2(n_394),
.B1(n_395),
.B2(n_393),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_561),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_597),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_562),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_592),
.A2(n_410),
.B1(n_411),
.B2(n_409),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_570),
.A2(n_421),
.B1(n_424),
.B2(n_417),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_576),
.B(n_427),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_584),
.B(n_428),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_431),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_595),
.A2(n_610),
.B1(n_622),
.B2(n_602),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_434),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_625),
.B(n_436),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_579),
.Y(n_710)
);

AND2x2_ASAP7_75t_SL g711 ( 
.A(n_625),
.B(n_441),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_603),
.A2(n_446),
.B1(n_448),
.B2(n_445),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_595),
.A2(n_452),
.B1(n_453),
.B2(n_449),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_619),
.B(n_460),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_602),
.A2(n_463),
.B1(n_469),
.B2(n_462),
.Y(n_715)
);

AOI22x1_ASAP7_75t_SL g716 ( 
.A1(n_574),
.A2(n_473),
.B1(n_478),
.B2(n_471),
.Y(n_716)
);

NAND3x1_ASAP7_75t_L g717 ( 
.A(n_610),
.B(n_18),
.C(n_20),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_622),
.A2(n_487),
.B1(n_488),
.B2(n_481),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_637),
.A2(n_495),
.B1(n_498),
.B2(n_490),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_603),
.A2(n_500),
.B1(n_501),
.B2(n_499),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_SL g722 ( 
.A1(n_635),
.A2(n_506),
.B1(n_507),
.B2(n_502),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_635),
.A2(n_511),
.B1(n_512),
.B2(n_509),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_644),
.A2(n_515),
.B1(n_516),
.B2(n_514),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_580),
.B(n_517),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_637),
.A2(n_524),
.B1(n_526),
.B2(n_518),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_550),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_665),
.B(n_666),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_678),
.B(n_586),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_648),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_655),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_657),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_657),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_645),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_666),
.B(n_580),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_664),
.B(n_614),
.Y(n_736)
);

AND2x6_ASAP7_75t_L g737 ( 
.A(n_654),
.B(n_652),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_707),
.B(n_573),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_718),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_679),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_679),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_710),
.B(n_619),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_694),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_694),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_646),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_710),
.B(n_626),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_693),
.B(n_573),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_693),
.B(n_691),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_714),
.B(n_626),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_651),
.B(n_579),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_658),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_706),
.B(n_615),
.Y(n_752)
);

XNOR2xp5_ASAP7_75t_L g753 ( 
.A(n_673),
.B(n_574),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_708),
.B(n_621),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_660),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_674),
.Y(n_756)
);

XNOR2xp5_ASAP7_75t_L g757 ( 
.A(n_700),
.B(n_577),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_656),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_718),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_R g760 ( 
.A(n_672),
.B(n_641),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_675),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_676),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_714),
.B(n_591),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_682),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_689),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_681),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_705),
.B(n_585),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_687),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_690),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_709),
.B(n_644),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_671),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_SL g773 ( 
.A(n_711),
.B(n_640),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_725),
.B(n_582),
.Y(n_774)
);

XOR2xp5_ASAP7_75t_L g775 ( 
.A(n_716),
.B(n_577),
.Y(n_775)
);

XOR2x2_ASAP7_75t_L g776 ( 
.A(n_661),
.B(n_597),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_695),
.A2(n_566),
.B(n_551),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_705),
.B(n_582),
.Y(n_778)
);

AND2x2_ASAP7_75t_SL g779 ( 
.A(n_668),
.B(n_550),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_688),
.B(n_618),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_696),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_699),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_701),
.Y(n_783)
);

XOR2xp5_ASAP7_75t_L g784 ( 
.A(n_716),
.B(n_608),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_703),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_667),
.A2(n_566),
.B(n_585),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_704),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_671),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_671),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_712),
.B(n_618),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_663),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_653),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_653),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_647),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_647),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_677),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_662),
.Y(n_797)
);

XNOR2xp5_ASAP7_75t_L g798 ( 
.A(n_659),
.B(n_553),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_670),
.A2(n_553),
.B(n_552),
.Y(n_799)
);

XOR2xp5_ASAP7_75t_L g800 ( 
.A(n_669),
.B(n_608),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_677),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_698),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_692),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_721),
.A2(n_565),
.B(n_543),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

AND2x6_ASAP7_75t_L g806 ( 
.A(n_680),
.B(n_583),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_650),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_723),
.B(n_608),
.Y(n_808)
);

XOR2xp5_ASAP7_75t_L g809 ( 
.A(n_669),
.B(n_611),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_683),
.B(n_684),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_722),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_685),
.A2(n_642),
.B(n_640),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_724),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_685),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_717),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_702),
.B(n_611),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_727),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_727),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_683),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_772),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_735),
.B(n_752),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_730),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_728),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_796),
.B(n_697),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_731),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_760),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_778),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_738),
.B(n_726),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_772),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_768),
.B(n_720),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_768),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_778),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_801),
.B(n_697),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_794),
.B(n_678),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_754),
.B(n_736),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_745),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_739),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_774),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_742),
.B(n_713),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_751),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_797),
.B(n_779),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_746),
.B(n_715),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_737),
.B(n_719),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_806),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_737),
.B(n_611),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_764),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_737),
.B(n_586),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_732),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_761),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_737),
.B(n_813),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_755),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_795),
.B(n_678),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_786),
.B(n_629),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_792),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_750),
.B(n_808),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_756),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_750),
.B(n_586),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_750),
.B(n_586),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_733),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_740),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_815),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_777),
.A2(n_804),
.B(n_799),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_771),
.B(n_594),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_773),
.B(n_632),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_814),
.B(n_594),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_750),
.B(n_616),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_787),
.B(n_632),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_799),
.B(n_632),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_791),
.B(n_632),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_806),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_793),
.B(n_636),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_805),
.B(n_636),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_747),
.B(n_616),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_743),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_744),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_758),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_749),
.B(n_628),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_804),
.A2(n_642),
.B(n_640),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_759),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_763),
.A2(n_642),
.B(n_640),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_748),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_798),
.B(n_628),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_807),
.B(n_636),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_762),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_766),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_817),
.B(n_636),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_767),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_818),
.B(n_591),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_773),
.B(n_591),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_816),
.B(n_412),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_757),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_753),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_802),
.B(n_591),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_812),
.A2(n_729),
.B(n_769),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_810),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_790),
.B(n_598),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_803),
.B(n_642),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_770),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_788),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_780),
.B(n_598),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_819),
.B(n_598),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_781),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_782),
.B(n_598),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_784),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_783),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_765),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_811),
.B(n_600),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_840),
.B(n_785),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_873),
.B(n_776),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_821),
.B(n_734),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_863),
.Y(n_915)
);

AND2x6_ASAP7_75t_L g916 ( 
.A(n_892),
.B(n_544),
.Y(n_916)
);

INVx8_ASAP7_75t_L g917 ( 
.A(n_873),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_843),
.B(n_600),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_833),
.B(n_600),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_828),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_841),
.B(n_528),
.Y(n_921)
);

NAND2x1_ASAP7_75t_SL g922 ( 
.A(n_846),
.B(n_800),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_821),
.B(n_809),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_850),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_857),
.B(n_775),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_894),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_836),
.B(n_600),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_843),
.B(n_607),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_826),
.B(n_607),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_823),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_867),
.B(n_607),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_889),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_844),
.B(n_607),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_867),
.B(n_21),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_832),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_873),
.B(n_824),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_824),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_829),
.B(n_530),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_895),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_846),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_850),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_846),
.B(n_532),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_899),
.B(n_536),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_828),
.Y(n_944)
);

BUFx8_ASAP7_75t_L g945 ( 
.A(n_824),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_899),
.B(n_539),
.Y(n_946)
);

AND2x2_ASAP7_75t_SL g947 ( 
.A(n_866),
.B(n_863),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_903),
.B(n_541),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_910),
.B(n_23),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_910),
.B(n_24),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_832),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_889),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_910),
.B(n_24),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_903),
.B(n_25),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_827),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_822),
.Y(n_956)
);

BUFx8_ASAP7_75t_SL g957 ( 
.A(n_911),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_825),
.Y(n_958)
);

AO21x2_ASAP7_75t_L g959 ( 
.A1(n_893),
.A2(n_413),
.B(n_412),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_874),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_867),
.B(n_25),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_874),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_836),
.B(n_549),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_837),
.B(n_911),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_837),
.B(n_549),
.Y(n_965)
);

NAND2x1_ASAP7_75t_L g966 ( 
.A(n_832),
.B(n_544),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_884),
.B(n_26),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_911),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_871),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_863),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_873),
.Y(n_971)
);

NAND2x1_ASAP7_75t_L g972 ( 
.A(n_862),
.B(n_544),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_861),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_834),
.B(n_852),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_871),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_848),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_820),
.B(n_549),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_834),
.B(n_562),
.Y(n_978)
);

BUFx4f_ASAP7_75t_L g979 ( 
.A(n_834),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_884),
.B(n_26),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_898),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_861),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_828),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_885),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_875),
.B(n_27),
.Y(n_985)
);

BUFx4f_ASAP7_75t_L g986 ( 
.A(n_904),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_917),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_945),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_984),
.B(n_845),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_917),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_947),
.B(n_855),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_934),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_956),
.Y(n_993)
);

INVx6_ASAP7_75t_L g994 ( 
.A(n_945),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_958),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_937),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_924),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_979),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_935),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_936),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_920),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_928),
.B(n_856),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_935),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_976),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_941),
.Y(n_1006)
);

BUFx2_ASAP7_75t_SL g1007 ( 
.A(n_939),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_973),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_982),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_926),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_934),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_936),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_967),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_928),
.B(n_869),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_957),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_964),
.B(n_869),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_967),
.Y(n_1017)
);

BUFx10_ASAP7_75t_L g1018 ( 
.A(n_949),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_970),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_981),
.Y(n_1020)
);

AND2x2_ASAP7_75t_SL g1021 ( 
.A(n_980),
.B(n_866),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_980),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_976),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_930),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_932),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_912),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_952),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_940),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_940),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_930),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_974),
.B(n_855),
.Y(n_1031)
);

CKINVDCx6p67_ASAP7_75t_R g1032 ( 
.A(n_978),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_986),
.Y(n_1033)
);

INVx3_ASAP7_75t_SL g1034 ( 
.A(n_912),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_951),
.B(n_831),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_969),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_951),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_971),
.B(n_820),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_914),
.A2(n_907),
.B1(n_854),
.B2(n_835),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_975),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_955),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_920),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_944),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_960),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_944),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_978),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_962),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_944),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_983),
.Y(n_1049)
);

INVx8_ASAP7_75t_L g1050 ( 
.A(n_974),
.Y(n_1050)
);

CKINVDCx11_ASAP7_75t_R g1051 ( 
.A(n_913),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_1015),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_1007),
.Y(n_1053)
);

CKINVDCx11_ASAP7_75t_R g1054 ( 
.A(n_1015),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_992),
.A2(n_950),
.B1(n_953),
.B2(n_954),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1021),
.A2(n_925),
.B1(n_923),
.B2(n_913),
.Y(n_1056)
);

OAI22xp33_ASAP7_75t_SL g1057 ( 
.A1(n_1034),
.A2(n_938),
.B1(n_919),
.B2(n_921),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_993),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_SL g1059 ( 
.A1(n_1021),
.A2(n_968),
.B1(n_942),
.B2(n_864),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_SL g1060 ( 
.A1(n_1026),
.A2(n_865),
.B1(n_961),
.B2(n_985),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_1026),
.A2(n_918),
.B1(n_879),
.B2(n_931),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_1029),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1039),
.A2(n_879),
.B1(n_931),
.B2(n_890),
.Y(n_1063)
);

CKINVDCx11_ASAP7_75t_R g1064 ( 
.A(n_988),
.Y(n_1064)
);

INVx6_ASAP7_75t_L g1065 ( 
.A(n_990),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_SL g1066 ( 
.A(n_988),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1024),
.A2(n_946),
.B1(n_948),
.B2(n_943),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_995),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_1010),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_1010),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1025),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1036),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1040),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1009),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1020),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_989),
.A2(n_870),
.B1(n_881),
.B2(n_847),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1034),
.A2(n_890),
.B1(n_901),
.B2(n_887),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_991),
.A2(n_915),
.B1(n_860),
.B2(n_859),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_1051),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1016),
.A2(n_1005),
.B1(n_1014),
.B2(n_1024),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1030),
.A2(n_862),
.B1(n_878),
.B2(n_872),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_991),
.A2(n_870),
.B1(n_892),
.B2(n_916),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1002),
.A2(n_901),
.B1(n_905),
.B2(n_887),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_1037),
.A2(n_933),
.B(n_849),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1030),
.B(n_922),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_1051),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1020),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_994),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1027),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_SL g1090 ( 
.A1(n_1013),
.A2(n_916),
.B1(n_886),
.B2(n_875),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_996),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1044),
.Y(n_1092)
);

CKINVDCx11_ASAP7_75t_R g1093 ( 
.A(n_996),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1009),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_994),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1044),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1017),
.A2(n_916),
.B1(n_886),
.B2(n_838),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1022),
.A2(n_842),
.B1(n_858),
.B2(n_853),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1047),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_998),
.B(n_983),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_994),
.Y(n_1101)
);

NAND2x1p5_ASAP7_75t_L g1102 ( 
.A(n_998),
.B(n_983),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_997),
.A2(n_905),
.B1(n_877),
.B2(n_929),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1047),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1023),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1006),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1008),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1011),
.A2(n_1031),
.B1(n_908),
.B2(n_888),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1062),
.A2(n_1023),
.B1(n_1028),
.B2(n_1041),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1058),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1062),
.A2(n_1032),
.B1(n_1028),
.B2(n_1046),
.Y(n_1111)
);

OAI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_1055),
.A2(n_882),
.B(n_862),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1056),
.A2(n_1018),
.B1(n_1032),
.B2(n_891),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1067),
.A2(n_1028),
.B1(n_1037),
.B2(n_999),
.Y(n_1114)
);

AOI211xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1057),
.A2(n_1049),
.B(n_868),
.C(n_830),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1080),
.A2(n_1033),
.B1(n_1018),
.B2(n_1019),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1068),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1056),
.A2(n_851),
.B1(n_902),
.B2(n_876),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1071),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1060),
.A2(n_1037),
.B1(n_999),
.B2(n_1003),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1096),
.Y(n_1121)
);

BUFx8_ASAP7_75t_L g1122 ( 
.A(n_1079),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1105),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1075),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1070),
.B(n_1019),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1081),
.A2(n_999),
.B1(n_1003),
.B2(n_987),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1059),
.A2(n_854),
.B1(n_835),
.B2(n_904),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1088),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1087),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1089),
.B(n_1000),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1063),
.A2(n_891),
.B1(n_1050),
.B2(n_1012),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1085),
.A2(n_1050),
.B1(n_1012),
.B2(n_1000),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1059),
.A2(n_839),
.B1(n_1050),
.B2(n_1035),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1072),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1064),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1082),
.A2(n_839),
.B1(n_1050),
.B2(n_1035),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1069),
.B(n_987),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1073),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1053),
.A2(n_990),
.B(n_965),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1077),
.A2(n_1003),
.B1(n_987),
.B2(n_972),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1099),
.A2(n_839),
.B1(n_900),
.B2(n_909),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1092),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1098),
.A2(n_1038),
.B1(n_990),
.B2(n_1049),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1101),
.A2(n_900),
.B1(n_927),
.B2(n_959),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1106),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1098),
.A2(n_900),
.B1(n_909),
.B2(n_906),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1076),
.A2(n_990),
.B(n_1038),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1076),
.A2(n_880),
.B(n_1049),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1061),
.A2(n_909),
.B1(n_963),
.B2(n_896),
.Y(n_1149)
);

AO22x1_ASAP7_75t_L g1150 ( 
.A1(n_1091),
.A2(n_990),
.B1(n_1042),
.B2(n_1045),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_SL g1151 ( 
.A1(n_1095),
.A2(n_909),
.B1(n_883),
.B2(n_1001),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1107),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1104),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1054),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1103),
.A2(n_909),
.B1(n_896),
.B2(n_897),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1097),
.A2(n_1038),
.B(n_1004),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1074),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1094),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1088),
.B(n_1042),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1100),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1083),
.A2(n_1048),
.B1(n_1045),
.B2(n_1004),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1097),
.A2(n_1004),
.B(n_1001),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1086),
.A2(n_1004),
.B1(n_1043),
.B2(n_1001),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1078),
.A2(n_1048),
.B1(n_1045),
.B2(n_830),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1090),
.A2(n_1004),
.B(n_1001),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1108),
.A2(n_1048),
.B1(n_1043),
.B2(n_1001),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1090),
.A2(n_1043),
.B1(n_413),
.B2(n_412),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1093),
.A2(n_1043),
.B1(n_413),
.B2(n_412),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1100),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1102),
.B(n_1043),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1102),
.B(n_830),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1066),
.A2(n_413),
.B1(n_412),
.B2(n_828),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1065),
.A2(n_966),
.B1(n_977),
.B2(n_31),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1052),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1065),
.Y(n_1175)
);

OAI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1116),
.A2(n_1084),
.B1(n_1065),
.B2(n_966),
.C(n_33),
.Y(n_1176)
);

AOI222xp33_ASAP7_75t_L g1177 ( 
.A1(n_1113),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.C1(n_34),
.C2(n_35),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1110),
.B(n_28),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1135),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1113),
.A2(n_413),
.B1(n_412),
.B2(n_562),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1167),
.A2(n_39),
.B1(n_36),
.B2(n_37),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1117),
.A2(n_572),
.B1(n_571),
.B2(n_569),
.C(n_547),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1119),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1134),
.B(n_36),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1115),
.B(n_547),
.C(n_544),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1118),
.A2(n_413),
.B1(n_563),
.B2(n_547),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1138),
.B(n_37),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1127),
.A2(n_563),
.B1(n_569),
.B2(n_547),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1131),
.A2(n_571),
.B1(n_572),
.B2(n_569),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1152),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1123),
.B(n_39),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1136),
.A2(n_557),
.B1(n_42),
.B2(n_41),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1125),
.B(n_44),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1158),
.A2(n_557),
.B1(n_47),
.B2(n_44),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1165),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1142),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1143),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1133),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1122),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1121),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1109),
.B(n_54),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1162),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_1202)
);

AOI222xp33_ASAP7_75t_L g1203 ( 
.A1(n_1148),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.C1(n_62),
.C2(n_63),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_L g1204 ( 
.A(n_1111),
.B(n_61),
.C(n_62),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1114),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1120),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1168),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1145),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1208)
);

OA222x2_ASAP7_75t_L g1209 ( 
.A1(n_1156),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.C1(n_75),
.C2(n_76),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1168),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1112),
.A2(n_1149),
.B1(n_1146),
.B2(n_1155),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1129),
.B(n_77),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1157),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1172),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1157),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_1215)
);

OAI222xp33_ASAP7_75t_L g1216 ( 
.A1(n_1132),
.A2(n_81),
.B1(n_83),
.B2(n_85),
.C1(n_86),
.C2(n_89),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1153),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1139),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1130),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1163),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1174),
.A2(n_1166),
.B1(n_1151),
.B2(n_1122),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1169),
.Y(n_1222)
);

OAI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1147),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1166),
.A2(n_114),
.B(n_116),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1154),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1175),
.B(n_123),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1137),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_1227)
);

OAI221xp5_ASAP7_75t_L g1228 ( 
.A1(n_1173),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.C(n_136),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1164),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.C(n_146),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1141),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_1230)
);

AOI222xp33_ASAP7_75t_L g1231 ( 
.A1(n_1124),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.C1(n_156),
.C2(n_157),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1160),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1144),
.A2(n_164),
.B1(n_166),
.B2(n_171),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1183),
.B(n_1128),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1202),
.A2(n_1128),
.B(n_1126),
.Y(n_1235)
);

NOR3xp33_ASAP7_75t_L g1236 ( 
.A(n_1195),
.B(n_1216),
.C(n_1204),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1190),
.B(n_1159),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1196),
.B(n_1150),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1203),
.B(n_1170),
.C(n_1171),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1193),
.B(n_1160),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1201),
.A2(n_1209),
.B(n_1177),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1195),
.B(n_1140),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1178),
.B(n_1160),
.Y(n_1243)
);

NOR3xp33_ASAP7_75t_L g1244 ( 
.A(n_1223),
.B(n_1176),
.C(n_1206),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1223),
.A2(n_1161),
.B(n_1160),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1211),
.A2(n_1161),
.B1(n_174),
.B2(n_175),
.Y(n_1246)
);

OAI221xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1197),
.A2(n_1198),
.B1(n_1213),
.B2(n_1215),
.C(n_1217),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1191),
.B(n_353),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1184),
.B(n_173),
.Y(n_1249)
);

NAND2xp33_ASAP7_75t_SL g1250 ( 
.A(n_1199),
.B(n_177),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1212),
.B(n_181),
.Y(n_1251)
);

AND2x2_ASAP7_75t_SL g1252 ( 
.A(n_1224),
.B(n_182),
.Y(n_1252)
);

AND2x2_ASAP7_75t_SL g1253 ( 
.A(n_1224),
.B(n_185),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1187),
.B(n_350),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1222),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1179),
.B(n_349),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1205),
.B(n_186),
.C(n_187),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1225),
.B(n_190),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1211),
.B(n_345),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1231),
.B(n_193),
.C(n_194),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1214),
.A2(n_197),
.B(n_198),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1226),
.B(n_200),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1221),
.B(n_344),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1221),
.B(n_202),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1218),
.B(n_203),
.Y(n_1265)
);

AOI211xp5_ASAP7_75t_L g1266 ( 
.A1(n_1181),
.A2(n_205),
.B(n_207),
.C(n_208),
.Y(n_1266)
);

NAND4xp25_ASAP7_75t_L g1267 ( 
.A(n_1208),
.B(n_343),
.C(n_211),
.D(n_214),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1207),
.A2(n_210),
.B(n_215),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1200),
.B(n_218),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1210),
.B(n_223),
.C(n_226),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1224),
.B(n_341),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1185),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1227),
.A2(n_233),
.B(n_234),
.Y(n_1273)
);

NAND4xp25_ASAP7_75t_SL g1274 ( 
.A(n_1192),
.B(n_235),
.C(n_238),
.D(n_240),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1180),
.B(n_241),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1188),
.Y(n_1276)
);

OAI221xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1180),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.C(n_247),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1229),
.B(n_248),
.C(n_253),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1256),
.B(n_1262),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1234),
.B(n_1194),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1238),
.B(n_1233),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1240),
.B(n_1220),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1237),
.B(n_1228),
.Y(n_1283)
);

NAND4xp75_ASAP7_75t_L g1284 ( 
.A(n_1241),
.B(n_1182),
.C(n_1232),
.D(n_1230),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1285)
);

NAND4xp75_ASAP7_75t_L g1286 ( 
.A(n_1258),
.B(n_1230),
.C(n_1219),
.D(n_1189),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1244),
.A2(n_1186),
.B1(n_259),
.B2(n_261),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1255),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1248),
.B(n_258),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1243),
.B(n_264),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1272),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1251),
.B(n_266),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1239),
.B(n_267),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1250),
.B(n_1235),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1272),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1242),
.B(n_269),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1245),
.B(n_270),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1236),
.B(n_272),
.C(n_273),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1252),
.B(n_274),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1236),
.B(n_275),
.C(n_276),
.Y(n_1300)
);

AOI211xp5_ASAP7_75t_L g1301 ( 
.A1(n_1261),
.A2(n_283),
.B(n_284),
.C(n_286),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1259),
.B(n_288),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1253),
.B(n_1271),
.Y(n_1303)
);

NAND4xp25_ASAP7_75t_L g1304 ( 
.A(n_1294),
.B(n_1247),
.C(n_1265),
.D(n_1273),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1279),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1295),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1291),
.B(n_1253),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1303),
.B(n_1265),
.Y(n_1308)
);

NAND4xp75_ASAP7_75t_SL g1309 ( 
.A(n_1283),
.B(n_1275),
.C(n_1260),
.D(n_1266),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1285),
.B(n_1276),
.Y(n_1310)
);

NOR3xp33_ASAP7_75t_L g1311 ( 
.A(n_1298),
.B(n_1274),
.C(n_1257),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1303),
.B(n_1268),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1280),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1288),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1280),
.B(n_1263),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1296),
.B(n_1246),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1289),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1293),
.Y(n_1318)
);

XOR2x2_ASAP7_75t_L g1319 ( 
.A(n_1284),
.B(n_1264),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1282),
.Y(n_1320)
);

NOR3xp33_ASAP7_75t_L g1321 ( 
.A(n_1300),
.B(n_1267),
.C(n_1270),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1281),
.B(n_1246),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1313),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1313),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1320),
.B(n_1281),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1314),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1306),
.B(n_1296),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1317),
.Y(n_1328)
);

XOR2x2_ASAP7_75t_L g1329 ( 
.A(n_1319),
.B(n_1286),
.Y(n_1329)
);

CKINVDCx8_ASAP7_75t_R g1330 ( 
.A(n_1305),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1320),
.B(n_1315),
.Y(n_1331)
);

XNOR2xp5_ASAP7_75t_L g1332 ( 
.A(n_1319),
.B(n_1292),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1314),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1322),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1331),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1334),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1330),
.A2(n_1305),
.B1(n_1317),
.B2(n_1318),
.Y(n_1337)
);

OAI22x1_ASAP7_75t_L g1338 ( 
.A1(n_1332),
.A2(n_1308),
.B1(n_1322),
.B2(n_1312),
.Y(n_1338)
);

XOR2x2_ASAP7_75t_L g1339 ( 
.A(n_1329),
.B(n_1309),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1334),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1324),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1327),
.Y(n_1342)
);

AOI22x1_ASAP7_75t_L g1343 ( 
.A1(n_1323),
.A2(n_1308),
.B1(n_1315),
.B2(n_1304),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1325),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1326),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1333),
.Y(n_1346)
);

AOI322xp5_ASAP7_75t_L g1347 ( 
.A1(n_1342),
.A2(n_1316),
.A3(n_1327),
.B1(n_1311),
.B2(n_1321),
.C1(n_1307),
.C2(n_1310),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1343),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1335),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1339),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1344),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1345),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1352),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1349),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1350),
.A2(n_1338),
.B1(n_1342),
.B2(n_1341),
.C(n_1337),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1352),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1348),
.A2(n_1335),
.B1(n_1336),
.B2(n_1340),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1355),
.A2(n_1347),
.B(n_1348),
.C(n_1357),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1356),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1354),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1353),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1358),
.B(n_1351),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1360),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1360),
.B(n_1351),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1361),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1359),
.B(n_1328),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1363),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1364),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1362),
.Y(n_1369)
);

NOR2xp67_ASAP7_75t_L g1370 ( 
.A(n_1366),
.B(n_1346),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1365),
.B(n_1301),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1367),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1369),
.B(n_1299),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1369),
.Y(n_1374)
);

AND4x1_ASAP7_75t_L g1375 ( 
.A(n_1368),
.B(n_1371),
.C(n_1370),
.D(n_1287),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1374),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1373),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1372),
.B(n_1297),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1375),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1374),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1374),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1381),
.A2(n_1302),
.B1(n_1278),
.B2(n_1277),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1379),
.A2(n_1290),
.B1(n_1269),
.B2(n_294),
.Y(n_1383)
);

AOI31xp33_ASAP7_75t_L g1384 ( 
.A1(n_1380),
.A2(n_290),
.A3(n_292),
.B(n_295),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1377),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1385),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1384),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1382),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1386),
.A2(n_1378),
.B1(n_1376),
.B2(n_1383),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1387),
.A2(n_337),
.B1(n_310),
.B2(n_313),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1389),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1391),
.A2(n_1388),
.B1(n_1390),
.B2(n_314),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1392),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1393),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.C(n_321),
.Y(n_1394)
);

AOI211xp5_ASAP7_75t_L g1395 ( 
.A1(n_1394),
.A2(n_323),
.B(n_326),
.C(n_331),
.Y(n_1395)
);


endmodule