module fake_jpeg_17229_n_112 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_21),
.B1(n_12),
.B2(n_20),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_26),
.C(n_27),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_48),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_34),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_28),
.B1(n_22),
.B2(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_11),
.C(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_26),
.B(n_14),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_60),
.B(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_11),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_18),
.B(n_2),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_31),
.B(n_30),
.C(n_32),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_32),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_39),
.C(n_47),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_73),
.C(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_30),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_73),
.A2(n_57),
.B(n_51),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_15),
.B(n_13),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_57),
.B(n_18),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_31),
.B1(n_13),
.B2(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_31),
.B1(n_59),
.B2(n_50),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_67),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_58),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_80),
.B(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_66),
.C(n_69),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_84),
.B1(n_85),
.B2(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_18),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_88),
.B1(n_71),
.B2(n_3),
.Y(n_98)
);

XOR2x2_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_93),
.C(n_71),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_65),
.C(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_83),
.Y(n_94)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_72),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_75),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_97),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_81),
.B1(n_72),
.B2(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_6),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_89),
.C(n_87),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_104),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_7),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_2),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_6),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_4),
.B1(n_100),
.B2(n_108),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_110),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_109),
.Y(n_112)
);


endmodule