module fake_jpeg_27109_n_309 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_32),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_23),
.B1(n_15),
.B2(n_18),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_54),
.Y(n_79)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_27),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_21),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_29),
.B1(n_14),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_29),
.B1(n_43),
.B2(n_40),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_39),
.B1(n_29),
.B2(n_34),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_43),
.B1(n_40),
.B2(n_34),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_35),
.C(n_41),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_77),
.Y(n_103)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_35),
.C(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_51),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_82),
.B1(n_95),
.B2(n_48),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_54),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_22),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_89),
.B(n_22),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_60),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_95),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_31),
.CI(n_24),
.CON(n_94),
.SN(n_94)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_71),
.B(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_24),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_35),
.B(n_10),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_81),
.B(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_100),
.Y(n_126)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_107),
.A2(n_15),
.B1(n_11),
.B2(n_21),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_22),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_86),
.B1(n_28),
.B2(n_46),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_89),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_113),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_71),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_121),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_20),
.B(n_21),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_133),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_80),
.B1(n_70),
.B2(n_69),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_120),
.B1(n_129),
.B2(n_28),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_80),
.B1(n_70),
.B2(n_69),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_24),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_30),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_30),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_19),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_52),
.B1(n_28),
.B2(n_15),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_8),
.B(n_10),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_6),
.B(n_10),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_87),
.B(n_96),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_19),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_18),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_17),
.C(n_18),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_94),
.B1(n_104),
.B2(n_99),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_137),
.A2(n_145),
.B1(n_164),
.B2(n_146),
.Y(n_188)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_156),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_6),
.B(n_7),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_101),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_144),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_102),
.B1(n_85),
.B2(n_92),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_92),
.B1(n_20),
.B2(n_85),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_149),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_91),
.B(n_86),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_163),
.B(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_155),
.Y(n_174)
);

CKINVDCx10_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_158),
.B(n_166),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_19),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_16),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_6),
.B(n_7),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_110),
.A2(n_15),
.B1(n_53),
.B2(n_46),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_19),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_170),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_17),
.C(n_11),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_12),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_119),
.B1(n_116),
.B2(n_117),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_178),
.B1(n_190),
.B2(n_199),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_113),
.B1(n_121),
.B2(n_112),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_136),
.C(n_135),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_187),
.C(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_159),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_33),
.C(n_25),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_147),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_15),
.B1(n_11),
.B2(n_16),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_165),
.C(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_143),
.A2(n_53),
.B1(n_11),
.B2(n_17),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_198),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_148),
.B(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_203),
.B(n_209),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_139),
.C(n_165),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_208),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_212),
.B1(n_184),
.B2(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_206),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_171),
.C(n_153),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_142),
.B(n_168),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_160),
.C(n_154),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_13),
.B1(n_33),
.B2(n_25),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_186),
.B1(n_181),
.B2(n_197),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_12),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_13),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_182),
.Y(n_227)
);

OA21x2_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_218),
.B(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_SL g232 ( 
.A(n_210),
.B(n_180),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_203),
.B(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_216),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_188),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_181),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_207),
.B1(n_197),
.B2(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_207),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_249),
.B1(n_252),
.B2(n_190),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_199),
.B1(n_174),
.B2(n_184),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_222),
.B1(n_200),
.B2(n_213),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_259),
.B1(n_229),
.B2(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_192),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_236),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_212),
.B(n_186),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_258),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_241),
.C(n_242),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_268),
.C(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_240),
.C(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_230),
.C(n_239),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_255),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_248),
.B1(n_227),
.B2(n_249),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_279),
.B1(n_280),
.B2(n_5),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_230),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_264),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_248),
.B1(n_33),
.B2(n_12),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_5),
.B1(n_7),
.B2(n_6),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_263),
.B(n_260),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_272),
.B(n_260),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_294),
.B(n_0),
.Y(n_298)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_12),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_289),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_5),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_292),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_33),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_293),
.A3(n_31),
.B1(n_280),
.B2(n_277),
.C1(n_279),
.C2(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_273),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_0),
.B(n_1),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_31),
.C(n_1),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_298),
.B(n_1),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_0),
.B(n_1),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_1),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_287),
.B(n_2),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.C(n_303),
.Y(n_304)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_300),
.B(n_295),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.C(n_31),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_3),
.B(n_4),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_3),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_3),
.B(n_4),
.Y(n_309)
);


endmodule