module fake_aes_4788_n_18 (n_1, n_2, n_4, n_3, n_5, n_0, n_18);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_17;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
OAI22xp5_ASAP7_75t_L g6 ( .A1(n_1), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_6) );
INVx3_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_1), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_9), .Y(n_10) );
OAI22xp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx2_ASAP7_75t_SL g14 ( .A(n_13), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_14), .B(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
endmodule