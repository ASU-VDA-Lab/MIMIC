module fake_jpeg_32116_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_3),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_13),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_22),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_14),
.B1(n_17),
.B2(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_18),
.B1(n_8),
.B2(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_36),
.B(n_37),
.Y(n_38)
);

XNOR2x2_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_15),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_10),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_31),
.B(n_25),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_26),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_26),
.B1(n_15),
.B2(n_5),
.Y(n_41)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_38),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_32),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_43),
.B1(n_2),
.B2(n_6),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_49),
.B(n_1),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_2),
.C(n_13),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_13),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);


endmodule