module fake_jpeg_8522_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_12),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_2),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_23),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_55),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_23),
.B1(n_35),
.B2(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_64),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_56),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_22),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_28),
.B(n_26),
.C(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_19),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_3),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_69),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_26),
.B1(n_19),
.B2(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_76),
.B1(n_50),
.B2(n_28),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_80),
.Y(n_114)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_87),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_31),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_93),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_32),
.B1(n_20),
.B2(n_26),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_99),
.B1(n_104),
.B2(n_90),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_34),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_95),
.B(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_96),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_2),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_48),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_28),
.B(n_29),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_26),
.B1(n_24),
.B2(n_19),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_3),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_28),
.B(n_5),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_59),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_28),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_34),
.B1(n_29),
.B2(n_5),
.Y(n_104)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_91),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_93),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_117),
.B(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_46),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_129),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_67),
.B1(n_49),
.B2(n_50),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_125),
.B1(n_134),
.B2(n_89),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_68),
.B1(n_71),
.B2(n_60),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_49),
.C(n_55),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_73),
.C(n_85),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_72),
.A3(n_71),
.B1(n_50),
.B2(n_34),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_93),
.B(n_107),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_50),
.B1(n_70),
.B2(n_29),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_95),
.B1(n_74),
.B2(n_102),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_103),
.B(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_75),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_28),
.B1(n_6),
.B2(n_9),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_16),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_4),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_142),
.B(n_127),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_156),
.B1(n_108),
.B2(n_131),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_73),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_124),
.B1(n_128),
.B2(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_139),
.C(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_85),
.B1(n_97),
.B2(n_75),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_157),
.B(n_160),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_107),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_100),
.B1(n_126),
.B2(n_132),
.C(n_129),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_189),
.B(n_149),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_165),
.B1(n_149),
.B2(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_190),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_152),
.B1(n_148),
.B2(n_150),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_184),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_108),
.C(n_126),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_145),
.C(n_160),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_100),
.C(n_80),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_158),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_154),
.C(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_163),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_192),
.C(n_195),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_201),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_142),
.B(n_155),
.C(n_166),
.D(n_143),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_179),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_161),
.B1(n_164),
.B2(n_140),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_204),
.B1(n_210),
.B2(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_213),
.B(n_216),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_146),
.B1(n_153),
.B2(n_151),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_211),
.B(n_174),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_206),
.B(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_209),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_122),
.B1(n_87),
.B2(n_83),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_R g211 ( 
.A(n_189),
.B(n_105),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_123),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_234),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_180),
.C(n_170),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_170),
.C(n_184),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_181),
.C(n_168),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_238),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_199),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_183),
.B(n_191),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_168),
.B(n_181),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_213),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_167),
.C(n_175),
.Y(n_238)
);

OAI31xp33_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_211),
.A3(n_207),
.B(n_203),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_247),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_216),
.B(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_204),
.Y(n_250)
);

AOI31xp67_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_202),
.A3(n_167),
.B(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_201),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_109),
.B1(n_81),
.B2(n_82),
.Y(n_265)
);

AOI321xp33_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_169),
.A3(n_185),
.B1(n_105),
.B2(n_10),
.C(n_11),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_238),
.B1(n_237),
.B2(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_263),
.B1(n_245),
.B2(n_6),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_265),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_226),
.C(n_236),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_264),
.C(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_248),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_235),
.B1(n_239),
.B2(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_81),
.C(n_82),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_249),
.B(n_242),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_278),
.B(n_10),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_250),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_274),
.C(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_240),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_16),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_245),
.C(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_277),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_267),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_4),
.B(n_9),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_11),
.C(n_13),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_281),
.B(n_282),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_264),
.C(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.C(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_283),
.B(n_272),
.CI(n_271),
.CON(n_288),
.SN(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_290),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_289),
.C(n_15),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_15),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_291),
.Y(n_295)
);


endmodule