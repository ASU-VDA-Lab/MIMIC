module fake_netlist_6_2234_n_1525 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1525);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1525;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1413;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1504;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_1408;
wire n_1196;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_212),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_123),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_173),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_79),
.B(n_181),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_53),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_247),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_80),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_213),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_137),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_46),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_301),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_12),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_355),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_18),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_297),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_124),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_359),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_153),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_241),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_107),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_239),
.Y(n_417)
);

CKINVDCx6p67_ASAP7_75t_R g418 ( 
.A(n_144),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_250),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_175),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_75),
.B(n_229),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_377),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_304),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_70),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_142),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_242),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_308),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_364),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_327),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_357),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_246),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_314),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_186),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_365),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_375),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_49),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_162),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_51),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_185),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_121),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_113),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_171),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_295),
.Y(n_444)
);

BUFx8_ASAP7_75t_SL g445 ( 
.A(n_202),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_248),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_107),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_252),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_183),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_249),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_362),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_149),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_141),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_138),
.Y(n_454)
);

BUFx8_ASAP7_75t_SL g455 ( 
.A(n_237),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_258),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_341),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_10),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_122),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_65),
.B(n_59),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_376),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_322),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_163),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_191),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_140),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_60),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_164),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_381),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_160),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_33),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_220),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_303),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_145),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_129),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_277),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_148),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_170),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_134),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_117),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_75),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_157),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_273),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_34),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_176),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_296),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_2),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_103),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_298),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_336),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_384),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_20),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_180),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_177),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_257),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_85),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_159),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_312),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_131),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_253),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_238),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_182),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_326),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_165),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_63),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_147),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_114),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_91),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_79),
.Y(n_508)
);

BUFx8_ASAP7_75t_SL g509 ( 
.A(n_267),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_271),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_234),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_200),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_317),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_392),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_203),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_86),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_211),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_259),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_174),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_260),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_119),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_373),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_255),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_44),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_231),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_187),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_172),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_372),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_156),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_190),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_233),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_315),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_51),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_88),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_206),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g536 ( 
.A(n_313),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_81),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_266),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_276),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_18),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_300),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_272),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_37),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_321),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_126),
.Y(n_545)
);

BUFx8_ASAP7_75t_SL g546 ( 
.A(n_154),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_192),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_60),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_76),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_47),
.B(n_299),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_113),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_179),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_47),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_29),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_112),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_284),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_8),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_58),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_61),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_351),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_11),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_374),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_268),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_281),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_150),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_24),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_136),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_31),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_235),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_59),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_42),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_240),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_388),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_209),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_523),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_570),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_477),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_553),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_410),
.B(n_0),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_416),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_400),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_570),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_495),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_570),
.Y(n_584)
);

BUFx12f_ASAP7_75t_L g585 ( 
.A(n_511),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_410),
.B(n_1),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_420),
.B(n_3),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_543),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_523),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_570),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_420),
.B(n_3),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_536),
.Y(n_594)
);

BUFx8_ASAP7_75t_L g595 ( 
.A(n_474),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_431),
.B(n_4),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_402),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_409),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_405),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_407),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_528),
.B(n_4),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

BUFx12f_ASAP7_75t_L g603 ( 
.A(n_511),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_442),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_536),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_422),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_444),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_438),
.B(n_5),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_523),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_523),
.B(n_118),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_424),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_441),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_543),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_441),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_536),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_441),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_444),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_536),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_458),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_469),
.B(n_6),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_450),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_438),
.B(n_120),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_483),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_450),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_490),
.B(n_7),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_548),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_548),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_506),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_437),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_439),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_447),
.Y(n_635)
);

NOR2x1_ASAP7_75t_L g636 ( 
.A(n_490),
.B(n_125),
.Y(n_636)
);

OAI22x1_ASAP7_75t_L g637 ( 
.A1(n_551),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_552),
.B(n_9),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_481),
.B(n_11),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_552),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_470),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_557),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_507),
.Y(n_644)
);

BUFx8_ASAP7_75t_L g645 ( 
.A(n_460),
.Y(n_645)
);

BUFx12f_ASAP7_75t_L g646 ( 
.A(n_487),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_519),
.B(n_13),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_481),
.B(n_13),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_566),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_491),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_482),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_482),
.B(n_14),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_480),
.B(n_15),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_396),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_576),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_575),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_598),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_619),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_644),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_644),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_598),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_599),
.B(n_613),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_R g664 ( 
.A(n_599),
.B(n_449),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_613),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_582),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_633),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_633),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_635),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_R g671 ( 
.A(n_650),
.B(n_465),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_650),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_R g673 ( 
.A(n_607),
.B(n_499),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_651),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_614),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_619),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_645),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_645),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_575),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_612),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_597),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_575),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_634),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_618),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_585),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_651),
.Y(n_686)
);

CKINVDCx16_ASAP7_75t_R g687 ( 
.A(n_603),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_642),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_646),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_619),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_627),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_R g692 ( 
.A(n_623),
.B(n_542),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_595),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_647),
.B(n_421),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_595),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_627),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_654),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_592),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_592),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_578),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_608),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_608),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_627),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_610),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_655),
.B(n_594),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_692),
.B(n_616),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_655),
.B(n_602),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_698),
.B(n_616),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_659),
.B(n_605),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_658),
.B(n_596),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_679),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_664),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_674),
.B(n_624),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_694),
.A2(n_601),
.B1(n_574),
.B2(n_567),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_681),
.B(n_683),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_686),
.B(n_624),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_699),
.A2(n_653),
.B1(n_577),
.B2(n_550),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_701),
.B(n_641),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_656),
.B(n_590),
.Y(n_719)
);

AND2x6_ASAP7_75t_SL g720 ( 
.A(n_700),
.B(n_399),
.Y(n_720)
);

AO221x1_ASAP7_75t_L g721 ( 
.A1(n_690),
.A2(n_637),
.B1(n_649),
.B2(n_419),
.C(n_423),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_702),
.B(n_641),
.Y(n_722)
);

NOR3xp33_ASAP7_75t_L g723 ( 
.A(n_665),
.B(n_586),
.C(n_579),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_656),
.B(n_590),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_663),
.B(n_580),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_658),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_697),
.B(n_580),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_667),
.B(n_586),
.C(n_579),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_682),
.B(n_590),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_668),
.B(n_593),
.C(n_587),
.Y(n_730)
);

INVxp33_ASAP7_75t_L g731 ( 
.A(n_671),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_670),
.B(n_630),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_676),
.B(n_587),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_659),
.B(n_606),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_672),
.B(n_596),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_676),
.B(n_593),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_703),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_679),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_666),
.B(n_611),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_704),
.B(n_628),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_704),
.B(n_628),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_669),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_691),
.B(n_638),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_703),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_696),
.B(n_583),
.Y(n_745)
);

AO221x1_ASAP7_75t_L g746 ( 
.A1(n_693),
.A2(n_427),
.B1(n_432),
.B2(n_406),
.C(n_397),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_680),
.Y(n_747)
);

OR2x2_ASAP7_75t_SL g748 ( 
.A(n_687),
.B(n_609),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_688),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_673),
.B(n_610),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_675),
.B(n_630),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_684),
.B(n_609),
.Y(n_752)
);

INVx8_ASAP7_75t_L g753 ( 
.A(n_689),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_685),
.B(n_648),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_695),
.B(n_512),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_657),
.B(n_583),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_662),
.B(n_522),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_677),
.B(n_532),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_660),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_678),
.B(n_556),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_661),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_658),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_694),
.A2(n_652),
.B(n_640),
.C(n_620),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_694),
.B(n_652),
.C(n_640),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_655),
.B(n_617),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_656),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_655),
.B(n_625),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_655),
.B(n_625),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_705),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_753),
.B(n_588),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_742),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_744),
.Y(n_773)
);

AND2x6_ASAP7_75t_SL g774 ( 
.A(n_758),
.B(n_600),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_723),
.B(n_398),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_728),
.A2(n_636),
.B1(n_403),
.B2(n_404),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_711),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_745),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_710),
.B(n_604),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_744),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_727),
.B(n_581),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_740),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_SL g783 ( 
.A(n_735),
.B(n_508),
.C(n_504),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_733),
.B(n_496),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_741),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_715),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_SL g787 ( 
.A(n_760),
.B(n_524),
.C(n_516),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_712),
.B(n_445),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_736),
.B(n_763),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_738),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_744),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_731),
.B(n_533),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_743),
.B(n_730),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_739),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_721),
.A2(n_625),
.B1(n_769),
.B2(n_768),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_739),
.Y(n_796)
);

INVx5_ASAP7_75t_L g797 ( 
.A(n_762),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_722),
.B(n_562),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_725),
.B(n_537),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_752),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_737),
.B(n_626),
.Y(n_801)
);

AND2x6_ASAP7_75t_SL g802 ( 
.A(n_757),
.B(n_632),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_769),
.A2(n_612),
.B1(n_563),
.B2(n_434),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_753),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_762),
.B(n_639),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_746),
.A2(n_612),
.B1(n_443),
.B2(n_454),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_705),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_751),
.B(n_588),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_714),
.B(n_540),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_707),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_756),
.Y(n_811)
);

NOR3x1_ASAP7_75t_L g812 ( 
.A(n_754),
.B(n_643),
.C(n_621),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_717),
.B(n_401),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_762),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_750),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_753),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_718),
.B(n_505),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_759),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_749),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_707),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_767),
.B(n_518),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_709),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_726),
.B(n_525),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_709),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_755),
.Y(n_825)
);

NAND2x1_ASAP7_75t_L g826 ( 
.A(n_747),
.B(n_527),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_734),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_706),
.B(n_408),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_708),
.B(n_622),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_748),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_734),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_766),
.B(n_544),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_713),
.A2(n_412),
.B1(n_413),
.B2(n_411),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_766),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_716),
.B(n_547),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_761),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_720),
.B(n_549),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_719),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_724),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_729),
.B(n_564),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_744),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_765),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_764),
.A2(n_573),
.B(n_565),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_742),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_744),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_742),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_742),
.Y(n_847)
);

AO22x1_ASAP7_75t_L g848 ( 
.A1(n_723),
.A2(n_555),
.B1(n_558),
.B2(n_554),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_742),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_742),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_725),
.B(n_589),
.Y(n_851)
);

OAI22xp33_ASAP7_75t_L g852 ( 
.A1(n_714),
.A2(n_418),
.B1(n_561),
.B2(n_559),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_726),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_740),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_733),
.B(n_414),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_733),
.B(n_415),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_710),
.B(n_615),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_764),
.A2(n_425),
.B1(n_426),
.B2(n_417),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_763),
.A2(n_429),
.B(n_430),
.C(n_428),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_725),
.B(n_631),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_732),
.B(n_433),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_710),
.B(n_629),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_744),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_733),
.B(n_435),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_765),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_733),
.B(n_436),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_732),
.B(n_440),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_732),
.B(n_446),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_SL g869 ( 
.A(n_727),
.B(n_571),
.C(n_568),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_737),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_800),
.B(n_455),
.Y(n_871)
);

AO32x2_ASAP7_75t_L g872 ( 
.A1(n_858),
.A2(n_19),
.A3(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_870),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_809),
.B(n_451),
.C(n_448),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_794),
.B(n_452),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_SL g876 ( 
.A1(n_781),
.A2(n_456),
.B1(n_457),
.B2(n_453),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_824),
.A2(n_461),
.B(n_459),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_777),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_SL g879 ( 
.A(n_804),
.B(n_509),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_827),
.A2(n_463),
.B(n_462),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_790),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_770),
.A2(n_467),
.B(n_464),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_811),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_796),
.B(n_468),
.Y(n_884)
);

INVx3_ASAP7_75t_SL g885 ( 
.A(n_771),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_770),
.A2(n_472),
.B(n_471),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_851),
.B(n_473),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_865),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_786),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_782),
.A2(n_476),
.B1(n_478),
.B2(n_475),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_822),
.A2(n_484),
.B(n_479),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_825),
.B(n_546),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_816),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_789),
.A2(n_488),
.B(n_489),
.C(n_485),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_SL g895 ( 
.A1(n_843),
.A2(n_493),
.B(n_494),
.C(n_492),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_780),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_799),
.A2(n_498),
.B(n_497),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_780),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_771),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_792),
.B(n_500),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_842),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_820),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_820),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_SL g904 ( 
.A1(n_837),
.A2(n_502),
.B1(n_503),
.B2(n_501),
.Y(n_904)
);

OA22x2_ASAP7_75t_L g905 ( 
.A1(n_778),
.A2(n_572),
.B1(n_513),
.B2(n_514),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_785),
.B(n_510),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_852),
.A2(n_517),
.B(n_520),
.C(n_515),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_780),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_808),
.B(n_521),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_857),
.B(n_127),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_854),
.B(n_526),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_862),
.B(n_128),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_822),
.A2(n_530),
.B1(n_531),
.B2(n_529),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_SL g914 ( 
.A1(n_807),
.A2(n_17),
.B(n_19),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_862),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_784),
.A2(n_21),
.B(n_22),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_815),
.B(n_535),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_810),
.B(n_538),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_831),
.A2(n_541),
.B(n_545),
.C(n_539),
.Y(n_919)
);

AO32x1_ASAP7_75t_L g920 ( 
.A1(n_838),
.A2(n_23),
.A3(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_834),
.A2(n_560),
.B1(n_569),
.B2(n_132),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_SL g922 ( 
.A1(n_859),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_795),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_834),
.B(n_27),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_779),
.B(n_130),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_853),
.B(n_28),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_860),
.B(n_30),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_818),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_772),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_841),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_R g931 ( 
.A(n_788),
.B(n_133),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_841),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_855),
.A2(n_139),
.B1(n_143),
.B2(n_135),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_779),
.B(n_32),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_836),
.B(n_35),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_774),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_856),
.B(n_36),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_864),
.B(n_38),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_866),
.A2(n_151),
.B1(n_152),
.B2(n_146),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_844),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_869),
.B(n_38),
.C(n_39),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_846),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_R g944 ( 
.A(n_841),
.B(n_155),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_801),
.Y(n_945)
);

NOR2xp67_ASAP7_75t_SL g946 ( 
.A(n_797),
.B(n_773),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_847),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_849),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_850),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_801),
.Y(n_950)
);

BUFx4f_ASAP7_75t_L g951 ( 
.A(n_805),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_776),
.A2(n_798),
.B(n_832),
.C(n_839),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_823),
.B(n_791),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_813),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_954)
);

OAI21xp33_ASAP7_75t_L g955 ( 
.A1(n_787),
.A2(n_40),
.B(n_41),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_797),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_775),
.B(n_42),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_819),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_791),
.B(n_43),
.Y(n_959)
);

OAI21xp33_ASAP7_75t_L g960 ( 
.A1(n_783),
.A2(n_43),
.B(n_44),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_829),
.A2(n_45),
.B(n_46),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_840),
.A2(n_49),
.B(n_45),
.C(n_48),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_797),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_803),
.A2(n_161),
.B(n_158),
.Y(n_964)
);

AO22x1_ASAP7_75t_L g965 ( 
.A1(n_812),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_830),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_829),
.B(n_54),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_835),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_814),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_845),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_845),
.A2(n_167),
.B1(n_168),
.B2(n_166),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_848),
.B(n_61),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_821),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_819),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_974)
);

OAI22x1_ASAP7_75t_L g975 ( 
.A1(n_802),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_817),
.B(n_66),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_828),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_833),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_863),
.B(n_169),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_863),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_861),
.B(n_69),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_867),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_982)
);

INVx3_ASAP7_75t_SL g983 ( 
.A(n_868),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_826),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_806),
.B(n_178),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_780),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_793),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_794),
.B(n_73),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_870),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_804),
.B(n_184),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_777),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_851),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_SL g993 ( 
.A1(n_781),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_993)
);

NOR2x1_ASAP7_75t_R g994 ( 
.A(n_804),
.B(n_74),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_794),
.B(n_77),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_777),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_857),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_809),
.A2(n_81),
.B1(n_78),
.B2(n_80),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_857),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_825),
.B(n_188),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_793),
.A2(n_83),
.B(n_78),
.C(n_82),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_786),
.B(n_83),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_777),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_R g1004 ( 
.A(n_804),
.B(n_189),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_800),
.B(n_84),
.Y(n_1005)
);

AND2x2_ASAP7_75t_SL g1006 ( 
.A(n_781),
.B(n_84),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_793),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_789),
.A2(n_194),
.B1(n_195),
.B2(n_193),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_L g1009 ( 
.A(n_809),
.B(n_87),
.C(n_88),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_782),
.A2(n_197),
.B1(n_198),
.B2(n_196),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_777),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_793),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_793),
.A2(n_93),
.B(n_89),
.C(n_92),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_789),
.A2(n_201),
.B(n_199),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_781),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_794),
.B(n_94),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_842),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_794),
.B(n_95),
.Y(n_1018)
);

OAI22x1_ASAP7_75t_L g1019 ( 
.A1(n_781),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_794),
.B(n_97),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_794),
.B(n_98),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_963),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_929),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_1017),
.B(n_99),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_888),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_938),
.A2(n_205),
.B(n_204),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_908),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_883),
.B(n_100),
.Y(n_1028)
);

BUFx2_ASAP7_75t_SL g1029 ( 
.A(n_908),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_1014),
.A2(n_208),
.B(n_207),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_878),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_901),
.B(n_100),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_939),
.A2(n_214),
.B(n_210),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_952),
.A2(n_216),
.B(n_215),
.Y(n_1034)
);

AOI22x1_ASAP7_75t_L g1035 ( 
.A1(n_973),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_943),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_881),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_924),
.A2(n_218),
.B(n_217),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_992),
.B(n_887),
.Y(n_1039)
);

AOI22x1_ASAP7_75t_L g1040 ( 
.A1(n_1019),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_900),
.B(n_104),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_928),
.Y(n_1042)
);

AO22x1_ASAP7_75t_L g1043 ( 
.A1(n_957),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_915),
.B(n_219),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_966),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_889),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

BUFx2_ASAP7_75t_SL g1048 ( 
.A(n_908),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_873),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_989),
.Y(n_1050)
);

INVx3_ASAP7_75t_SL g1051 ( 
.A(n_893),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_936),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1006),
.B(n_950),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_871),
.B(n_105),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_967),
.B(n_106),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_948),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_1002),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_894),
.A2(n_222),
.B(n_221),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_885),
.Y(n_1059)
);

BUFx10_ASAP7_75t_L g1060 ( 
.A(n_892),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_988),
.A2(n_224),
.B(n_223),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_963),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_902),
.B(n_108),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_923),
.A2(n_226),
.B(n_225),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_953),
.A2(n_228),
.B(n_227),
.Y(n_1065)
);

BUFx4_ASAP7_75t_SL g1066 ( 
.A(n_958),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_991),
.Y(n_1067)
);

BUFx2_ASAP7_75t_R g1068 ( 
.A(n_937),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_986),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_876),
.A2(n_316),
.B1(n_394),
.B2(n_393),
.Y(n_1070)
);

OA21x2_ASAP7_75t_L g1071 ( 
.A1(n_995),
.A2(n_232),
.B(n_230),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_996),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_896),
.B(n_236),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_986),
.Y(n_1074)
);

AOI22x1_ASAP7_75t_L g1075 ( 
.A1(n_1003),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_934),
.B(n_109),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1011),
.Y(n_1077)
);

BUFx2_ASAP7_75t_SL g1078 ( 
.A(n_956),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_899),
.Y(n_1079)
);

INVxp67_ASAP7_75t_SL g1080 ( 
.A(n_986),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_903),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_932),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_949),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_899),
.Y(n_1084)
);

AO21x2_ASAP7_75t_L g1085 ( 
.A1(n_985),
.A2(n_244),
.B(n_243),
.Y(n_1085)
);

NAND2x1_ASAP7_75t_L g1086 ( 
.A(n_946),
.B(n_245),
.Y(n_1086)
);

CKINVDCx6p67_ASAP7_75t_R g1087 ( 
.A(n_899),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_SL g1088 ( 
.A1(n_916),
.A2(n_323),
.B(n_391),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_956),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_967),
.B(n_110),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_941),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1016),
.A2(n_325),
.B(n_390),
.Y(n_1092)
);

AO21x2_ASAP7_75t_L g1093 ( 
.A1(n_874),
.A2(n_320),
.B(n_389),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_932),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_979),
.B(n_898),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_930),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_919),
.A2(n_918),
.B(n_1018),
.Y(n_1097)
);

BUFx2_ASAP7_75t_SL g1098 ( 
.A(n_979),
.Y(n_1098)
);

BUFx2_ASAP7_75t_R g1099 ( 
.A(n_983),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_947),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_990),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_972),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_976),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_910),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_875),
.B(n_111),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_910),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_1004),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1005),
.B(n_112),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_912),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_1020),
.A2(n_1021),
.B(n_959),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_SL g1111 ( 
.A1(n_954),
.A2(n_319),
.B(n_387),
.Y(n_1111)
);

BUFx2_ASAP7_75t_R g1112 ( 
.A(n_1000),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_927),
.A2(n_318),
.B(n_386),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_931),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_912),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_997),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_906),
.B(n_114),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_SL g1118 ( 
.A1(n_977),
.A2(n_981),
.B(n_964),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_935),
.B(n_115),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_999),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_905),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_951),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_925),
.B(n_969),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_884),
.B(n_115),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_980),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_882),
.A2(n_329),
.B(n_251),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_SL g1127 ( 
.A1(n_926),
.A2(n_116),
.B1(n_254),
.B2(n_256),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_925),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_984),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_970),
.Y(n_1130)
);

BUFx4_ASAP7_75t_SL g1131 ( 
.A(n_942),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_911),
.B(n_116),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_922),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_975),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_917),
.B(n_909),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_944),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_872),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_879),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_886),
.A2(n_261),
.B(n_262),
.Y(n_1139)
);

AO21x2_ASAP7_75t_L g1140 ( 
.A1(n_895),
.A2(n_263),
.B(n_264),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_872),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_914),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_872),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_891),
.A2(n_265),
.B(n_269),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_965),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1008),
.A2(n_270),
.B(n_274),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_974),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_961),
.B(n_275),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_904),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1009),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_920),
.Y(n_1151)
);

BUFx2_ASAP7_75t_SL g1152 ( 
.A(n_971),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_933),
.A2(n_278),
.B(n_279),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_877),
.A2(n_280),
.B(n_282),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1010),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_890),
.Y(n_1156)
);

CKINVDCx6p67_ASAP7_75t_R g1157 ( 
.A(n_994),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_940),
.A2(n_921),
.B(n_907),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_982),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_897),
.A2(n_283),
.B(n_285),
.Y(n_1160)
);

CKINVDCx14_ASAP7_75t_R g1161 ( 
.A(n_913),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_920),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_960),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_955),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_978),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1015),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_880),
.B(n_993),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_962),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_998),
.A2(n_286),
.B(n_287),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_987),
.Y(n_1170)
);

BUFx2_ASAP7_75t_SL g1171 ( 
.A(n_1001),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1007),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1012),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1091),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1166),
.A2(n_1013),
.B1(n_968),
.B2(n_290),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1128),
.B(n_395),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1141),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1148),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_1178)
);

INVx6_ASAP7_75t_L g1179 ( 
.A(n_1079),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1040),
.A2(n_1143),
.B1(n_1141),
.B2(n_1169),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1031),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1100),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1074),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1101),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1031),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1042),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_SL g1187 ( 
.A(n_1084),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1141),
.A2(n_302),
.B1(n_305),
.B2(n_306),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1034),
.A2(n_309),
.B(n_310),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1148),
.A2(n_311),
.B1(n_328),
.B2(n_330),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1046),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_1025),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1037),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1045),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1053),
.B(n_331),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1047),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1082),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1089),
.B(n_1074),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1067),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1133),
.A2(n_332),
.B(n_333),
.Y(n_1200)
);

BUFx2_ASAP7_75t_R g1201 ( 
.A(n_1051),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1094),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1167),
.A2(n_334),
.B1(n_335),
.B2(n_337),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1041),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1039),
.B(n_342),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1103),
.B(n_343),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1072),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1058),
.A2(n_344),
.B(n_345),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1164),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1077),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1040),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1118),
.A2(n_349),
.B(n_350),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1077),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1023),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1143),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1030),
.A2(n_356),
.B(n_358),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1036),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1108),
.A2(n_360),
.B1(n_361),
.B2(n_363),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1094),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_SL g1220 ( 
.A1(n_1088),
.A2(n_366),
.B(n_367),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1035),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1089),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1056),
.Y(n_1223)
);

BUFx2_ASAP7_75t_R g1224 ( 
.A(n_1149),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1114),
.A2(n_371),
.B1(n_378),
.B2(n_379),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1089),
.B(n_380),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1083),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1081),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1163),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1130),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1158),
.A2(n_1146),
.B(n_1168),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_1059),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1142),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1123),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1049),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_1028),
.Y(n_1236)
);

BUFx2_ASAP7_75t_R g1237 ( 
.A(n_1052),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1063),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1109),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1168),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1150),
.A2(n_382),
.B1(n_383),
.B2(n_385),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1109),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1170),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1022),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1122),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1105),
.A2(n_1124),
.B(n_1153),
.Y(n_1246)
);

INVx8_ASAP7_75t_L g1247 ( 
.A(n_1074),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1050),
.Y(n_1248)
);

OAI21xp33_ASAP7_75t_L g1249 ( 
.A1(n_1119),
.A2(n_1117),
.B(n_1054),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1170),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_SL g1251 ( 
.A(n_1024),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1095),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1159),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1022),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1043),
.A2(n_1156),
.B1(n_1152),
.B2(n_1161),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1159),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1145),
.A2(n_1055),
.B1(n_1090),
.B2(n_1136),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1069),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1080),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1057),
.Y(n_1260)
);

OAI22x1_ASAP7_75t_L g1261 ( 
.A1(n_1147),
.A2(n_1035),
.B1(n_1075),
.B2(n_1121),
.Y(n_1261)
);

AO21x1_ASAP7_75t_L g1262 ( 
.A1(n_1026),
.A2(n_1033),
.B(n_1092),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1098),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1022),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1087),
.Y(n_1265)
);

INVxp33_ASAP7_75t_SL g1266 ( 
.A(n_1066),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1076),
.B(n_1134),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1165),
.B(n_1098),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1110),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1062),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1172),
.A2(n_1173),
.B1(n_1155),
.B2(n_1171),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1044),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1044),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1062),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1151),
.A2(n_1162),
.B(n_1154),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1062),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1155),
.A2(n_1171),
.B1(n_1127),
.B2(n_1135),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1132),
.B(n_1099),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1055),
.A2(n_1090),
.B1(n_1075),
.B2(n_1024),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1096),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1152),
.A2(n_1135),
.B1(n_1128),
.B2(n_1120),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1096),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1025),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1125),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1107),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1128),
.B(n_1106),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1116),
.A2(n_1106),
.B1(n_1104),
.B2(n_1115),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1129),
.Y(n_1288)
);

CKINVDCx6p67_ASAP7_75t_R g1289 ( 
.A(n_1157),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1027),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1115),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1065),
.A2(n_1126),
.B(n_1144),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1255),
.A2(n_1102),
.B1(n_1138),
.B2(n_1113),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1232),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1186),
.B(n_1032),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1174),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1184),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1266),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1271),
.A2(n_1112),
.B1(n_1115),
.B2(n_1138),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1262),
.A2(n_1162),
.A3(n_1151),
.B(n_1137),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1271),
.B(n_1060),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_R g1302 ( 
.A(n_1285),
.B(n_1247),
.Y(n_1302)
);

AND4x1_ASAP7_75t_L g1303 ( 
.A(n_1178),
.B(n_1070),
.C(n_1139),
.D(n_1061),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1277),
.A2(n_1281),
.B1(n_1209),
.B2(n_1255),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1196),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1192),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1247),
.B(n_1027),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1182),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1289),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1249),
.A2(n_1097),
.B1(n_1111),
.B2(n_1160),
.Y(n_1310)
);

INVxp33_ASAP7_75t_SL g1311 ( 
.A(n_1278),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1247),
.B(n_1029),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1254),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1267),
.B(n_1068),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1191),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1238),
.B(n_1209),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_R g1317 ( 
.A(n_1187),
.B(n_1029),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1181),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1233),
.B(n_1078),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1195),
.B(n_1048),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1205),
.B(n_1048),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1206),
.B(n_1078),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1236),
.B(n_1073),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1243),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1194),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1260),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1201),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1288),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_SL g1329 ( 
.A(n_1279),
.B(n_1131),
.C(n_1086),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1265),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1201),
.Y(n_1331)
);

OR2x2_ASAP7_75t_SL g1332 ( 
.A(n_1283),
.B(n_1179),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1283),
.B(n_1064),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1250),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1183),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_SL g1336 ( 
.A(n_1257),
.B(n_1093),
.C(n_1140),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1198),
.B(n_1071),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1272),
.B(n_1038),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1193),
.B(n_1199),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1273),
.B(n_1085),
.Y(n_1340)
);

CKINVDCx16_ASAP7_75t_R g1341 ( 
.A(n_1251),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_R g1342 ( 
.A(n_1222),
.B(n_1245),
.Y(n_1342)
);

CKINVDCx16_ASAP7_75t_R g1343 ( 
.A(n_1251),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1236),
.Y(n_1344)
);

CKINVDCx16_ASAP7_75t_R g1345 ( 
.A(n_1235),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1185),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1180),
.A2(n_1268),
.B1(n_1279),
.B2(n_1287),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1177),
.A2(n_1188),
.B1(n_1208),
.B2(n_1189),
.Y(n_1348)
);

NOR4xp25_ASAP7_75t_SL g1349 ( 
.A(n_1253),
.B(n_1256),
.C(n_1240),
.D(n_1263),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1292),
.A2(n_1231),
.B(n_1246),
.Y(n_1350)
);

NAND2xp33_ASAP7_75t_R g1351 ( 
.A(n_1176),
.B(n_1222),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1237),
.Y(n_1352)
);

OAI222xp33_ASAP7_75t_L g1353 ( 
.A1(n_1211),
.A2(n_1190),
.B1(n_1215),
.B2(n_1221),
.C1(n_1177),
.C2(n_1188),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1230),
.B(n_1214),
.Y(n_1354)
);

OR2x6_ASAP7_75t_L g1355 ( 
.A(n_1198),
.B(n_1183),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1211),
.A2(n_1175),
.B1(n_1208),
.B2(n_1261),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1179),
.Y(n_1357)
);

BUFx4f_ASAP7_75t_L g1358 ( 
.A(n_1254),
.Y(n_1358)
);

INVxp33_ASAP7_75t_SL g1359 ( 
.A(n_1264),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1217),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1203),
.A2(n_1218),
.B1(n_1176),
.B2(n_1204),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1284),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1254),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1225),
.B(n_1246),
.C(n_1290),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_SL g1365 ( 
.A(n_1215),
.B(n_1221),
.C(n_1241),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1274),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1276),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1244),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1223),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1237),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1227),
.B(n_1213),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1229),
.A2(n_1239),
.B1(n_1242),
.B2(n_1259),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1220),
.A2(n_1231),
.B(n_1269),
.C(n_1252),
.Y(n_1373)
);

NAND2xp33_ASAP7_75t_L g1374 ( 
.A(n_1234),
.B(n_1286),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1224),
.Y(n_1375)
);

XNOR2xp5_ASAP7_75t_L g1376 ( 
.A(n_1286),
.B(n_1248),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1244),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1258),
.A2(n_1212),
.B1(n_1210),
.B2(n_1207),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1270),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1324),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1324),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1305),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1334),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1316),
.B(n_1228),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1325),
.B(n_1354),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1300),
.B(n_1275),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1300),
.B(n_1296),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1328),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1318),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1362),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1326),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1346),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1301),
.B(n_1200),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1365),
.A2(n_1226),
.B1(n_1291),
.B2(n_1252),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1311),
.B(n_1224),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1338),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1371),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1366),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1353),
.A2(n_1282),
.B1(n_1280),
.B2(n_1270),
.C(n_1226),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1360),
.Y(n_1400)
);

BUFx4f_ASAP7_75t_L g1401 ( 
.A(n_1307),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1369),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1361),
.A2(n_1197),
.B1(n_1202),
.B2(n_1219),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1339),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1295),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1297),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1308),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1333),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1304),
.B(n_1216),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1347),
.B(n_1320),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1340),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1373),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1350),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1321),
.B(n_1348),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1310),
.B(n_1378),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1333),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1337),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1364),
.B(n_1356),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1315),
.B(n_1322),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1396),
.B(n_1345),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1404),
.B(n_1293),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1418),
.A2(n_1299),
.B1(n_1329),
.B2(n_1323),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1390),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1383),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1408),
.B(n_1337),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1414),
.B(n_1367),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1383),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1396),
.B(n_1349),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1404),
.B(n_1319),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1390),
.B(n_1344),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1387),
.B(n_1336),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1416),
.B(n_1312),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1389),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1416),
.B(n_1417),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1389),
.Y(n_1436)
);

NOR2xp67_ASAP7_75t_SL g1437 ( 
.A(n_1388),
.B(n_1341),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1418),
.A2(n_1303),
.B1(n_1370),
.B2(n_1375),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1403),
.B(n_1372),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1405),
.B(n_1368),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1414),
.B(n_1314),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1382),
.B(n_1376),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1401),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1385),
.B(n_1332),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_1379),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1363),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1391),
.B(n_1359),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1410),
.B(n_1343),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1408),
.B(n_1307),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1417),
.B(n_1355),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1430),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1434),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1432),
.B(n_1413),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1425),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1427),
.B(n_1398),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1432),
.B(n_1413),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1436),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1424),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1426),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1428),
.B(n_1386),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1450),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1445),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1431),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1440),
.B(n_1397),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1411),
.Y(n_1466)
);

AND3x2_ASAP7_75t_L g1467 ( 
.A(n_1454),
.B(n_1395),
.C(n_1448),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1453),
.B(n_1444),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1464),
.A2(n_1439),
.B1(n_1438),
.B2(n_1422),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1462),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1458),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1458),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1463),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1453),
.B(n_1420),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1462),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1452),
.Y(n_1476)
);

OA222x2_ASAP7_75t_L g1477 ( 
.A1(n_1461),
.A2(n_1425),
.B1(n_1449),
.B2(n_1412),
.C1(n_1409),
.C2(n_1393),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1429),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1457),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1460),
.Y(n_1480)
);

NAND4xp75_ASAP7_75t_L g1481 ( 
.A(n_1456),
.B(n_1439),
.C(n_1429),
.D(n_1421),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1456),
.B(n_1441),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1466),
.Y(n_1483)
);

AOI211xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1477),
.A2(n_1412),
.B(n_1450),
.C(n_1459),
.Y(n_1484)
);

OAI211xp5_ASAP7_75t_L g1485 ( 
.A1(n_1469),
.A2(n_1438),
.B(n_1422),
.C(n_1465),
.Y(n_1485)
);

OAI31xp33_ASAP7_75t_L g1486 ( 
.A1(n_1469),
.A2(n_1454),
.A3(n_1415),
.B(n_1433),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1474),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1470),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1481),
.A2(n_1351),
.B1(n_1450),
.B2(n_1433),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1468),
.A2(n_1401),
.B1(n_1449),
.B2(n_1394),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1468),
.A2(n_1401),
.B1(n_1449),
.B2(n_1443),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1489),
.A2(n_1467),
.B1(n_1478),
.B2(n_1482),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1488),
.B(n_1467),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1484),
.A2(n_1442),
.B(n_1455),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1487),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1486),
.B(n_1482),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1492),
.A2(n_1485),
.B(n_1490),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1495),
.B(n_1306),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1494),
.A2(n_1491),
.B1(n_1476),
.B2(n_1473),
.C(n_1447),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1496),
.A2(n_1443),
.B(n_1406),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1493),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1495),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1502),
.B(n_1471),
.Y(n_1503)
);

NOR3xp33_ASAP7_75t_L g1504 ( 
.A(n_1501),
.B(n_1327),
.C(n_1331),
.Y(n_1504)
);

NAND4xp25_ASAP7_75t_L g1505 ( 
.A(n_1497),
.B(n_1419),
.C(n_1388),
.D(n_1399),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1503),
.A2(n_1352),
.B(n_1499),
.Y(n_1506)
);

NOR2xp67_ASAP7_75t_L g1507 ( 
.A(n_1505),
.B(n_1500),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1506),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1508),
.A2(n_1507),
.B1(n_1504),
.B2(n_1498),
.Y(n_1509)
);

CKINVDCx14_ASAP7_75t_R g1510 ( 
.A(n_1509),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1509),
.Y(n_1511)
);

OR3x1_ASAP7_75t_L g1512 ( 
.A(n_1510),
.B(n_1437),
.C(n_1309),
.Y(n_1512)
);

XNOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1511),
.B(n_1298),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1512),
.A2(n_1294),
.B1(n_1357),
.B2(n_1330),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1513),
.Y(n_1515)
);

AO22x2_ASAP7_75t_L g1516 ( 
.A1(n_1515),
.A2(n_1335),
.B1(n_1317),
.B2(n_1475),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1514),
.A2(n_1443),
.B1(n_1449),
.B2(n_1472),
.Y(n_1517)
);

AOI222xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1517),
.A2(n_1302),
.B1(n_1342),
.B2(n_1483),
.C1(n_1480),
.C2(n_1479),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1516),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1519),
.A2(n_1358),
.B(n_1335),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1518),
.A2(n_1355),
.B(n_1374),
.C(n_1384),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1520),
.A2(n_1443),
.B1(n_1358),
.B2(n_1313),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_R g1523 ( 
.A1(n_1521),
.A2(n_1400),
.B1(n_1402),
.B2(n_1407),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1522),
.A2(n_1313),
.B1(n_1377),
.B2(n_1433),
.C(n_1392),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1524),
.A2(n_1523),
.B1(n_1313),
.B2(n_1446),
.Y(n_1525)
);


endmodule