module fake_jpeg_21266_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_25),
.B1(n_22),
.B2(n_18),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_36),
.B1(n_17),
.B2(n_22),
.Y(n_80)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_39),
.B1(n_36),
.B2(n_19),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_88),
.B1(n_18),
.B2(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_86),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_44),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_92),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_91),
.B1(n_77),
.B2(n_25),
.Y(n_132)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_64),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_104),
.B(n_85),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_64),
.B1(n_60),
.B2(n_53),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_105),
.B1(n_111),
.B2(n_112),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_35),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_70),
.B1(n_79),
.B2(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_50),
.B1(n_38),
.B2(n_35),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_50),
.B1(n_38),
.B2(n_30),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_29),
.C(n_28),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_92),
.C(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_20),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_73),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_66),
.A2(n_30),
.B1(n_32),
.B2(n_24),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_22),
.B1(n_25),
.B2(n_16),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_32),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_30),
.B1(n_89),
.B2(n_76),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_113),
.B(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_128),
.B(n_133),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_16),
.B1(n_33),
.B2(n_31),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_87),
.B1(n_71),
.B2(n_77),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_149),
.B1(n_116),
.B2(n_97),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_134),
.B1(n_140),
.B2(n_130),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_86),
.CI(n_72),
.CON(n_133),
.SN(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_69),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_74),
.C(n_29),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_142),
.C(n_115),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_85),
.B(n_73),
.C(n_74),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_17),
.B1(n_31),
.B2(n_18),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_107),
.B1(n_119),
.B2(n_95),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_158),
.B1(n_162),
.B2(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_164),
.C(n_143),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_115),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_167),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_124),
.B(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_101),
.B1(n_113),
.B2(n_116),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_168),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_101),
.C(n_96),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_97),
.B1(n_99),
.B2(n_108),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_99),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_110),
.B1(n_100),
.B2(n_102),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_171),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_109),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_177),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_102),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_184),
.C(n_198),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_186),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_178),
.B1(n_176),
.B2(n_28),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_132),
.CI(n_148),
.CON(n_188),
.SN(n_188)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_188),
.B(n_28),
.Y(n_231)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_195),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_94),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_145),
.B(n_127),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_191),
.B(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_127),
.C(n_123),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_20),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_151),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_123),
.C(n_29),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_26),
.C(n_1),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_33),
.B1(n_31),
.B2(n_16),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_158),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_28),
.B1(n_26),
.B2(n_17),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_228),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_175),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_214),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_167),
.B1(n_168),
.B2(n_163),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_160),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_198),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_153),
.B1(n_150),
.B2(n_159),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_195),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_159),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_225),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_155),
.B1(n_151),
.B2(n_177),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_206),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_205),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_203),
.C(n_191),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_238),
.C(n_241),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_197),
.B(n_181),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_179),
.C(n_181),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_179),
.C(n_194),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_209),
.C(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_243),
.C(n_247),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_187),
.C(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_188),
.C(n_189),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_253),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_225),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_189),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_229),
.B1(n_222),
.B2(n_219),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_220),
.CI(n_224),
.CON(n_256),
.SN(n_256)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_256),
.B(n_258),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_208),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_212),
.B1(n_222),
.B2(n_232),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_249),
.B1(n_252),
.B2(n_234),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_228),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_0),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_26),
.C(n_15),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_241),
.C(n_236),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_243),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_11),
.B(n_1),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_14),
.B(n_13),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_273),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_256),
.B1(n_3),
.B2(n_4),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_233),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_275),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_235),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_235),
.C(n_12),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_266),
.C(n_270),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_278),
.B1(n_261),
.B2(n_263),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_254),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_285),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_269),
.C(n_3),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_262),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_0),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_290),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_280),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_294),
.B(n_297),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_268),
.B(n_257),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_0),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_274),
.C(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_304),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_279),
.B(n_281),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_303),
.B(n_7),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_3),
.B(n_4),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_5),
.C(n_7),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_290),
.B(n_287),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_292),
.C(n_7),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_311),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_5),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_314),
.C(n_300),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_315),
.B(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_7),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_8),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_304),
.B(n_9),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_310),
.B(n_309),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_316),
.Y(n_323)
);

OAI321xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_321),
.C(n_322),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_8),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_10),
.Y(n_326)
);


endmodule