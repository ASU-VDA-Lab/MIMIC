module fake_netlist_6_2481_n_356 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_356);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_356;

wire n_326;
wire n_256;
wire n_209;
wire n_223;
wire n_278;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_168;
wire n_125;
wire n_297;
wire n_342;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_350;
wire n_142;
wire n_143;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_280;
wire n_287;
wire n_353;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_183;
wire n_338;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_352;
wire n_272;
wire n_185;
wire n_348;
wire n_293;
wire n_334;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_166;
wire n_184;
wire n_216;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_346;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx2_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_32),
.Y(n_110)
);

INVxp33_ASAP7_75t_SL g111 ( 
.A(n_40),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_15),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_29),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_28),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_26),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVxp33_ASAP7_75t_SL g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_31),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_82),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_21),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_18),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_46),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_2),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_24),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_11),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_3),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_10),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_54),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_0),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_74),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_104),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_17),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_8),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_62),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_23),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_5),
.B(n_6),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

CKINVDCx11_ASAP7_75t_R g176 ( 
.A(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2x1p5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_118),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_141),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_116),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_147),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_151),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_111),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_112),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_146),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_171),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_166),
.B1(n_125),
.B2(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_135),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

OR2x6_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_148),
.B1(n_123),
.B2(n_144),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_177),
.B(n_175),
.C(n_178),
.Y(n_215)
);

OR2x6_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_177),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_114),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_158),
.B1(n_157),
.B2(n_119),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_156),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_115),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_131),
.B1(n_121),
.B2(n_124),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_140),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_126),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_194),
.B(n_200),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_155),
.B1(n_154),
.B2(n_128),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_122),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_153),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_127),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_152),
.B1(n_150),
.B2(n_129),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_130),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_132),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_134),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_180),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_195),
.B(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_187),
.B1(n_120),
.B2(n_195),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_195),
.B(n_179),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

NAND2x1p5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_196),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_187),
.B(n_120),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_187),
.B(n_7),
.C(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_6),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_55),
.B1(n_9),
.B2(n_12),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_56),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_7),
.B1(n_14),
.B2(n_16),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_19),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_20),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_211),
.A2(n_22),
.B(n_25),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_27),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_30),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_33),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_231),
.B(n_225),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_222),
.Y(n_264)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_215),
.B(n_234),
.C(n_232),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_227),
.B1(n_235),
.B2(n_221),
.Y(n_266)
);

AO31x2_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_208),
.A3(n_230),
.B(n_36),
.Y(n_267)
);

AO31x2_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_34),
.A3(n_35),
.B(n_37),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_38),
.B(n_41),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_42),
.B(n_43),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_44),
.B(n_45),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_47),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_247),
.B(n_242),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_48),
.B(n_49),
.Y(n_274)
);

NAND2x1p5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_251),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_51),
.B(n_52),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_53),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_237),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_63),
.B(n_64),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_65),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_67),
.Y(n_281)
);

NAND3xp33_ASAP7_75t_SL g282 ( 
.A(n_254),
.B(n_69),
.C(n_71),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_243),
.B(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

AO21x2_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_258),
.B(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_246),
.B(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_240),
.B(n_239),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_72),
.B(n_73),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_271),
.B(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_291),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

AO21x2_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_282),
.B(n_270),
.Y(n_300)
);

OR2x6_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_274),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_269),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_276),
.B(n_268),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_268),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_283),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_283),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_292),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_300),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_300),
.Y(n_322)
);

NOR2x1_ASAP7_75t_R g323 ( 
.A(n_312),
.B(n_300),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_303),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_312),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_310),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_316),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_326),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_322),
.B1(n_318),
.B2(n_328),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_331),
.B(n_334),
.C(n_332),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_333),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_336),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_318),
.B1(n_327),
.B2(n_324),
.Y(n_342)
);

OAI221xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_278),
.B1(n_323),
.B2(n_78),
.C(n_80),
.Y(n_343)
);

NAND4xp25_ASAP7_75t_SL g344 ( 
.A(n_342),
.B(n_75),
.C(n_76),
.D(n_81),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_SL g345 ( 
.A(n_343),
.B(n_86),
.C(n_92),
.Y(n_345)
);

NAND5xp2_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_94),
.C(n_95),
.D(n_96),
.E(n_98),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_347),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_344),
.B(n_295),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_99),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_350),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_350),
.A2(n_295),
.B(n_328),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_102),
.Y(n_354)
);

OR2x6_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_353),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_356)
);


endmodule