module real_aes_8811_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g508 ( .A(n_1), .Y(n_508) );
INVx1_ASAP7_75t_L g160 ( .A(n_2), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_3), .A2(n_102), .B1(n_111), .B2(n_743), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_4), .A2(n_38), .B1(n_185), .B2(n_464), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g204 ( .A1(n_5), .A2(n_176), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_6), .B(n_174), .Y(n_519) );
AND2x6_ASAP7_75t_L g153 ( .A(n_7), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_8), .A2(n_258), .B(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_9), .B(n_39), .Y(n_110) );
INVx1_ASAP7_75t_L g210 ( .A(n_10), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_11), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_13), .B(n_166), .Y(n_472) );
INVx1_ASAP7_75t_L g264 ( .A(n_14), .Y(n_264) );
INVx1_ASAP7_75t_L g502 ( .A(n_15), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_16), .B(n_141), .Y(n_524) );
AO32x2_ASAP7_75t_L g491 ( .A1(n_17), .A2(n_140), .A3(n_174), .B1(n_466), .B2(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_18), .B(n_185), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_19), .B(n_181), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_20), .B(n_141), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_21), .A2(n_31), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_21), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_22), .A2(n_50), .B1(n_185), .B2(n_464), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_23), .B(n_176), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_24), .A2(n_77), .B1(n_166), .B2(n_185), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_25), .B(n_185), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_26), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_27), .A2(n_262), .B(n_263), .C(n_265), .Y(n_261) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_29), .B(n_171), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_30), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_31), .Y(n_741) );
INVx1_ASAP7_75t_L g199 ( .A(n_32), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_33), .B(n_171), .Y(n_489) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_35), .B(n_185), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_36), .B(n_171), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_37), .A2(n_153), .B(n_156), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g197 ( .A(n_40), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_41), .B(n_164), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_42), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_43), .B(n_185), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_44), .A2(n_87), .B1(n_228), .B2(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_45), .B(n_185), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_46), .B(n_185), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_47), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_48), .B(n_507), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_49), .B(n_176), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_51), .A2(n_61), .B1(n_166), .B2(n_185), .Y(n_528) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_52), .A2(n_125), .B1(n_128), .B2(n_728), .C1(n_729), .C2(n_731), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_53), .A2(n_156), .B1(n_166), .B2(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_54), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_55), .B(n_185), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_56), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_57), .B(n_185), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_58), .A2(n_184), .B(n_208), .C(n_209), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_59), .Y(n_255) );
INVx1_ASAP7_75t_L g206 ( .A(n_60), .Y(n_206) );
INVx1_ASAP7_75t_L g154 ( .A(n_62), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_63), .B(n_185), .Y(n_509) );
INVx1_ASAP7_75t_L g144 ( .A(n_64), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_65), .Y(n_115) );
AO32x2_ASAP7_75t_L g461 ( .A1(n_66), .A2(n_174), .A3(n_233), .B1(n_462), .B2(n_466), .Y(n_461) );
INVx1_ASAP7_75t_L g541 ( .A(n_67), .Y(n_541) );
INVx1_ASAP7_75t_L g484 ( .A(n_68), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_69), .A2(n_76), .B1(n_126), .B2(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_69), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_SL g180 ( .A1(n_70), .A2(n_181), .B(n_182), .C(n_184), .Y(n_180) );
INVxp67_ASAP7_75t_L g183 ( .A(n_71), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_72), .B(n_166), .Y(n_485) );
INVx1_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_74), .Y(n_202) );
INVx1_ASAP7_75t_L g248 ( .A(n_75), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_76), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_78), .A2(n_153), .B(n_156), .C(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_79), .B(n_464), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_80), .B(n_166), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_81), .B(n_161), .Y(n_224) );
INVx2_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_83), .B(n_181), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_84), .B(n_166), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_85), .A2(n_153), .B(n_156), .C(n_159), .Y(n_155) );
INVx2_ASAP7_75t_L g105 ( .A(n_86), .Y(n_105) );
OR2x2_ASAP7_75t_L g119 ( .A(n_86), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g131 ( .A(n_86), .B(n_121), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_88), .A2(n_100), .B1(n_166), .B2(n_167), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_89), .B(n_171), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_90), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_91), .A2(n_153), .B(n_156), .C(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_92), .Y(n_243) );
INVx1_ASAP7_75t_L g179 ( .A(n_93), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_94), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_95), .B(n_161), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_96), .B(n_166), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_97), .B(n_174), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_98), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_99), .A2(n_176), .B(n_177), .Y(n_175) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_103), .Y(n_744) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_109), .Y(n_103) );
OR2x2_ASAP7_75t_L g452 ( .A(n_105), .B(n_121), .Y(n_452) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_105), .B(n_120), .Y(n_733) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g121 ( .A(n_110), .B(n_122), .Y(n_121) );
AOI22x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_124), .B1(n_734), .B2(n_736), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g735 ( .A(n_115), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_116), .A2(n_737), .B(n_742), .Y(n_736) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_123), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_119), .Y(n_742) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g728 ( .A(n_125), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B1(n_450), .B2(n_453), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_129), .A2(n_133), .B1(n_454), .B2(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_132), .A2(n_133), .B1(n_738), .B2(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR4x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_339), .C(n_399), .D(n_426), .Y(n_133) );
NAND4xp25_ASAP7_75t_SL g134 ( .A(n_135), .B(n_287), .C(n_318), .D(n_335), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_212), .B(n_214), .C(n_267), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_190), .Y(n_136) );
INVx1_ASAP7_75t_L g329 ( .A(n_137), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_137), .A2(n_370), .B1(n_418), .B2(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_172), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_138), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g280 ( .A(n_138), .B(n_192), .Y(n_280) );
AND2x2_ASAP7_75t_L g322 ( .A(n_138), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_138), .B(n_213), .Y(n_334) );
INVx1_ASAP7_75t_L g374 ( .A(n_138), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_138), .B(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g302 ( .A(n_139), .B(n_192), .Y(n_302) );
INVx3_ASAP7_75t_L g306 ( .A(n_139), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_139), .B(n_364), .Y(n_363) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_168), .Y(n_139) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_140), .A2(n_193), .B(n_201), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_140), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g229 ( .A(n_140), .Y(n_229) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_142), .B(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_155), .Y(n_146) );
OAI22xp33_ASAP7_75t_L g193 ( .A1(n_148), .A2(n_186), .B1(n_194), .B2(n_200), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_148), .A2(n_248), .B(n_249), .Y(n_247) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
AND2x4_ASAP7_75t_L g176 ( .A(n_149), .B(n_153), .Y(n_176) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g507 ( .A(n_150), .Y(n_507) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx1_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx3_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_152), .Y(n_164) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVx4_ASAP7_75t_SL g186 ( .A(n_153), .Y(n_186) );
BUFx3_ASAP7_75t_L g466 ( .A(n_153), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_153), .A2(n_470), .B(n_474), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_153), .A2(n_483), .B(n_486), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_153), .A2(n_501), .B(n_505), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_153), .A2(n_513), .B(n_516), .Y(n_512) );
INVx5_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
BUFx3_ASAP7_75t_L g228 ( .A(n_157), .Y(n_228) );
INVx1_ASAP7_75t_L g464 ( .A(n_157), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_163), .C(n_165), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_SL g483 ( .A1(n_161), .A2(n_184), .B(n_484), .C(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g494 ( .A(n_161), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_161), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_161), .A2(n_538), .B(n_539), .Y(n_537) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_162), .B(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_162), .B(n_210), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_162), .A2(n_164), .B1(n_463), .B2(n_465), .Y(n_462) );
INVx2_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
INVx4_ASAP7_75t_L g239 ( .A(n_164), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_164), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_164), .A2(n_494), .B1(n_527), .B2(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_165), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_170), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_170), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_171), .A2(n_257), .B(n_266), .Y(n_256) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_171), .A2(n_469), .B(n_477), .Y(n_468) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_171), .A2(n_482), .B(n_489), .Y(n_481) );
AND2x2_ASAP7_75t_L g393 ( .A(n_172), .B(n_203), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_172), .B(n_306), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_172), .B(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g213 ( .A(n_173), .B(n_192), .Y(n_213) );
INVx1_ASAP7_75t_L g275 ( .A(n_173), .Y(n_275) );
BUFx2_ASAP7_75t_L g279 ( .A(n_173), .Y(n_279) );
AND2x2_ASAP7_75t_L g323 ( .A(n_173), .B(n_191), .Y(n_323) );
OR2x2_ASAP7_75t_L g362 ( .A(n_173), .B(n_191), .Y(n_362) );
AND2x2_ASAP7_75t_L g387 ( .A(n_173), .B(n_203), .Y(n_387) );
AND2x2_ASAP7_75t_L g446 ( .A(n_173), .B(n_276), .Y(n_446) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_187), .Y(n_173) );
INVx4_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_174), .A2(n_512), .B(n_519), .Y(n_511) );
BUFx2_ASAP7_75t_L g258 ( .A(n_176), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .C(n_186), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_178), .A2(n_186), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_178), .A2(n_186), .B(n_260), .C(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g473 ( .A(n_181), .Y(n_473) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_185), .Y(n_240) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_188), .A2(n_204), .B(n_211), .Y(n_203) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_189), .B(n_231), .Y(n_230) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_189), .B(n_466), .C(n_526), .Y(n_525) );
AO21x1_ASAP7_75t_L g572 ( .A1(n_189), .A2(n_526), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g421 ( .A(n_190), .Y(n_421) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_203), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_191), .B(n_203), .Y(n_307) );
AND2x2_ASAP7_75t_L g317 ( .A(n_191), .B(n_306), .Y(n_317) );
BUFx2_ASAP7_75t_L g328 ( .A(n_191), .Y(n_328) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g350 ( .A(n_192), .B(n_203), .Y(n_350) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_192), .Y(n_405) );
OAI22xp5_ASAP7_75t_SL g195 ( .A1(n_196), .A2(n_197), .B1(n_198), .B2(n_199), .Y(n_195) );
INVx2_ASAP7_75t_L g198 ( .A(n_196), .Y(n_198) );
INVx4_ASAP7_75t_L g262 ( .A(n_196), .Y(n_262) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_203), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_SL g276 ( .A(n_203), .Y(n_276) );
BUFx2_ASAP7_75t_L g301 ( .A(n_203), .Y(n_301) );
INVx2_ASAP7_75t_L g320 ( .A(n_203), .Y(n_320) );
AND2x2_ASAP7_75t_L g382 ( .A(n_203), .B(n_306), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_208), .A2(n_475), .B(n_476), .Y(n_474) );
O2A1O1Ixp5_ASAP7_75t_L g540 ( .A1(n_208), .A2(n_506), .B(n_541), .C(n_542), .Y(n_540) );
AOI321xp33_ASAP7_75t_L g401 ( .A1(n_212), .A2(n_402), .A3(n_403), .B1(n_404), .B2(n_406), .C(n_407), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_213), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_213), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g395 ( .A(n_213), .B(n_374), .Y(n_395) );
AND2x2_ASAP7_75t_L g428 ( .A(n_213), .B(n_320), .Y(n_428) );
INVx1_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_244), .Y(n_215) );
OR2x2_ASAP7_75t_L g330 ( .A(n_216), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_232), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g282 ( .A(n_219), .Y(n_282) );
AND2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_246), .Y(n_292) );
AND2x2_ASAP7_75t_L g297 ( .A(n_219), .B(n_272), .Y(n_297) );
INVx1_ASAP7_75t_L g314 ( .A(n_219), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_219), .B(n_295), .Y(n_333) );
AND2x2_ASAP7_75t_L g338 ( .A(n_219), .B(n_271), .Y(n_338) );
OR2x2_ASAP7_75t_L g370 ( .A(n_219), .B(n_359), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_219), .B(n_283), .Y(n_409) );
AND2x2_ASAP7_75t_L g443 ( .A(n_219), .B(n_269), .Y(n_443) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_230), .Y(n_219) );
AOI21xp5_ASAP7_75t_SL g220 ( .A1(n_221), .A2(n_222), .B(n_229), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_226), .A2(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
INVx1_ASAP7_75t_L g253 ( .A(n_229), .Y(n_253) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_229), .A2(n_500), .B(n_510), .Y(n_499) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_229), .A2(n_536), .B(n_543), .Y(n_535) );
INVx1_ASAP7_75t_L g270 ( .A(n_232), .Y(n_270) );
INVx2_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
AND2x2_ASAP7_75t_L g325 ( .A(n_232), .B(n_296), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_232), .B(n_272), .Y(n_347) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_242), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g431 ( .A(n_245), .B(n_282), .Y(n_431) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_256), .Y(n_245) );
INVx2_ASAP7_75t_L g272 ( .A(n_246), .Y(n_272) );
AND2x2_ASAP7_75t_L g425 ( .A(n_246), .B(n_285), .Y(n_425) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_253), .B(n_254), .Y(n_246) );
AND2x2_ASAP7_75t_L g271 ( .A(n_256), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
INVx1_ASAP7_75t_L g296 ( .A(n_256), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_262), .B(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_262), .A2(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g504 ( .A(n_262), .Y(n_504) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_273), .B1(n_277), .B2(n_281), .Y(n_267) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_268), .A2(n_386), .B1(n_423), .B2(n_424), .Y(n_422) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_271), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_272), .B(n_285), .Y(n_359) );
INVx1_ASAP7_75t_L g375 ( .A(n_272), .Y(n_375) );
AND2x2_ASAP7_75t_L g316 ( .A(n_274), .B(n_317), .Y(n_316) );
INVx3_ASAP7_75t_SL g355 ( .A(n_274), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_274), .B(n_280), .Y(n_432) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g441 ( .A(n_277), .Y(n_441) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_278), .B(n_374), .Y(n_416) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx3_ASAP7_75t_SL g321 ( .A(n_280), .Y(n_321) );
NAND2x1_ASAP7_75t_SL g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g342 ( .A(n_282), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g349 ( .A(n_282), .B(n_286), .Y(n_349) );
AND2x2_ASAP7_75t_L g354 ( .A(n_282), .B(n_295), .Y(n_354) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_282), .Y(n_403) );
OAI311xp33_ASAP7_75t_L g426 ( .A1(n_283), .A2(n_427), .A3(n_429), .B1(n_430), .C1(n_440), .Y(n_426) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g439 ( .A(n_284), .B(n_312), .Y(n_439) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g295 ( .A(n_285), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g343 ( .A(n_285), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g398 ( .A(n_285), .Y(n_398) );
INVx1_ASAP7_75t_L g291 ( .A(n_286), .Y(n_291) );
INVx1_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_286), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g344 ( .A(n_286), .Y(n_344) );
AOI221xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_290), .B1(n_298), .B2(n_303), .C(n_308), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_293), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx4_ASAP7_75t_L g312 ( .A(n_292), .Y(n_312) );
AND2x2_ASAP7_75t_L g406 ( .A(n_292), .B(n_325), .Y(n_406) );
AND2x2_ASAP7_75t_L g413 ( .A(n_292), .B(n_295), .Y(n_413) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_295), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g324 ( .A(n_297), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_300), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g449 ( .A(n_302), .B(n_393), .Y(n_449) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g434 ( .A(n_306), .B(n_362), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_307), .A2(n_400), .B(n_401), .C(n_414), .Y(n_399) );
AOI21xp33_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_313), .B(n_315), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g378 ( .A(n_312), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_313), .A2(n_408), .B1(n_409), .B2(n_410), .C(n_411), .Y(n_407) );
AND2x2_ASAP7_75t_L g384 ( .A(n_314), .B(n_325), .Y(n_384) );
AND2x2_ASAP7_75t_L g437 ( .A(n_314), .B(n_332), .Y(n_437) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_317), .B(n_355), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_324), .C(n_326), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_323), .Y(n_365) );
OR2x2_ASAP7_75t_L g408 ( .A(n_320), .B(n_362), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_321), .B(n_387), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_321), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g352 ( .A(n_322), .Y(n_352) );
INVx1_ASAP7_75t_L g418 ( .A(n_325), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_333), .B2(n_334), .Y(n_326) );
INVx1_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_328), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g404 ( .A(n_329), .B(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_332), .B(n_418), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_333), .A2(n_392), .B1(n_394), .B2(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g400 ( .A(n_336), .Y(n_400) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g442 ( .A(n_337), .B(n_437), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_338), .A2(n_372), .B1(n_375), .B2(n_376), .C1(n_379), .C2(n_380), .Y(n_371) );
NAND4xp25_ASAP7_75t_SL g339 ( .A(n_340), .B(n_360), .C(n_371), .D(n_383), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_345), .B2(n_350), .C(n_351), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_343), .B(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_345), .A2(n_415), .B1(n_417), .B2(n_419), .C(n_422), .Y(n_414) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g357 ( .A(n_349), .B(n_358), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_350), .A2(n_412), .B(n_413), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_355), .B2(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_366), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g402 ( .A(n_373), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_374), .B(n_393), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_374), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_378), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g410 ( .A(n_382), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_388), .B2(n_390), .C(n_391), .Y(n_383) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI222xp33_ASAP7_75t_L g430 ( .A1(n_393), .A2(n_431), .B1(n_432), .B2(n_433), .C1(n_435), .C2(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_397), .B(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp33_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_444), .C(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g730 ( .A(n_451), .Y(n_730) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND3x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_648), .C(n_696), .Y(n_455) );
NOR4xp25_ASAP7_75t_L g456 ( .A(n_457), .B(n_576), .C(n_621), .D(n_635), .Y(n_456) );
OAI311xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_496), .A3(n_520), .B1(n_529), .C1(n_544), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_467), .Y(n_458) );
OAI21xp33_ASAP7_75t_L g529 ( .A1(n_459), .A2(n_530), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g637 ( .A(n_459), .B(n_564), .Y(n_637) );
AND2x2_ASAP7_75t_L g694 ( .A(n_459), .B(n_580), .Y(n_694) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g587 ( .A(n_460), .B(n_490), .Y(n_587) );
AND2x2_ASAP7_75t_L g644 ( .A(n_460), .B(n_592), .Y(n_644) );
INVx1_ASAP7_75t_L g685 ( .A(n_460), .Y(n_685) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_461), .Y(n_553) );
AND2x2_ASAP7_75t_L g594 ( .A(n_461), .B(n_490), .Y(n_594) );
AND2x2_ASAP7_75t_L g598 ( .A(n_461), .B(n_491), .Y(n_598) );
INVx1_ASAP7_75t_L g610 ( .A(n_461), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_466), .A2(n_537), .B(n_540), .Y(n_536) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g531 ( .A(n_468), .B(n_490), .Y(n_531) );
INVx2_ASAP7_75t_L g565 ( .A(n_468), .Y(n_565) );
AND2x2_ASAP7_75t_L g580 ( .A(n_468), .B(n_491), .Y(n_580) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_468), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_468), .B(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g600 ( .A(n_468), .B(n_563), .Y(n_600) );
INVx1_ASAP7_75t_L g612 ( .A(n_468), .Y(n_612) );
INVx1_ASAP7_75t_L g653 ( .A(n_468), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_468), .B(n_553), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_473), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g478 ( .A(n_479), .B(n_490), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g530 ( .A(n_480), .B(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
AND2x2_ASAP7_75t_SL g611 ( .A(n_480), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g615 ( .A(n_480), .B(n_490), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_480), .B(n_610), .Y(n_673) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g563 ( .A(n_481), .Y(n_563) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_481), .Y(n_579) );
OR2x2_ASAP7_75t_L g652 ( .A(n_481), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g559 ( .A(n_491), .Y(n_559) );
AND2x2_ASAP7_75t_L g564 ( .A(n_491), .B(n_565), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_494), .A2(n_506), .B(n_508), .C(n_509), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_494), .A2(n_517), .B(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_496), .B(n_547), .Y(n_710) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g680 ( .A(n_497), .B(n_522), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_511), .Y(n_497) );
AND2x2_ASAP7_75t_L g556 ( .A(n_498), .B(n_547), .Y(n_556) );
INVx2_ASAP7_75t_L g568 ( .A(n_498), .Y(n_568) );
AND2x2_ASAP7_75t_L g602 ( .A(n_498), .B(n_550), .Y(n_602) );
AND2x2_ASAP7_75t_L g669 ( .A(n_498), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_499), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g549 ( .A(n_499), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g589 ( .A(n_499), .B(n_511), .Y(n_589) );
AND2x2_ASAP7_75t_L g606 ( .A(n_499), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g532 ( .A(n_511), .B(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g550 ( .A(n_511), .Y(n_550) );
AND2x2_ASAP7_75t_L g555 ( .A(n_511), .B(n_535), .Y(n_555) );
AND2x2_ASAP7_75t_L g628 ( .A(n_511), .B(n_607), .Y(n_628) );
AND2x2_ASAP7_75t_L g693 ( .A(n_511), .B(n_683), .Y(n_693) );
OAI311xp33_ASAP7_75t_L g576 ( .A1(n_520), .A2(n_577), .A3(n_581), .B1(n_583), .C1(n_603), .Y(n_576) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g588 ( .A(n_521), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g647 ( .A(n_521), .B(n_555), .Y(n_647) );
AND2x2_ASAP7_75t_L g721 ( .A(n_521), .B(n_602), .Y(n_721) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_522), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g656 ( .A(n_522), .Y(n_656) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g547 ( .A(n_523), .Y(n_547) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_523), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g676 ( .A(n_523), .B(n_550), .Y(n_676) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
AND2x2_ASAP7_75t_L g551 ( .A(n_531), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g604 ( .A(n_531), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g684 ( .A(n_531), .B(n_685), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_532), .A2(n_564), .B1(n_584), .B2(n_588), .C(n_590), .Y(n_583) );
INVx1_ASAP7_75t_L g708 ( .A(n_533), .Y(n_708) );
OR2x2_ASAP7_75t_L g674 ( .A(n_534), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g569 ( .A(n_535), .B(n_550), .Y(n_569) );
OR2x2_ASAP7_75t_L g571 ( .A(n_535), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g596 ( .A(n_535), .Y(n_596) );
INVx2_ASAP7_75t_L g607 ( .A(n_535), .Y(n_607) );
AND2x2_ASAP7_75t_L g634 ( .A(n_535), .B(n_572), .Y(n_634) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_535), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_551), .B1(n_554), .B2(n_557), .C(n_560), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g645 ( .A(n_547), .B(n_555), .Y(n_645) );
AND2x2_ASAP7_75t_L g695 ( .A(n_547), .B(n_549), .Y(n_695) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g582 ( .A(n_549), .B(n_553), .Y(n_582) );
AND2x2_ASAP7_75t_L g661 ( .A(n_549), .B(n_634), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_550), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g620 ( .A(n_550), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_551), .A2(n_631), .B(n_633), .Y(n_630) );
OR2x2_ASAP7_75t_L g574 ( .A(n_552), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g640 ( .A(n_552), .B(n_600), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_552), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g617 ( .A(n_553), .B(n_586), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_553), .B(n_700), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_554), .B(n_580), .Y(n_690) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g613 ( .A(n_555), .B(n_568), .Y(n_613) );
INVx1_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_566), .B1(n_570), .B2(n_574), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g592 ( .A(n_563), .Y(n_592) );
INVx1_ASAP7_75t_L g605 ( .A(n_563), .Y(n_605) );
INVx1_ASAP7_75t_L g575 ( .A(n_564), .Y(n_575) );
AND2x2_ASAP7_75t_L g646 ( .A(n_564), .B(n_592), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_564), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
OR2x2_ASAP7_75t_L g570 ( .A(n_567), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_567), .B(n_683), .Y(n_682) );
NOR2xp67_ASAP7_75t_L g714 ( .A(n_567), .B(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g717 ( .A(n_569), .B(n_669), .Y(n_717) );
INVx1_ASAP7_75t_SL g683 ( .A(n_571), .Y(n_683) );
AND2x2_ASAP7_75t_L g623 ( .A(n_572), .B(n_607), .Y(n_623) );
INVx1_ASAP7_75t_L g670 ( .A(n_572), .Y(n_670) );
OAI222xp33_ASAP7_75t_L g711 ( .A1(n_577), .A2(n_667), .B1(n_712), .B2(n_713), .C1(n_716), .C2(n_718), .Y(n_711) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g632 ( .A(n_579), .Y(n_632) );
AND2x2_ASAP7_75t_L g643 ( .A(n_580), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_580), .B(n_685), .Y(n_712) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_582), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g687 ( .A(n_584), .Y(n_687) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g625 ( .A(n_587), .Y(n_625) );
AND2x2_ASAP7_75t_L g704 ( .A(n_587), .B(n_665), .Y(n_704) );
AND2x2_ASAP7_75t_L g727 ( .A(n_587), .B(n_611), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_589), .B(n_623), .Y(n_622) );
OAI32xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .A3(n_595), .B1(n_597), .B2(n_601), .Y(n_590) );
BUFx2_ASAP7_75t_L g665 ( .A(n_592), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_593), .B(n_611), .Y(n_692) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g631 ( .A(n_594), .B(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g699 ( .A(n_594), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g688 ( .A(n_595), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g659 ( .A(n_598), .B(n_632), .Y(n_659) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_600), .A2(n_622), .B1(n_624), .B2(n_626), .C(n_630), .Y(n_621) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g633 ( .A(n_602), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g639 ( .A(n_602), .B(n_623), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_608), .B2(n_613), .C(n_614), .Y(n_603) );
INVx1_ASAP7_75t_L g722 ( .A(n_604), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_605), .B(n_699), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_606), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_611), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g677 ( .A(n_611), .Y(n_677) );
BUFx3_ASAP7_75t_L g700 ( .A(n_612), .Y(n_700) );
INVx1_ASAP7_75t_SL g641 ( .A(n_613), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_613), .B(n_655), .Y(n_654) );
AOI21xp33_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_616), .B(n_618), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_615), .A2(n_716), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g662 ( .A(n_620), .B(n_623), .Y(n_662) );
INVx1_ASAP7_75t_L g726 ( .A(n_620), .Y(n_726) );
INVx2_ASAP7_75t_L g715 ( .A(n_623), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_623), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g668 ( .A(n_628), .B(n_669), .Y(n_668) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_638), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_646), .B2(n_647), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_644), .A2(n_706), .B1(n_707), .B2(n_709), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_647), .A2(n_724), .B(n_727), .Y(n_723) );
NOR4xp25_ASAP7_75t_SL g648 ( .A(n_649), .B(n_657), .C(n_666), .D(n_686), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_663), .B2(n_664), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g702 ( .A(n_662), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B1(n_674), .B2(n_677), .C(n_678), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g689 ( .A(n_669), .Y(n_689) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_681), .B(n_684), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B(n_690), .C(n_691), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_691) );
CKINVDCx14_ASAP7_75t_R g701 ( .A(n_695), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_711), .C(n_719), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B1(n_702), .B2(n_703), .C(n_705), .Y(n_697) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
CKINVDCx16_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
endmodule