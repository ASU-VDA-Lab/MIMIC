module fake_netlist_1_5798_n_30 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
INVx4_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx6_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
NAND3xp33_ASAP7_75t_SL g17 ( .A(n_12), .B(n_0), .C(n_1), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_2), .B(n_3), .Y(n_18) );
OAI21xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_16), .B(n_13), .Y(n_19) );
AO21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_13), .B(n_16), .Y(n_20) );
INVx4_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_15), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_15), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B1(n_14), .B2(n_7), .Y(n_24) );
NAND3xp33_ASAP7_75t_L g25 ( .A(n_24), .B(n_14), .C(n_5), .Y(n_25) );
AOI211xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_14), .B(n_9), .C(n_10), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
OA21x2_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_26), .B(n_4), .Y(n_30) );
endmodule