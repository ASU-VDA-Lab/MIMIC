module fake_jpeg_16313_n_148 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_47),
.B1(n_23),
.B2(n_31),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_24),
.C(n_21),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_24),
.C(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_21),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_49),
.Y(n_77)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_16),
.A2(n_11),
.B1(n_12),
.B2(n_8),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_21),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_53),
.Y(n_63)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_33),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_68),
.Y(n_87)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_20),
.B1(n_26),
.B2(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_36),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_28),
.B1(n_41),
.B2(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_42),
.B(n_19),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_71),
.C(n_80),
.Y(n_117)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_28),
.B1(n_17),
.B2(n_29),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_95),
.B(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_29),
.B1(n_9),
.B2(n_11),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_29),
.B1(n_9),
.B2(n_25),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_32),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_96),
.Y(n_107)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_118),
.B(n_97),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_67),
.C(n_73),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_62),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_98),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_66),
.C(n_55),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_84),
.B1(n_105),
.B2(n_86),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_100),
.C(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_85),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_102),
.B(n_97),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_125),
.B1(n_128),
.B2(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_130),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_92),
.B1(n_83),
.B2(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_58),
.B1(n_65),
.B2(n_55),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_131),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_133),
.B1(n_122),
.B2(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_140),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_126),
.Y(n_140)
);

OAI321xp33_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_125),
.A3(n_128),
.B1(n_127),
.B2(n_121),
.C(n_132),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

BUFx4f_ASAP7_75t_SL g142 ( 
.A(n_135),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_59),
.A3(n_71),
.B1(n_80),
.B2(n_106),
.C1(n_109),
.C2(n_145),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_143),
.Y(n_148)
);


endmodule