module fake_jpeg_2956_n_617 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_617);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_617;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_57),
.Y(n_168)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_23),
.Y(n_62)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_91),
.Y(n_139)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g98 ( 
.A(n_24),
.B(n_11),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_99),
.B(n_0),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_27),
.A2(n_37),
.B(n_55),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_22),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_109),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_28),
.Y(n_125)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_112),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_68),
.B1(n_73),
.B2(n_65),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_113),
.A2(n_128),
.B1(n_140),
.B2(n_154),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_125),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_27),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_135),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_28),
.B1(n_48),
.B2(n_49),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_134),
.A2(n_16),
.B(n_19),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_37),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_84),
.A2(n_20),
.B1(n_54),
.B2(n_49),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_85),
.A2(n_56),
.B1(n_47),
.B2(n_20),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_141),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_42),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_144),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_56),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_42),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_145),
.B(n_158),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_89),
.A2(n_55),
.B1(n_29),
.B2(n_31),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_35),
.B1(n_29),
.B2(n_31),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_94),
.A2(n_54),
.B1(n_22),
.B2(n_49),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_32),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_32),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_161),
.B(n_162),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_33),
.Y(n_162)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g283 ( 
.A(n_179),
.Y(n_283)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_181),
.Y(n_271)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_187),
.Y(n_276)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_191),
.A2(n_192),
.B1(n_214),
.B2(n_223),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_123),
.A2(n_79),
.B1(n_62),
.B2(n_69),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_156),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_193),
.B(n_212),
.Y(n_264)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_197),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_72),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_208),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_209),
.A2(n_227),
.B1(n_138),
.B2(n_30),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_78),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_210),
.B(n_216),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_113),
.A2(n_107),
.B1(n_57),
.B2(n_58),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_211),
.A2(n_230),
.B(n_232),
.C(n_34),
.Y(n_289)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_134),
.A2(n_50),
.B1(n_39),
.B2(n_108),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_146),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_215),
.B(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_147),
.B(n_50),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_217),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_152),
.B(n_100),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_218),
.B(n_234),
.Y(n_265)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_221),
.B(n_222),
.Y(n_288)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_128),
.A2(n_140),
.B1(n_154),
.B2(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_229),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_153),
.B(n_112),
.C(n_109),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_225),
.B(n_52),
.C(n_41),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_168),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_141),
.A2(n_106),
.B1(n_71),
.B2(n_83),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_115),
.B(n_105),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_233),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_130),
.B(n_30),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_236),
.Y(n_282)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_115),
.B(n_64),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_238),
.Y(n_287)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_139),
.A2(n_20),
.B1(n_22),
.B2(n_54),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_34),
.B(n_30),
.Y(n_261)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_240),
.B(n_241),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_170),
.B(n_129),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_114),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_243),
.B(n_251),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_249),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_166),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_185),
.B(n_166),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_266),
.Y(n_321)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_186),
.A2(n_129),
.B1(n_173),
.B2(n_163),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_258),
.B(n_289),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_261),
.A2(n_298),
.B(n_0),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_165),
.B1(n_175),
.B2(n_164),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_263),
.A2(n_267),
.B1(n_284),
.B2(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_183),
.B(n_176),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_191),
.A2(n_165),
.B1(n_175),
.B2(n_167),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_199),
.B(n_169),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_269),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_180),
.B(n_138),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_167),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_273),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_173),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_211),
.A2(n_138),
.B1(n_76),
.B2(n_59),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_274),
.A2(n_262),
.B1(n_292),
.B2(n_245),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_225),
.A2(n_126),
.B1(n_34),
.B2(n_163),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_209),
.B(n_133),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_291),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_202),
.B(n_133),
.Y(n_293)
);

OAI22x1_ASAP7_75t_SL g294 ( 
.A1(n_239),
.A2(n_126),
.B1(n_52),
.B2(n_41),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_296),
.B(n_203),
.Y(n_325)
);

OR2x4_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_0),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_243),
.A2(n_230),
.B1(n_238),
.B2(n_206),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_299),
.A2(n_300),
.B1(n_306),
.B2(n_307),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_229),
.B1(n_217),
.B2(n_204),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_264),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_344),
.Y(n_350)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_265),
.A2(n_179),
.B1(n_237),
.B2(n_241),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_253),
.A2(n_236),
.B1(n_201),
.B2(n_215),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_222),
.B1(n_192),
.B2(n_208),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_308),
.A2(n_323),
.B1(n_324),
.B2(n_336),
.Y(n_365)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_266),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_311),
.B(n_312),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_268),
.B(n_227),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_256),
.A2(n_182),
.B1(n_178),
.B2(n_194),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_315),
.A2(n_328),
.B(n_333),
.Y(n_376)
);

OAI21xp33_ASAP7_75t_SL g367 ( 
.A1(n_317),
.A2(n_293),
.B(n_252),
.Y(n_367)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_193),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_337),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_233),
.B1(n_196),
.B2(n_213),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_256),
.A2(n_203),
.B1(n_197),
.B2(n_52),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_325),
.B(n_276),
.C(n_286),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_254),
.A2(n_197),
.B(n_52),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_341),
.B(n_333),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_298),
.A2(n_52),
.B1(n_41),
.B2(n_3),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_329),
.A2(n_245),
.B1(n_257),
.B2(n_279),
.Y(n_388)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_330),
.Y(n_366)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_19),
.B1(n_11),
.B2(n_3),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_275),
.B1(n_292),
.B2(n_287),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_251),
.A2(n_1),
.B(n_2),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_289),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_5),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_269),
.B(n_5),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_342),
.Y(n_352)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_261),
.A2(n_6),
.B(n_8),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_277),
.B(n_6),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_343),
.A2(n_283),
.B1(n_242),
.B2(n_259),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_288),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_246),
.B(n_8),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_246),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_288),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_295),
.Y(n_372)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_296),
.B(n_9),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_279),
.C(n_271),
.Y(n_373)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_264),
.Y(n_349)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_354),
.A2(n_355),
.B1(n_359),
.B2(n_378),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_339),
.A2(n_258),
.B1(n_280),
.B2(n_244),
.Y(n_355)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_311),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_357),
.B(n_394),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_321),
.A2(n_258),
.B1(n_248),
.B2(n_247),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_363),
.A2(n_371),
.B(n_395),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_322),
.B(n_258),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_369),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_370),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_326),
.B(n_252),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_372),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_373),
.B(n_301),
.Y(n_405)
);

OAI22x1_ASAP7_75t_L g374 ( 
.A1(n_339),
.A2(n_259),
.B1(n_257),
.B2(n_283),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_374),
.A2(n_323),
.B(n_308),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_337),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_384),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_342),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_345),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_391),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_339),
.A2(n_242),
.B1(n_255),
.B2(n_250),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_386),
.A2(n_389),
.B1(n_300),
.B2(n_299),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_388),
.A2(n_315),
.B1(n_328),
.B2(n_332),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_322),
.A2(n_276),
.B1(n_271),
.B2(n_286),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_320),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_320),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_348),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_312),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_325),
.A2(n_281),
.B(n_10),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_316),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_396),
.B(n_406),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_301),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_397),
.B(n_408),
.C(n_414),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_391),
.A2(n_327),
.B1(n_316),
.B2(n_321),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_399),
.A2(n_382),
.B1(n_375),
.B2(n_366),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_363),
.A2(n_302),
.B(n_346),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_400),
.A2(n_402),
.B(n_404),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_371),
.A2(n_343),
.B(n_341),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_405),
.B(n_318),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_389),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_375),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_381),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_370),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_421),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_392),
.A2(n_327),
.B1(n_307),
.B2(n_344),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_411),
.A2(n_416),
.B1(n_418),
.B2(n_360),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_348),
.C(n_338),
.Y(n_414)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_355),
.A2(n_336),
.B1(n_306),
.B2(n_331),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_365),
.A2(n_334),
.B1(n_330),
.B2(n_303),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_383),
.B(n_347),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_422),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_381),
.B(n_305),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_423),
.B(n_352),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_349),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_428),
.C(n_433),
.Y(n_471)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_362),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_432),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_383),
.B(n_340),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_429),
.A2(n_374),
.B1(n_386),
.B2(n_385),
.Y(n_449)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_366),
.B(n_309),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_382),
.C(n_379),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_374),
.A2(n_324),
.B(n_313),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_435),
.A2(n_358),
.B(n_368),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_413),
.A2(n_369),
.B1(n_365),
.B2(n_361),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_436),
.A2(n_437),
.B1(n_450),
.B2(n_467),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_413),
.A2(n_369),
.B1(n_361),
.B2(n_387),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_438),
.A2(n_440),
.B1(n_447),
.B2(n_449),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_441),
.B(n_468),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_434),
.B(n_377),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_443),
.B(n_454),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_397),
.B(n_351),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_461),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_411),
.B1(n_418),
.B2(n_406),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_419),
.A2(n_369),
.B1(n_379),
.B2(n_384),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_402),
.A2(n_354),
.B1(n_351),
.B2(n_378),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_451),
.A2(n_459),
.B1(n_462),
.B2(n_415),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_432),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_396),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_417),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_422),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_456),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_422),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_390),
.Y(n_458)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_395),
.B(n_376),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_460),
.A2(n_469),
.B(n_435),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_405),
.B(n_407),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_412),
.A2(n_352),
.B1(n_364),
.B2(n_360),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_364),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_461),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_419),
.A2(n_376),
.B1(n_380),
.B2(n_368),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_401),
.B(n_380),
.Y(n_472)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_472),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_447),
.A2(n_410),
.B1(n_416),
.B2(n_404),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_473),
.A2(n_498),
.B1(n_446),
.B2(n_450),
.Y(n_510)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_474),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_433),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_475),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_441),
.B(n_398),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_478),
.B(n_479),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_472),
.Y(n_479)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_480),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_488),
.Y(n_505)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_439),
.Y(n_485)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_485),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_414),
.C(n_425),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_489),
.C(n_490),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_444),
.B(n_398),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_487),
.B(n_500),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_468),
.B(n_421),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_428),
.C(n_424),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_396),
.C(n_431),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_442),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_501),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_431),
.C(n_409),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_457),
.C(n_467),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_496),
.A2(n_358),
.B(n_362),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_430),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_497),
.B(n_481),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_445),
.A2(n_460),
.B(n_466),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_442),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_436),
.A2(n_446),
.B1(n_437),
.B2(n_451),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_502),
.A2(n_449),
.B1(n_466),
.B2(n_452),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_445),
.B(n_335),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_470),
.Y(n_507)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_439),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_310),
.Y(n_521)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_507),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_509),
.B(n_512),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_510),
.A2(n_515),
.B1(n_517),
.B2(n_523),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_497),
.Y(n_511)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_511),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_457),
.C(n_438),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_513),
.A2(n_532),
.B1(n_483),
.B2(n_482),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_476),
.B(n_304),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_514),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_494),
.A2(n_470),
.B1(n_465),
.B2(n_452),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_469),
.C(n_465),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_528),
.C(n_505),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_473),
.A2(n_426),
.B1(n_420),
.B2(n_403),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g519 ( 
.A(n_490),
.B(n_403),
.CI(n_427),
.CON(n_519),
.SN(n_519)
);

FAx1_ASAP7_75t_SL g551 ( 
.A(n_519),
.B(n_480),
.CI(n_488),
.CON(n_551),
.SN(n_551)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_520),
.A2(n_501),
.B(n_499),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_521),
.B(n_475),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_484),
.A2(n_362),
.B1(n_313),
.B2(n_304),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_281),
.C(n_10),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_531),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_9),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_502),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_495),
.B(n_496),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_540),
.Y(n_556)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_526),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_538),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_536),
.B(n_14),
.Y(n_573)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_519),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_548),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_512),
.B(n_489),
.C(n_493),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_544),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_530),
.C(n_509),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_524),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_545),
.B(n_546),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_508),
.B(n_499),
.C(n_477),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_483),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_547),
.B(n_549),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_516),
.B(n_477),
.C(n_482),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_551),
.A2(n_529),
.B(n_522),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_504),
.C(n_485),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_552),
.Y(n_566)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_519),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_553),
.A2(n_528),
.B(n_518),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_555),
.B(n_17),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_558),
.B(n_573),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_549),
.B(n_505),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_564),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_539),
.A2(n_522),
.B1(n_525),
.B2(n_506),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_561),
.A2(n_570),
.B1(n_571),
.B2(n_572),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_545),
.A2(n_520),
.B(n_510),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_562),
.B(n_533),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_536),
.B(n_513),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_569),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_515),
.C(n_517),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_537),
.A2(n_532),
.B1(n_521),
.B2(n_523),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_554),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_551),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_572)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_574),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_550),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_577),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_569),
.B(n_563),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_535),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_578),
.B(n_581),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_559),
.A2(n_548),
.B1(n_541),
.B2(n_551),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_564),
.B(n_542),
.C(n_546),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_583),
.C(n_588),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_560),
.B(n_552),
.C(n_543),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_534),
.Y(n_584)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_584),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_557),
.B(n_573),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_585),
.A2(n_18),
.B(n_583),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_14),
.Y(n_586)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_586),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_16),
.C(n_17),
.Y(n_588)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_589),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_581),
.A2(n_556),
.B(n_572),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_591),
.A2(n_589),
.B(n_587),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_575),
.B(n_556),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_580),
.Y(n_607)
);

OA21x2_ASAP7_75t_L g593 ( 
.A1(n_574),
.A2(n_571),
.B(n_17),
.Y(n_593)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_593),
.Y(n_602)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_600),
.Y(n_605)
);

AO21x1_ASAP7_75t_L g608 ( 
.A1(n_601),
.A2(n_603),
.B(n_606),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_599),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_595),
.B(n_582),
.Y(n_604)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_604),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_580),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_607),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_603),
.B(n_594),
.C(n_596),
.Y(n_609)
);

AOI31xp33_ASAP7_75t_L g612 ( 
.A1(n_609),
.A2(n_591),
.A3(n_590),
.B(n_602),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_612),
.A2(n_613),
.B(n_611),
.Y(n_614)
);

AOI321xp33_ASAP7_75t_L g613 ( 
.A1(n_610),
.A2(n_598),
.A3(n_605),
.B1(n_579),
.B2(n_593),
.C(n_597),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_614),
.A2(n_608),
.B(n_593),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_615),
.B(n_588),
.C(n_18),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_18),
.Y(n_617)
);


endmodule