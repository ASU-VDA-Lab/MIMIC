module fake_jpeg_20462_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_59),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_33),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_38),
.B1(n_44),
.B2(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_80),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_71),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_52),
.C(n_53),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_87),
.C(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_75),
.B1(n_81),
.B2(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_37),
.B1(n_25),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_82),
.B1(n_21),
.B2(n_20),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_25),
.B1(n_34),
.B2(n_30),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_86),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx6f_ASAP7_75t_SL g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_22),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_44),
.C(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_34),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_29),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_95),
.B1(n_21),
.B2(n_26),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_104),
.B1(n_109),
.B2(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_41),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_27),
.B(n_22),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_117),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_41),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_42),
.B1(n_29),
.B2(n_26),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_123),
.B1(n_32),
.B2(n_30),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_27),
.B1(n_89),
.B2(n_94),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_63),
.C(n_74),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_39),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_36),
.B1(n_39),
.B2(n_21),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_36),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_80),
.Y(n_130)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_131),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_154),
.B(n_83),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_24),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_45),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_103),
.B(n_83),
.C(n_31),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_137),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_36),
.B1(n_64),
.B2(n_67),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_149),
.B1(n_100),
.B2(n_115),
.Y(n_160)
);

CKINVDCx10_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_64),
.B1(n_45),
.B2(n_39),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_78),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_22),
.C(n_39),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_65),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_22),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_45),
.B1(n_16),
.B2(n_13),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_96),
.B(n_91),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_151),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_22),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_153),
.B(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_70),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_101),
.B(n_11),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_98),
.B(n_106),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_164),
.B(n_165),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_109),
.B1(n_99),
.B2(n_125),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_162),
.B1(n_178),
.B2(n_184),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_106),
.A3(n_124),
.B1(n_115),
.B2(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_31),
.B1(n_7),
.B2(n_8),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_149),
.B1(n_144),
.B2(n_131),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_107),
.B1(n_111),
.B2(n_100),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_105),
.C(n_111),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_173),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_17),
.B(n_98),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_132),
.B(n_134),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_17),
.B(n_33),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_167),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_17),
.B(n_33),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_24),
.B(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_181),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_24),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_171),
.B(n_31),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_0),
.B(n_2),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_141),
.C(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_202),
.C(n_218),
.Y(n_239)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_191),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_198),
.Y(n_236)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_154),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_143),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_204),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_151),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_16),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_16),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_16),
.B1(n_31),
.B2(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_174),
.B1(n_181),
.B2(n_169),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_0),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_178),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_14),
.B(n_12),
.C(n_10),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_186),
.B(n_179),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_220),
.B(n_232),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_186),
.B(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_173),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_201),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_165),
.B(n_161),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_176),
.C(n_166),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_235),
.C(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_192),
.Y(n_245)
);

XNOR2x2_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_234),
.B1(n_192),
.B2(n_213),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_193),
.A2(n_160),
.B(n_167),
.C(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_182),
.C(n_10),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_182),
.B1(n_7),
.B2(n_4),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_241),
.B1(n_218),
.B2(n_217),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_2),
.B(n_3),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_237),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_245),
.A2(n_262),
.B1(n_226),
.B2(n_234),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_190),
.Y(n_248)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_199),
.Y(n_278)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_194),
.C(n_209),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_237),
.C(n_235),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_225),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_260),
.Y(n_270)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_229),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_200),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_227),
.B(n_226),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_250),
.B(n_264),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_261),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_229),
.C(n_220),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_275),
.C(n_244),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_209),
.C(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_263),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_290),
.Y(n_308)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

NOR2x1_ASAP7_75t_R g293 ( 
.A(n_266),
.B(n_239),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_258),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_239),
.C(n_233),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_275),
.C(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_278),
.C(n_265),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_268),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_309),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_277),
.B(n_272),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_296),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_280),
.Y(n_309)
);

INVx11_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_311),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_271),
.B1(n_297),
.B2(n_290),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.C(n_311),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_291),
.B1(n_283),
.B2(n_294),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_276),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_317),
.B(n_281),
.C(n_286),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_304),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_323),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_303),
.C(n_309),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_316),
.A3(n_285),
.B1(n_314),
.B2(n_313),
.C1(n_310),
.C2(n_232),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_321),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_321),
.B(n_322),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_325),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_327),
.C(n_303),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_306),
.B1(n_234),
.B2(n_214),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_234),
.B(n_5),
.C(n_6),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_6),
.Y(n_334)
);


endmodule