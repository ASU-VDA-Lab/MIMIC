module fake_netlist_6_3303_n_5550 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_694, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5550);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_694;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5550;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_890;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_5534;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_5541;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_5485;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_5519;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5471;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_5508;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_3147;
wire n_2662;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_5509;
wire n_5382;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1517;
wire n_1867;
wire n_1393;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_5492;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_5499;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_5507;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3777;
wire n_3641;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5387;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5531;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_957;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4845;
wire n_4104;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_5478;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_3910;
wire n_3812;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5425;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_5454;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_5369;
wire n_975;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_5527;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_SL g699 ( 
.A(n_654),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_105),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_376),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_635),
.Y(n_703)
);

INVx4_ASAP7_75t_R g704 ( 
.A(n_551),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_219),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_332),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_91),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_346),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_362),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_559),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_265),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_634),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_114),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_149),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_670),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_42),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_596),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_178),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_377),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_99),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_555),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_138),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_552),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_636),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_604),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_656),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_441),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_280),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_564),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_540),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_221),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_452),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_71),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_245),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_337),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_59),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_233),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_202),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_691),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_214),
.Y(n_740)
);

BUFx8_ASAP7_75t_SL g741 ( 
.A(n_532),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_598),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_16),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_403),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_178),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_528),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_90),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_496),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_402),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_140),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_190),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_564),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_260),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_411),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_351),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_444),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_457),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_409),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_640),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_686),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_77),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_547),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_386),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_57),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_203),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_295),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_671),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_630),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_692),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_32),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_330),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_277),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_412),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_50),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_643),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_88),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_305),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_261),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_115),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_634),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_438),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_315),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_26),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_663),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_321),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_509),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_274),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_510),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_395),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_179),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_358),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_330),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_453),
.Y(n_793)
);

CKINVDCx14_ASAP7_75t_R g794 ( 
.A(n_17),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_463),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_602),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_135),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_519),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_626),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_281),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_70),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_262),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_400),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_641),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_57),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_515),
.Y(n_806)
);

BUFx2_ASAP7_75t_R g807 ( 
.A(n_334),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_242),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_536),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_483),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_155),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_42),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_306),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_176),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_434),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_493),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_230),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_262),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_135),
.Y(n_819)
);

CKINVDCx14_ASAP7_75t_R g820 ( 
.A(n_219),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_450),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_193),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_343),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_642),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_327),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_193),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_173),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_34),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_49),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_506),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_474),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_56),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_123),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_578),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_609),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_51),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_55),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_256),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_276),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_500),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_616),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_343),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_493),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_449),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_233),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_369),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_319),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_102),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_535),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_659),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_124),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_621),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_584),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_354),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_132),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_666),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_102),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_276),
.Y(n_858)
);

BUFx5_ASAP7_75t_L g859 ( 
.A(n_625),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_52),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_11),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_236),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_51),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_264),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_444),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_12),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_571),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_192),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_247),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_207),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_647),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_355),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_591),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_115),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_52),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_639),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_293),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_285),
.Y(n_878)
);

BUFx2_ASAP7_75t_SL g879 ( 
.A(n_652),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_26),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_453),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_501),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_175),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_461),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_575),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_423),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_131),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_100),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_388),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_129),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_667),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_198),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_309),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_625),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_397),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_185),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_103),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_176),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_88),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_32),
.Y(n_900)
);

BUFx10_ASAP7_75t_L g901 ( 
.A(n_134),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_658),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_230),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_214),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_59),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_474),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_200),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_141),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_278),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_236),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_482),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_539),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_477),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_133),
.Y(n_914)
);

BUFx10_ASAP7_75t_L g915 ( 
.A(n_323),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_370),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_490),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_469),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_357),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_384),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_426),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_36),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_431),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_383),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_523),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_187),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_147),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_516),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_30),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_673),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_619),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_690),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_296),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_352),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_452),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_638),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_117),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_237),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_82),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_484),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_235),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_608),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_400),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_660),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_558),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_92),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_561),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_17),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_528),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_247),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_251),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_156),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_255),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_694),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_356),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_675),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_510),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_393),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_661),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_317),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_556),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_38),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_305),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_286),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_415),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_525),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_332),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_231),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_669),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_111),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_311),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_527),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_514),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_436),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_295),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_384),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_172),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_177),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_482),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_425),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_563),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_118),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_131),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_194),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_585),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_614),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_608),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_218),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_284),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_40),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_696),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_216),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_620),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_337),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_592),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_392),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_45),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_110),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_479),
.Y(n_999)
);

CKINVDCx14_ASAP7_75t_R g1000 ( 
.A(n_296),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_22),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_571),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_590),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_261),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_197),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_246),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_120),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_587),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_637),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_209),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_44),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_0),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_252),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_133),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_433),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_449),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_210),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_99),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_58),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_258),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_129),
.Y(n_1021)
);

BUFx10_ASAP7_75t_L g1022 ( 
.A(n_622),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_6),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_170),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_137),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_98),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_136),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_537),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_547),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_447),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_87),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_191),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_512),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_239),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_583),
.Y(n_1035)
);

CKINVDCx14_ASAP7_75t_R g1036 ( 
.A(n_794),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_859),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_979),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_716),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_741),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_767),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_784),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_762),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_850),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_956),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_859),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_859),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_969),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_859),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_859),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_820),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_859),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1000),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_717),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_753),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_859),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_832),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_756),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_717),
.Y(n_1061)
);

INVx4_ASAP7_75t_R g1062 ( 
.A(n_745),
.Y(n_1062)
);

BUFx10_ASAP7_75t_L g1063 ( 
.A(n_703),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_771),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_726),
.Y(n_1065)
);

BUFx8_ASAP7_75t_SL g1066 ( 
.A(n_701),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_771),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_832),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_832),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_775),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_758),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_775),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_761),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_765),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_760),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_766),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_783),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_783),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_848),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_714),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_848),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_L g1082 ( 
.A(n_748),
.B(n_0),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_768),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_770),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_774),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_885),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_776),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_777),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_778),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_724),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_885),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_779),
.Y(n_1092)
);

BUFx5_ASAP7_75t_L g1093 ( 
.A(n_769),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_780),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_781),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_832),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_786),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_856),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_787),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_790),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_832),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_791),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_894),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_792),
.Y(n_1104)
);

BUFx5_ASAP7_75t_L g1105 ( 
.A(n_932),
.Y(n_1105)
);

INVxp33_ASAP7_75t_SL g1106 ( 
.A(n_817),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_888),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_796),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_798),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_799),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_894),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_965),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_800),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_965),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_801),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_802),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_881),
.B(n_1),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_803),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1025),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_804),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1025),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_899),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_809),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_951),
.Y(n_1124)
);

CKINVDCx11_ASAP7_75t_R g1125 ( 
.A(n_710),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_757),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_888),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_810),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_944),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_813),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_888),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_764),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_888),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_866),
.B(n_1),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_888),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_948),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_814),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_948),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_948),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_948),
.Y(n_1140)
);

BUFx5_ASAP7_75t_L g1141 ( 
.A(n_954),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_815),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_948),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_974),
.Y(n_1144)
);

XNOR2xp5_ASAP7_75t_L g1145 ( 
.A(n_772),
.B(n_2),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_974),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_1003),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_974),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_819),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_974),
.Y(n_1150)
);

BUFx10_ASAP7_75t_L g1151 ( 
.A(n_1020),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_823),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_974),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_976),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_824),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_976),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_808),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_710),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_976),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_976),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_825),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_827),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_829),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_831),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_833),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_834),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_836),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_976),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_891),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_818),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_702),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_838),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_713),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_839),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_727),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_730),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_700),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_732),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_733),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_737),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_840),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_720),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_738),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_740),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_959),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_742),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_844),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_746),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_891),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_845),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_750),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_751),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_752),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_849),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_755),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_851),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_991),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_759),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_857),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_715),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_858),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_763),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_700),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_891),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_860),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_861),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_865),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_867),
.Y(n_1208)
);

CKINVDCx14_ASAP7_75t_R g1209 ( 
.A(n_710),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_871),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_785),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_705),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_789),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_793),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_891),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_795),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_715),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_872),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_875),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_797),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_739),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_805),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_891),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_878),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_806),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_880),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_811),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_812),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_822),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_882),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_884),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_826),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_720),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_837),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_886),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_830),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_835),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_843),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_887),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_816),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_863),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_889),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_892),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_893),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_841),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_897),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_904),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_906),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_846),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_907),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_908),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_847),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_912),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_736),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_913),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_852),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_963),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_964),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_966),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_705),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_853),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_967),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_890),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_896),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_855),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_862),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_873),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_864),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_971),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_868),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_911),
.B(n_2),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_972),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_869),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_870),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_975),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_977),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_736),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_981),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_816),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_773),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_739),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_922),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_883),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_895),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_898),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_699),
.B(n_4),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_706),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_903),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_982),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_910),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_983),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_917),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_L g1293 ( 
.A(n_978),
.B(n_3),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_990),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_992),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_919),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_933),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_993),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_984),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_920),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_924),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_925),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_773),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_928),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_994),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_935),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_936),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_782),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_938),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_782),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_939),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_996),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_999),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1002),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_943),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_945),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_947),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_949),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_958),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_788),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1004),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_961),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1006),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_998),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_968),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_973),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1007),
.Y(n_1327)
);

BUFx8_ASAP7_75t_SL g1328 ( 
.A(n_1008),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1013),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_788),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_930),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_980),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_985),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1009),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_986),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_816),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_988),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_989),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_930),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1017),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_821),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_821),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_995),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_997),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1012),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_901),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1005),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1010),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1011),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_842),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1019),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1014),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1015),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1026),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1029),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1034),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_901),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_842),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1018),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1021),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_854),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_854),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1030),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_877),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_877),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_706),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_909),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_745),
.B(n_3),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1023),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_909),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_931),
.Y(n_1371)
);

BUFx2_ASAP7_75t_SL g1372 ( 
.A(n_902),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_901),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1035),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_879),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_931),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_915),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_955),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_707),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_955),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_707),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_970),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_708),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_708),
.Y(n_1384)
);

BUFx2_ASAP7_75t_R g1385 ( 
.A(n_709),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_709),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_970),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1016),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_711),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1016),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_915),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_711),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_876),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_915),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_876),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_712),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_987),
.Y(n_1397)
);

CKINVDCx14_ASAP7_75t_R g1398 ( 
.A(n_987),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_987),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1127),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1042),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1133),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1080),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1065),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1043),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1045),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1046),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1135),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1065),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1372),
.B(n_929),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1080),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1050),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1044),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1136),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1126),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_1200),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1138),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1139),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1099),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1098),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1100),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1140),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1102),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1126),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1143),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1104),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1108),
.B(n_929),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1144),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1132),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1132),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1146),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1148),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_1109),
.B(n_1110),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1113),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1150),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1153),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1115),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1154),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1156),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1168),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1116),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1118),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1170),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1170),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1120),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1123),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1128),
.Y(n_1447)
);

CKINVDCx16_ASAP7_75t_R g1448 ( 
.A(n_1039),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1330),
.Y(n_1449)
);

INVxp33_ASAP7_75t_SL g1450 ( 
.A(n_1053),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1159),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1130),
.B(n_653),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1234),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1159),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1075),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1234),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1059),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1137),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1142),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1159),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1209),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1059),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1068),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1068),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1203),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1069),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1069),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1149),
.B(n_1001),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1152),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1096),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1096),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1101),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1155),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1238),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1161),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1101),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1107),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1107),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1162),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1131),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1131),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1160),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1163),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1238),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1160),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1169),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1171),
.Y(n_1487)
);

CKINVDCx16_ASAP7_75t_R g1488 ( 
.A(n_1398),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1164),
.Y(n_1489)
);

CKINVDCx16_ASAP7_75t_R g1490 ( 
.A(n_1036),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1165),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1166),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1063),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1173),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1175),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1241),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1167),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1176),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1172),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1178),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1287),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1174),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1241),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1181),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1280),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1194),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1386),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1205),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1179),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1200),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1180),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1183),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_1217),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1206),
.B(n_1001),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1184),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1207),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1186),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1208),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1210),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1217),
.B(n_1022),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1263),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1219),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1224),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1226),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1188),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1191),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1192),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1263),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1230),
.B(n_712),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1193),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1221),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1221),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1195),
.Y(n_1533)
);

INVxp33_ASAP7_75t_L g1534 ( 
.A(n_1122),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1231),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1282),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1198),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1202),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1235),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1239),
.B(n_718),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1177),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1211),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1242),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1212),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1366),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1282),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1213),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1243),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1244),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1246),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1281),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1299),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1247),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1214),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1216),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1220),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1222),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1225),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1227),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1281),
.B(n_1331),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1248),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1250),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1299),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1228),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1229),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1312),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1236),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1251),
.B(n_718),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1253),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1255),
.B(n_719),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1312),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1257),
.Y(n_1572)
);

INVxp33_ASAP7_75t_SL g1573 ( 
.A(n_1053),
.Y(n_1573)
);

INVxp33_ASAP7_75t_SL g1574 ( 
.A(n_1055),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1237),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1340),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1245),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1258),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1259),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1262),
.Y(n_1580)
);

CKINVDCx16_ASAP7_75t_R g1581 ( 
.A(n_1279),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1340),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1269),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1272),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1249),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1252),
.Y(n_1586)
);

NOR2xp67_ASAP7_75t_L g1587 ( 
.A(n_1275),
.B(n_655),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1280),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1276),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1256),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1261),
.Y(n_1591)
);

INVxp33_ASAP7_75t_SL g1592 ( 
.A(n_1055),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1265),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1280),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1260),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1278),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1289),
.B(n_719),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1266),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1268),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1270),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1273),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1291),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1274),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1283),
.Y(n_1604)
);

INVxp67_ASAP7_75t_SL g1605 ( 
.A(n_1331),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1284),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1285),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1079),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1288),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1290),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1292),
.Y(n_1611)
);

CKINVDCx16_ASAP7_75t_R g1612 ( 
.A(n_1336),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1296),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1280),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1066),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1300),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1294),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1066),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1339),
.B(n_1395),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1328),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1301),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1328),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1295),
.Y(n_1623)
);

XNOR2xp5_ASAP7_75t_L g1624 ( 
.A(n_1040),
.B(n_1145),
.Y(n_1624)
);

CKINVDCx20_ASAP7_75t_R g1625 ( 
.A(n_1125),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1302),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1125),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1304),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1298),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1305),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1306),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1339),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1377),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1307),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1309),
.Y(n_1635)
);

INVxp33_ASAP7_75t_SL g1636 ( 
.A(n_1399),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1311),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1357),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1267),
.B(n_721),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1341),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1366),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1313),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1315),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1357),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1056),
.B(n_754),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1373),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1373),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1314),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1384),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1384),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1316),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1317),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1341),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1056),
.B(n_721),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1057),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1040),
.Y(n_1656)
);

BUFx10_ASAP7_75t_L g1657 ( 
.A(n_1057),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1060),
.B(n_657),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1060),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1318),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1319),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1341),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1391),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1071),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1075),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1071),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1322),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1041),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1157),
.Y(n_1669)
);

INVxp33_ASAP7_75t_SL g1670 ( 
.A(n_1073),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1124),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1232),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1325),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1326),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1332),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1333),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1335),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1337),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1073),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1074),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1338),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1074),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1076),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1343),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1076),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_1264),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1129),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1297),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1083),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1083),
.Y(n_1690)
);

CKINVDCx14_ASAP7_75t_R g1691 ( 
.A(n_1084),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1169),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1344),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1324),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1084),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1085),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1169),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1085),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1347),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1329),
.Y(n_1700)
);

NOR2xp67_ASAP7_75t_L g1701 ( 
.A(n_1087),
.B(n_662),
.Y(n_1701)
);

INVxp33_ASAP7_75t_SL g1702 ( 
.A(n_1087),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1363),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1348),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1169),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1487),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1457),
.B(n_1037),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1404),
.B(n_1061),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1486),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1505),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1457),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1486),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1494),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1633),
.B(n_1088),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1495),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1480),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1505),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1588),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1658),
.B(n_1088),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1608),
.B(n_1089),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1520),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1588),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1480),
.B(n_1047),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1404),
.B(n_1064),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1498),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1500),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1509),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1511),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1481),
.B(n_1048),
.Y(n_1729)
);

INVx6_ASAP7_75t_L g1730 ( 
.A(n_1490),
.Y(n_1730)
);

BUFx8_ASAP7_75t_L g1731 ( 
.A(n_1545),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1512),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1515),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1645),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1486),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1481),
.B(n_1049),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1594),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1701),
.B(n_1089),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1619),
.A2(n_1052),
.B(n_1051),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1486),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1462),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1409),
.B(n_1067),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1594),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1560),
.B(n_1410),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1669),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1517),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1525),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1526),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1409),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1527),
.Y(n_1750)
);

OAI22x1_ASAP7_75t_SL g1751 ( 
.A1(n_1641),
.A2(n_1106),
.B1(n_722),
.B2(n_725),
.Y(n_1751)
);

INVx6_ASAP7_75t_L g1752 ( 
.A(n_1455),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1614),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1703),
.B(n_1092),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1614),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1466),
.B(n_1054),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1455),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1467),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1451),
.A2(n_1058),
.B(n_1182),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1640),
.Y(n_1761)
);

AND2x6_ASAP7_75t_L g1762 ( 
.A(n_1427),
.B(n_1129),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1640),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1530),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1470),
.B(n_1093),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1653),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1533),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1653),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1403),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1454),
.A2(n_1233),
.B(n_1182),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1662),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1662),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1400),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1665),
.B(n_1070),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1402),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1408),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1537),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1665),
.B(n_1072),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1414),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1460),
.A2(n_1254),
.B(n_1233),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1538),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_L g1782 ( 
.A(n_1654),
.B(n_1093),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1417),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1534),
.B(n_1092),
.Y(n_1784)
);

NAND2xp33_ASAP7_75t_L g1785 ( 
.A(n_1639),
.B(n_1093),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1418),
.Y(n_1786)
);

OAI21x1_ASAP7_75t_L g1787 ( 
.A1(n_1416),
.A2(n_1277),
.B(n_1254),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1529),
.A2(n_1106),
.B1(n_1286),
.B2(n_1094),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1468),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1542),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1471),
.B(n_1093),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1547),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1422),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1472),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_SL g1795 ( 
.A(n_1461),
.B(n_1385),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1554),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1555),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1401),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1476),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1477),
.B(n_1093),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1425),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1405),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1428),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1431),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1510),
.A2(n_1303),
.B(n_1277),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1556),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1557),
.Y(n_1807)
);

BUFx8_ASAP7_75t_L g1808 ( 
.A(n_1493),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1558),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1478),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1403),
.Y(n_1811)
);

XNOR2xp5_ASAP7_75t_L g1812 ( 
.A(n_1624),
.B(n_1094),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1559),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1449),
.B(n_1095),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1687),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1687),
.B(n_1077),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1564),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1565),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1567),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1432),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1433),
.B(n_1185),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1575),
.Y(n_1822)
);

INVx5_ASAP7_75t_L g1823 ( 
.A(n_1657),
.Y(n_1823)
);

AND2x2_ASAP7_75t_SL g1824 ( 
.A(n_1514),
.B(n_1117),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1577),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1435),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1436),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1513),
.B(n_1095),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1438),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1534),
.B(n_1097),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1439),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1440),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1482),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1485),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1540),
.B(n_1097),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1568),
.B(n_1187),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1570),
.A2(n_1187),
.B1(n_1196),
.B2(n_1190),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1531),
.B(n_1078),
.Y(n_1838)
);

OA21x2_ASAP7_75t_L g1839 ( 
.A1(n_1692),
.A2(n_1308),
.B(n_1303),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1585),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1452),
.B(n_1185),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1586),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1697),
.B(n_1093),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1668),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1590),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1591),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1705),
.B(n_1093),
.Y(n_1847)
);

INVx3_ASAP7_75t_L g1848 ( 
.A(n_1593),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1704),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1597),
.B(n_1190),
.Y(n_1850)
);

AND2x6_ASAP7_75t_L g1851 ( 
.A(n_1598),
.B(n_1197),
.Y(n_1851)
);

BUFx8_ASAP7_75t_L g1852 ( 
.A(n_1493),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1488),
.B(n_1196),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1599),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1587),
.B(n_1199),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1532),
.B(n_1081),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1600),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1601),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1465),
.A2(n_1368),
.B1(n_1090),
.B2(n_1038),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1603),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1604),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1669),
.A2(n_722),
.B1(n_725),
.B2(n_723),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1606),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1607),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1406),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1671),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1609),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1407),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1551),
.B(n_1199),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1605),
.B(n_1086),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1610),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1611),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1613),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1632),
.B(n_1105),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1616),
.B(n_1105),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1621),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1626),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1628),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1412),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1631),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1634),
.Y(n_1881)
);

BUFx12f_ASAP7_75t_L g1882 ( 
.A(n_1618),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1638),
.B(n_1091),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1672),
.A2(n_723),
.B1(n_729),
.B2(n_728),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1635),
.B(n_1105),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1420),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1637),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1643),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1651),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1652),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1501),
.B(n_1201),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1660),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1421),
.B(n_1201),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1644),
.B(n_1103),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1661),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1667),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1507),
.B(n_1218),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1673),
.Y(n_1898)
);

BUFx12f_ASAP7_75t_L g1899 ( 
.A(n_1618),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1541),
.A2(n_1218),
.B1(n_1323),
.B2(n_1321),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1691),
.B(n_1321),
.Y(n_1901)
);

AND2x6_ASAP7_75t_L g1902 ( 
.A(n_1674),
.B(n_1197),
.Y(n_1902)
);

AOI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1544),
.A2(n_1327),
.B1(n_1334),
.B2(n_1323),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1675),
.Y(n_1904)
);

AND2x6_ASAP7_75t_L g1905 ( 
.A(n_1676),
.B(n_1349),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1677),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1678),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1681),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1646),
.B(n_1111),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1684),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1693),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1699),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1647),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1657),
.Y(n_1914)
);

NOR2x1_ASAP7_75t_L g1915 ( 
.A(n_1672),
.B(n_1394),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1595),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1419),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1441),
.B(n_1112),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1458),
.B(n_1114),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1483),
.B(n_1119),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1499),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1413),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1657),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1670),
.B(n_1327),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1423),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1686),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1426),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1553),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1434),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1589),
.A2(n_1345),
.B1(n_1352),
.B2(n_1334),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1695),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1437),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1442),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1445),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1446),
.B(n_1105),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1447),
.B(n_1121),
.Y(n_1936)
);

INVx3_ASAP7_75t_L g1937 ( 
.A(n_1459),
.Y(n_1937)
);

OA21x2_ASAP7_75t_L g1938 ( 
.A1(n_1469),
.A2(n_1310),
.B(n_1308),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1473),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1655),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1659),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1475),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1479),
.B(n_1105),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1489),
.Y(n_1944)
);

BUFx8_ASAP7_75t_SL g1945 ( 
.A(n_1615),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1491),
.B(n_1351),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1492),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1497),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_SL g1949 ( 
.A1(n_1686),
.A2(n_728),
.B1(n_731),
.B2(n_729),
.Y(n_1949)
);

AND2x6_ASAP7_75t_L g1950 ( 
.A(n_1450),
.B(n_1354),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1502),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1504),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1670),
.A2(n_1352),
.B1(n_1353),
.B2(n_1345),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1506),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1702),
.A2(n_900),
.B1(n_905),
.B2(n_874),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1508),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1516),
.B(n_1105),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1518),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1519),
.B(n_1355),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1522),
.B(n_1353),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1523),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1524),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1535),
.B(n_1105),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1664),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1539),
.B(n_1359),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1543),
.Y(n_1966)
);

CKINVDCx20_ASAP7_75t_R g1967 ( 
.A(n_1411),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1702),
.A2(n_1360),
.B1(n_1369),
.B2(n_1359),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1548),
.B(n_1141),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1549),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1550),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1666),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1561),
.B(n_1141),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1562),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1679),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1569),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1572),
.B(n_1360),
.Y(n_1977)
);

CKINVDCx16_ASAP7_75t_R g1978 ( 
.A(n_1448),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1680),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1578),
.A2(n_1374),
.B1(n_1369),
.B2(n_1375),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1579),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1580),
.B(n_1356),
.Y(n_1982)
);

INVxp67_ASAP7_75t_L g1983 ( 
.A(n_1682),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1683),
.A2(n_731),
.B1(n_735),
.B2(n_734),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1583),
.B(n_1374),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1584),
.Y(n_1986)
);

BUFx8_ASAP7_75t_L g1987 ( 
.A(n_1615),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1596),
.B(n_1375),
.Y(n_1988)
);

INVx5_ASAP7_75t_L g1989 ( 
.A(n_1581),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_SL g1990 ( 
.A(n_1636),
.B(n_807),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1602),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1617),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1623),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_L g1994 ( 
.A(n_1629),
.B(n_1141),
.Y(n_1994)
);

INVx6_ASAP7_75t_L g1995 ( 
.A(n_1612),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1789),
.B(n_1630),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1744),
.B(n_1642),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1714),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1770),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1770),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1873),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1770),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1873),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1780),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1745),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1935),
.B(n_1648),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1945),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1926),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1876),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1734),
.B(n_1379),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1876),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1935),
.B(n_1141),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1749),
.B(n_1358),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1844),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1887),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1780),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1887),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1780),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1734),
.B(n_1379),
.Y(n_2019)
);

CKINVDCx11_ASAP7_75t_R g2020 ( 
.A(n_1769),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1760),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1706),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1713),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1874),
.B(n_1685),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1715),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1760),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1760),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1725),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1787),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1839),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1874),
.B(n_1689),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1805),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1840),
.Y(n_2033)
);

BUFx2_ASAP7_75t_L g2034 ( 
.A(n_1844),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1839),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1839),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1945),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1824),
.B(n_1381),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1726),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1727),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1728),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1943),
.B(n_1141),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1752),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1866),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1824),
.B(n_1690),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1943),
.B(n_1696),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1732),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1711),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1711),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1733),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1716),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1716),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1746),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1840),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1752),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1753),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1749),
.B(n_1361),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_1754),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1747),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1784),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1748),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1750),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1741),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1764),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1767),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1741),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1957),
.B(n_1141),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1777),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1759),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1957),
.B(n_1141),
.Y(n_2070)
);

OA21x2_ASAP7_75t_L g2071 ( 
.A1(n_1739),
.A2(n_1320),
.B(n_1310),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1840),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1781),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1963),
.B(n_1698),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1840),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1759),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1866),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_SL g2078 ( 
.A1(n_1812),
.A2(n_1649),
.B1(n_1650),
.B2(n_1641),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1753),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1790),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1794),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_1753),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1963),
.B(n_1969),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1886),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1857),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_1830),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1789),
.B(n_1450),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1857),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1792),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_1814),
.B(n_1573),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1796),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1797),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1814),
.B(n_1573),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1838),
.B(n_1381),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1794),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1799),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_1753),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1806),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1807),
.Y(n_2099)
);

INVx3_ASAP7_75t_L g2100 ( 
.A(n_1756),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1809),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1838),
.B(n_1383),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1813),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1799),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1817),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_1913),
.A2(n_1592),
.B1(n_1574),
.B2(n_1636),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1818),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1752),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_1756),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1856),
.B(n_1383),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1756),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1857),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_1762),
.A2(n_1592),
.B1(n_1574),
.B2(n_1688),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1969),
.B(n_1389),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1857),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1856),
.B(n_1870),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1810),
.Y(n_2117)
);

HB1xp67_ASAP7_75t_L g2118 ( 
.A(n_1918),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1819),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1822),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1825),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1973),
.B(n_1389),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1845),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1846),
.Y(n_2124)
);

OA21x2_ASAP7_75t_L g2125 ( 
.A1(n_1875),
.A2(n_1342),
.B(n_1320),
.Y(n_2125)
);

INVx4_ASAP7_75t_L g2126 ( 
.A(n_1938),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_SL g2127 ( 
.A(n_1865),
.B(n_1620),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1871),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1878),
.Y(n_2129)
);

INVxp67_ASAP7_75t_L g2130 ( 
.A(n_1891),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1810),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1881),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_1918),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1870),
.B(n_1392),
.Y(n_2134)
);

BUFx2_ASAP7_75t_L g2135 ( 
.A(n_1916),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_1861),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1938),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1890),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_1758),
.B(n_1362),
.Y(n_2139)
);

OA21x2_ASAP7_75t_L g2140 ( 
.A1(n_1875),
.A2(n_1350),
.B(n_1342),
.Y(n_2140)
);

INVxp33_ASAP7_75t_SL g2141 ( 
.A(n_1795),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1919),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1973),
.B(n_1392),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1938),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1756),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1758),
.B(n_1364),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_1919),
.Y(n_2147)
);

OA21x2_ASAP7_75t_L g2148 ( 
.A1(n_1885),
.A2(n_1388),
.B(n_1350),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1710),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1763),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1892),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1861),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1895),
.Y(n_2153)
);

BUFx8_ASAP7_75t_L g2154 ( 
.A(n_1914),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_1920),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1896),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1906),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1717),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_SL g2159 ( 
.A(n_1721),
.B(n_1396),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1861),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1815),
.B(n_1365),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1883),
.B(n_1396),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1762),
.B(n_1341),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1842),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1861),
.B(n_1189),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1718),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1883),
.B(n_1397),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1849),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1889),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1858),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1889),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1864),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1872),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1722),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1763),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1737),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1889),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1894),
.B(n_1158),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1894),
.B(n_1240),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1815),
.B(n_1367),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1898),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1889),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1908),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1904),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1907),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1911),
.Y(n_2186)
);

NAND3xp33_ASAP7_75t_L g2187 ( 
.A(n_1891),
.B(n_1134),
.C(n_1082),
.Y(n_2187)
);

INVx3_ASAP7_75t_L g2188 ( 
.A(n_1763),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1768),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_1920),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1762),
.B(n_1189),
.Y(n_2191)
);

CKINVDCx8_ASAP7_75t_R g2192 ( 
.A(n_1978),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1755),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1771),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1755),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_1922),
.Y(n_2196)
);

INVxp67_ASAP7_75t_L g2197 ( 
.A(n_1897),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1772),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1848),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1762),
.B(n_1189),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1743),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1848),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1743),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1854),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1761),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1854),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1908),
.B(n_1189),
.Y(n_2207)
);

OA21x2_ASAP7_75t_L g2208 ( 
.A1(n_1885),
.A2(n_1390),
.B(n_1388),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1762),
.B(n_1204),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_1763),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1761),
.Y(n_2211)
);

INVxp67_ASAP7_75t_L g2212 ( 
.A(n_1897),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1863),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1863),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1867),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1766),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1867),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1877),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1877),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1766),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_1708),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_1931),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_1909),
.B(n_1346),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1888),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1888),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1912),
.B(n_1204),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1912),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1766),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1766),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1860),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1860),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1833),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1793),
.B(n_1801),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_1880),
.B(n_1708),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1880),
.Y(n_2235)
);

NAND2xp33_ASAP7_75t_SL g2236 ( 
.A(n_1835),
.B(n_734),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_1709),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1724),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1834),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1909),
.B(n_1393),
.Y(n_2240)
);

NOR2x1_ASAP7_75t_L g2241 ( 
.A(n_1923),
.B(n_1271),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1724),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_1742),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_1720),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1707),
.Y(n_2245)
);

AND2x6_ASAP7_75t_L g2246 ( 
.A(n_1914),
.B(n_1393),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1908),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1707),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1742),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1793),
.B(n_1204),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_1774),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1774),
.B(n_1063),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1778),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1778),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1816),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1816),
.B(n_1063),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_1908),
.B(n_1204),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1723),
.Y(n_2258)
);

OA21x2_ASAP7_75t_L g2259 ( 
.A1(n_1843),
.A2(n_1390),
.B(n_1371),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1723),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1801),
.B(n_1215),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_1836),
.B(n_1147),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1828),
.B(n_1215),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1850),
.B(n_1147),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1783),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1729),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1820),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1831),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_1946),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1729),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1832),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1757),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1828),
.B(n_1215),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1757),
.Y(n_2274)
);

BUFx2_ASAP7_75t_L g2275 ( 
.A(n_1769),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1736),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1736),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1910),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1773),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1773),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1910),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1910),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1869),
.B(n_1215),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1910),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_1709),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1869),
.B(n_1994),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1994),
.B(n_1773),
.Y(n_2287)
);

BUFx8_ASAP7_75t_L g2288 ( 
.A(n_1914),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1765),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_1811),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_1946),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_1959),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1765),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1773),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1791),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_1924),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1775),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_1709),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1775),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1791),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1775),
.B(n_1223),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1800),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1709),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1775),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1800),
.Y(n_2305)
);

INVx6_ASAP7_75t_L g2306 ( 
.A(n_1776),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_1730),
.Y(n_2307)
);

INVx4_ASAP7_75t_L g2308 ( 
.A(n_1905),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_1712),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_1712),
.Y(n_2310)
);

OA21x2_ASAP7_75t_L g2311 ( 
.A1(n_1843),
.A2(n_1847),
.B(n_1738),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1776),
.Y(n_2312)
);

HB1xp67_ASAP7_75t_L g2313 ( 
.A(n_1959),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1776),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1776),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1779),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1779),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2063),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_2307),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2027),
.Y(n_2320)
);

OR2x2_ASAP7_75t_L g2321 ( 
.A(n_2034),
.B(n_1921),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2063),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2130),
.B(n_1924),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2066),
.Y(n_2324)
);

AOI22xp33_ASAP7_75t_L g2325 ( 
.A1(n_2245),
.A2(n_1955),
.B1(n_1785),
.B2(n_1884),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2034),
.B(n_1921),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2066),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2027),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2286),
.B(n_1914),
.Y(n_2329)
);

INVx4_ASAP7_75t_L g2330 ( 
.A(n_2054),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2272),
.B(n_1958),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2285),
.Y(n_2332)
);

NOR2x1p5_ASAP7_75t_L g2333 ( 
.A(n_2307),
.B(n_1923),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2069),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2069),
.Y(n_2335)
);

BUFx10_ASAP7_75t_L g2336 ( 
.A(n_1996),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2048),
.Y(n_2337)
);

NAND3xp33_ASAP7_75t_L g2338 ( 
.A(n_2090),
.B(n_1788),
.C(n_1837),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2193),
.B(n_1950),
.Y(n_2339)
);

INVxp67_ASAP7_75t_SL g2340 ( 
.A(n_2030),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2086),
.B(n_2044),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2197),
.B(n_1977),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2048),
.Y(n_2343)
);

AO22x2_ASAP7_75t_L g2344 ( 
.A1(n_2038),
.A2(n_1955),
.B1(n_1859),
.B2(n_1984),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2076),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2033),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2005),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2076),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2212),
.B(n_2296),
.Y(n_2349)
);

INVxp67_ASAP7_75t_SL g2350 ( 
.A(n_2030),
.Y(n_2350)
);

AND2x4_ASAP7_75t_L g2351 ( 
.A(n_2043),
.B(n_2055),
.Y(n_2351)
);

INVx8_ASAP7_75t_L g2352 ( 
.A(n_2246),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2049),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2081),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2081),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2095),
.Y(n_2356)
);

NAND2xp33_ASAP7_75t_L g2357 ( 
.A(n_2246),
.B(n_1950),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2274),
.B(n_1929),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2033),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2049),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2060),
.B(n_1977),
.Y(n_2361)
);

INVx6_ASAP7_75t_L g2362 ( 
.A(n_2154),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2095),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_2087),
.B(n_1972),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2090),
.B(n_1903),
.C(n_1900),
.Y(n_2365)
);

INVx4_ASAP7_75t_L g2366 ( 
.A(n_2054),
.Y(n_2366)
);

INVxp67_ASAP7_75t_SL g2367 ( 
.A(n_2035),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2051),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2096),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2154),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2077),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2195),
.B(n_1950),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2096),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2104),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2051),
.Y(n_2375)
);

CKINVDCx16_ASAP7_75t_R g2376 ( 
.A(n_2078),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2052),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2276),
.B(n_1950),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2052),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2104),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2117),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2043),
.B(n_1823),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_2087),
.B(n_1972),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2117),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1999),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1999),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2000),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2000),
.Y(n_2388)
);

NAND3xp33_ASAP7_75t_L g2389 ( 
.A(n_2093),
.B(n_1968),
.C(n_1953),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2002),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_1998),
.B(n_1983),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2245),
.A2(n_2248),
.B1(n_2260),
.B2(n_2258),
.Y(n_2392)
);

BUFx3_ASAP7_75t_L g2393 ( 
.A(n_2154),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2006),
.B(n_1929),
.Y(n_2394)
);

AOI22xp33_ASAP7_75t_L g2395 ( 
.A1(n_2248),
.A2(n_2258),
.B1(n_2266),
.B2(n_2260),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2277),
.B(n_1950),
.Y(n_2396)
);

INVx1_ASAP7_75t_SL g2397 ( 
.A(n_2014),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2074),
.B(n_1929),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2131),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_2033),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2005),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2054),
.B(n_1929),
.Y(n_2402)
);

INVx11_ASAP7_75t_L g2403 ( 
.A(n_2288),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_2033),
.Y(n_2404)
);

INVx3_ASAP7_75t_L g2405 ( 
.A(n_2075),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2058),
.B(n_1983),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_L g2407 ( 
.A(n_2093),
.B(n_1980),
.C(n_1930),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2131),
.Y(n_2408)
);

INVxp67_ASAP7_75t_L g2409 ( 
.A(n_2178),
.Y(n_2409)
);

INVxp67_ASAP7_75t_L g2410 ( 
.A(n_2178),
.Y(n_2410)
);

NAND3xp33_ASAP7_75t_L g2411 ( 
.A(n_2010),
.B(n_1859),
.C(n_1984),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2002),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2004),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2054),
.B(n_1958),
.Y(n_2414)
);

OAI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2266),
.A2(n_1990),
.B1(n_1823),
.B2(n_1961),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2001),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2003),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2004),
.Y(n_2418)
);

BUFx2_ASAP7_75t_L g2419 ( 
.A(n_2008),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_2244),
.B(n_1865),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2016),
.Y(n_2421)
);

AOI22xp33_ASAP7_75t_L g2422 ( 
.A1(n_2270),
.A2(n_1785),
.B1(n_1862),
.B2(n_1851),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_L g2423 ( 
.A(n_2010),
.B(n_1985),
.C(n_1893),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_2054),
.B(n_1961),
.Y(n_2424)
);

INVx4_ASAP7_75t_L g2425 ( 
.A(n_2072),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2016),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_2013),
.Y(n_2427)
);

BUFx3_ASAP7_75t_L g2428 ( 
.A(n_2288),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2009),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2075),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2018),
.Y(n_2431)
);

INVx4_ASAP7_75t_L g2432 ( 
.A(n_2072),
.Y(n_2432)
);

AO22x2_ASAP7_75t_L g2433 ( 
.A1(n_2038),
.A2(n_1933),
.B1(n_1954),
.B2(n_1952),
.Y(n_2433)
);

INVx1_ASAP7_75t_SL g2434 ( 
.A(n_2008),
.Y(n_2434)
);

INVx4_ASAP7_75t_L g2435 ( 
.A(n_2072),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2018),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2222),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2270),
.B(n_1719),
.Y(n_2438)
);

OAI22xp33_ASAP7_75t_SL g2439 ( 
.A1(n_2045),
.A2(n_1738),
.B1(n_1719),
.B2(n_1855),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2026),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2026),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2026),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2011),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_2072),
.B(n_1958),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2122),
.B(n_1855),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2143),
.A2(n_1782),
.B1(n_1982),
.B2(n_1936),
.Y(n_2446)
);

CKINVDCx11_ASAP7_75t_R g2447 ( 
.A(n_2192),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2149),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2075),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2015),
.Y(n_2450)
);

INVx1_ASAP7_75t_SL g2451 ( 
.A(n_2222),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_2084),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_2086),
.B(n_1879),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2149),
.Y(n_2454)
);

AOI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2114),
.A2(n_1782),
.B1(n_1982),
.B2(n_1936),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2158),
.Y(n_2456)
);

XOR2xp5_ASAP7_75t_L g2457 ( 
.A(n_2084),
.B(n_1411),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2158),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2017),
.Y(n_2459)
);

BUFx10_ASAP7_75t_L g2460 ( 
.A(n_1996),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2019),
.B(n_1893),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2289),
.A2(n_1902),
.B1(n_1851),
.B2(n_1905),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2075),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2262),
.B(n_1988),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2022),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2023),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2072),
.B(n_1958),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2166),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2166),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2019),
.B(n_1985),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_SL g2471 ( 
.A(n_2192),
.B(n_1798),
.Y(n_2471)
);

AND2x6_ASAP7_75t_L g2472 ( 
.A(n_2137),
.B(n_1961),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_1997),
.B(n_1879),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2293),
.B(n_1821),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2112),
.B(n_1961),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2025),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_2295),
.A2(n_1902),
.B1(n_1851),
.B2(n_1905),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2288),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2028),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2174),
.Y(n_2480)
);

AOI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2114),
.A2(n_1902),
.B1(n_1851),
.B2(n_1933),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2174),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2300),
.B(n_1952),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2039),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2176),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2040),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2176),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2302),
.B(n_1954),
.Y(n_2488)
);

BUFx8_ASAP7_75t_SL g2489 ( 
.A(n_2007),
.Y(n_2489)
);

INVx4_ASAP7_75t_L g2490 ( 
.A(n_2112),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2262),
.B(n_1927),
.Y(n_2491)
);

AND2x6_ASAP7_75t_L g2492 ( 
.A(n_2137),
.B(n_1962),
.Y(n_2492)
);

INVx2_ASAP7_75t_SL g2493 ( 
.A(n_2013),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2189),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_2285),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2041),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2035),
.Y(n_2497)
);

INVx2_ASAP7_75t_SL g2498 ( 
.A(n_2013),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2055),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2047),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2036),
.Y(n_2501)
);

BUFx4f_ASAP7_75t_L g2502 ( 
.A(n_2246),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_2057),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2050),
.Y(n_2504)
);

BUFx8_ASAP7_75t_SL g2505 ( 
.A(n_2007),
.Y(n_2505)
);

INVx3_ASAP7_75t_L g2506 ( 
.A(n_2085),
.Y(n_2506)
);

BUFx2_ASAP7_75t_L g2507 ( 
.A(n_2275),
.Y(n_2507)
);

BUFx10_ASAP7_75t_L g2508 ( 
.A(n_2037),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2135),
.B(n_1986),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_2135),
.B(n_2046),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2112),
.B(n_1962),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2036),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2021),
.Y(n_2513)
);

INVxp33_ASAP7_75t_SL g2514 ( 
.A(n_2127),
.Y(n_2514)
);

INVx1_ASAP7_75t_SL g2515 ( 
.A(n_2275),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2053),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2305),
.A2(n_1902),
.B1(n_1851),
.B2(n_1905),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2059),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2057),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2083),
.B(n_2233),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2021),
.Y(n_2521)
);

OAI21xp33_ASAP7_75t_SL g2522 ( 
.A1(n_2287),
.A2(n_1966),
.B(n_1956),
.Y(n_2522)
);

INVx4_ASAP7_75t_L g2523 ( 
.A(n_2112),
.Y(n_2523)
);

OAI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2083),
.A2(n_2163),
.B1(n_2308),
.B2(n_2116),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2108),
.B(n_1823),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2264),
.B(n_1917),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2108),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2061),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2112),
.B(n_1962),
.Y(n_2529)
);

AND2x2_ASAP7_75t_SL g2530 ( 
.A(n_2126),
.B(n_1962),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2021),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2021),
.Y(n_2532)
);

BUFx4f_ASAP7_75t_L g2533 ( 
.A(n_2246),
.Y(n_2533)
);

AO21x2_ASAP7_75t_L g2534 ( 
.A1(n_2191),
.A2(n_1847),
.B(n_1956),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_2115),
.B(n_1971),
.Y(n_2535)
);

OR2x6_ASAP7_75t_L g2536 ( 
.A(n_2290),
.B(n_1730),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2046),
.B(n_1927),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2021),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2062),
.Y(n_2539)
);

OR2x2_ASAP7_75t_L g2540 ( 
.A(n_2264),
.B(n_1928),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2064),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2126),
.A2(n_1902),
.B1(n_1905),
.B2(n_1293),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2144),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2045),
.B(n_1986),
.Y(n_2544)
);

AO21x2_ASAP7_75t_L g2545 ( 
.A1(n_2200),
.A2(n_1966),
.B(n_1941),
.Y(n_2545)
);

INVx4_ASAP7_75t_L g2546 ( 
.A(n_2115),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2144),
.Y(n_2547)
);

OR2x2_ASAP7_75t_L g2548 ( 
.A(n_2290),
.B(n_1960),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2065),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2115),
.B(n_2136),
.Y(n_2550)
);

BUFx4f_ASAP7_75t_L g2551 ( 
.A(n_2246),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2259),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2259),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2068),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2259),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2085),
.Y(n_2556)
);

INVx4_ASAP7_75t_L g2557 ( 
.A(n_2115),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2073),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2020),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2080),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2089),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2189),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2091),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2179),
.B(n_1934),
.Y(n_2564)
);

AND2x6_ASAP7_75t_L g2565 ( 
.A(n_2116),
.B(n_1971),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2092),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2098),
.Y(n_2567)
);

AOI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_2024),
.A2(n_1965),
.B1(n_1979),
.B2(n_1940),
.Y(n_2568)
);

INVxp67_ASAP7_75t_SL g2569 ( 
.A(n_2285),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2099),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2263),
.B(n_1823),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_2285),
.Y(n_2572)
);

BUFx2_ASAP7_75t_L g2573 ( 
.A(n_2118),
.Y(n_2573)
);

BUFx10_ASAP7_75t_L g2574 ( 
.A(n_2037),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2194),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2101),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2103),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2194),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2115),
.B(n_1971),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2198),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2126),
.A2(n_1022),
.B1(n_735),
.B2(n_744),
.Y(n_2581)
);

AO22x2_ASAP7_75t_L g2582 ( 
.A1(n_2187),
.A2(n_1975),
.B1(n_1964),
.B2(n_1942),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2136),
.B(n_1971),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2136),
.B(n_1974),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2105),
.Y(n_2585)
);

AOI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2024),
.A2(n_1944),
.B1(n_1947),
.B2(n_1939),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2273),
.B(n_1841),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2031),
.B(n_1934),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2198),
.Y(n_2589)
);

INVx8_ASAP7_75t_L g2590 ( 
.A(n_2246),
.Y(n_2590)
);

INVxp33_ASAP7_75t_L g2591 ( 
.A(n_2133),
.Y(n_2591)
);

AND2x6_ASAP7_75t_L g2592 ( 
.A(n_2209),
.B(n_1974),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2107),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2136),
.B(n_1974),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2283),
.B(n_1951),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2199),
.B(n_1970),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2119),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2057),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2202),
.B(n_2204),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2234),
.B(n_1974),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2125),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2139),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2179),
.B(n_1937),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2125),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2120),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2206),
.B(n_1981),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2125),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2121),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2140),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2140),
.Y(n_2610)
);

BUFx6f_ASAP7_75t_SL g2611 ( 
.A(n_2234),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2123),
.Y(n_2612)
);

AND2x6_ASAP7_75t_L g2613 ( 
.A(n_2029),
.B(n_1976),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2124),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2020),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2140),
.Y(n_2616)
);

BUFx3_ASAP7_75t_L g2617 ( 
.A(n_2234),
.Y(n_2617)
);

BUFx10_ASAP7_75t_L g2618 ( 
.A(n_2139),
.Y(n_2618)
);

AND2x2_ASAP7_75t_SL g2619 ( 
.A(n_2311),
.B(n_1976),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2148),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2285),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2148),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2128),
.Y(n_2623)
);

INVx2_ASAP7_75t_SL g2624 ( 
.A(n_2139),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2148),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2303),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2213),
.B(n_1993),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2208),
.Y(n_2628)
);

BUFx2_ASAP7_75t_L g2629 ( 
.A(n_2142),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2214),
.B(n_1779),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2215),
.B(n_1779),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2129),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2311),
.A2(n_1022),
.B1(n_743),
.B2(n_747),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2132),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2138),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2151),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2153),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2156),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2146),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2232),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2217),
.B(n_1786),
.Y(n_2641)
);

INVx2_ASAP7_75t_SL g2642 ( 
.A(n_2146),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2157),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2232),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2031),
.B(n_1937),
.Y(n_2645)
);

AOI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2311),
.A2(n_743),
.B1(n_747),
.B2(n_744),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_2196),
.B(n_1948),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2239),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2236),
.A2(n_749),
.B1(n_914),
.B2(n_828),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2239),
.Y(n_2650)
);

INVxp67_ASAP7_75t_L g2651 ( 
.A(n_2223),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2146),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2218),
.B(n_1786),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2161),
.Y(n_2654)
);

AOI21x1_ASAP7_75t_L g2655 ( 
.A1(n_2012),
.A2(n_1915),
.B(n_1376),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2201),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2223),
.B(n_1948),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2208),
.Y(n_2658)
);

AO22x2_ASAP7_75t_L g2659 ( 
.A1(n_2094),
.A2(n_1932),
.B1(n_1925),
.B2(n_1949),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2161),
.Y(n_2660)
);

BUFx10_ASAP7_75t_L g2661 ( 
.A(n_2161),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2208),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2180),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2180),
.Y(n_2664)
);

INVx5_ASAP7_75t_L g2665 ( 
.A(n_2308),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2094),
.B(n_1976),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2180),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2164),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2230),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2201),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2203),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2203),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2452),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2337),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2491),
.B(n_1976),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_2323),
.B(n_1688),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2323),
.B(n_1694),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2337),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2392),
.B(n_2395),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2392),
.B(n_2395),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2464),
.B(n_2102),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2342),
.B(n_1694),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2340),
.B(n_2219),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2375),
.Y(n_2684)
);

INVx3_ASAP7_75t_L g2685 ( 
.A(n_2330),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2318),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_2489),
.Y(n_2687)
);

AND2x2_ASAP7_75t_SL g2688 ( 
.A(n_2581),
.B(n_1991),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2375),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2340),
.B(n_2224),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2350),
.B(n_2225),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2350),
.B(n_2227),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2377),
.Y(n_2693)
);

NAND3xp33_ASAP7_75t_SL g2694 ( 
.A(n_2338),
.B(n_1700),
.C(n_1650),
.Y(n_2694)
);

CKINVDCx20_ASAP7_75t_R g2695 ( 
.A(n_2447),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2367),
.B(n_2240),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_L g2697 ( 
.A(n_2342),
.B(n_1700),
.Y(n_2697)
);

BUFx3_ASAP7_75t_L g2698 ( 
.A(n_2347),
.Y(n_2698)
);

NOR2xp67_ASAP7_75t_SL g2699 ( 
.A(n_2665),
.B(n_1991),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2364),
.B(n_1802),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2322),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2324),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2367),
.B(n_2445),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_2389),
.A2(n_2236),
.B1(n_2235),
.B2(n_2231),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2341),
.B(n_2147),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2377),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2364),
.B(n_2102),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2509),
.B(n_1991),
.Y(n_2708)
);

INVxp33_ASAP7_75t_L g2709 ( 
.A(n_2507),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2327),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2383),
.B(n_2110),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2379),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2483),
.B(n_2240),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_2509),
.B(n_1991),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2383),
.B(n_2110),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2473),
.B(n_1992),
.Y(n_2716)
);

BUFx6f_ASAP7_75t_L g2717 ( 
.A(n_2626),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2401),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2379),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2670),
.Y(n_2720)
);

BUFx2_ASAP7_75t_R g2721 ( 
.A(n_2489),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2488),
.B(n_2134),
.Y(n_2722)
);

NOR2xp67_ASAP7_75t_L g2723 ( 
.A(n_2423),
.B(n_1989),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2473),
.B(n_2134),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2361),
.B(n_2162),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2657),
.B(n_1992),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2361),
.B(n_2162),
.Y(n_2727)
);

INVx3_ASAP7_75t_L g2728 ( 
.A(n_2330),
.Y(n_2728)
);

INVxp67_ASAP7_75t_SL g2729 ( 
.A(n_2569),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2588),
.B(n_2167),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2657),
.B(n_1992),
.Y(n_2731)
);

CKINVDCx14_ASAP7_75t_R g2732 ( 
.A(n_2457),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2349),
.B(n_2365),
.Y(n_2733)
);

INVx2_ASAP7_75t_SL g2734 ( 
.A(n_2419),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2670),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2588),
.B(n_2167),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2645),
.B(n_2241),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2645),
.B(n_1992),
.Y(n_2738)
);

INVx5_ASAP7_75t_L g2739 ( 
.A(n_2472),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2334),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_L g2741 ( 
.A(n_2349),
.B(n_1868),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_SL g2742 ( 
.A(n_2564),
.B(n_1925),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_SL g2743 ( 
.A(n_2370),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2526),
.B(n_2155),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2505),
.Y(n_2745)
);

BUFx6f_ASAP7_75t_L g2746 ( 
.A(n_2626),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2438),
.B(n_2279),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2407),
.B(n_1932),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2520),
.B(n_2279),
.Y(n_2749)
);

NOR2xp67_ASAP7_75t_L g2750 ( 
.A(n_2409),
.B(n_1989),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2461),
.B(n_1649),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2335),
.Y(n_2752)
);

NAND3xp33_ASAP7_75t_L g2753 ( 
.A(n_2510),
.B(n_2113),
.C(n_2106),
.Y(n_2753)
);

NOR2xp67_ASAP7_75t_L g2754 ( 
.A(n_2409),
.B(n_1989),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2671),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2540),
.B(n_2190),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2470),
.B(n_1415),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_SL g2758 ( 
.A(n_2603),
.B(n_2269),
.Y(n_2758)
);

HB1xp67_ASAP7_75t_L g2759 ( 
.A(n_2437),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2543),
.B(n_2280),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2391),
.B(n_1415),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2345),
.Y(n_2762)
);

HB1xp67_ASAP7_75t_L g2763 ( 
.A(n_2451),
.Y(n_2763)
);

INVx2_ASAP7_75t_SL g2764 ( 
.A(n_2321),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2600),
.B(n_2291),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2600),
.B(n_2292),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2671),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2391),
.B(n_1424),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2537),
.B(n_2595),
.Y(n_2769)
);

OAI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2524),
.A2(n_2067),
.B(n_2042),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2537),
.B(n_2168),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2348),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2354),
.Y(n_2773)
);

NOR3xp33_ASAP7_75t_L g2774 ( 
.A(n_2666),
.B(n_1853),
.C(n_2313),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2355),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2672),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2510),
.B(n_2141),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2544),
.B(n_2170),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2356),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2406),
.B(n_1424),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2544),
.B(n_2325),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2410),
.B(n_2252),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2672),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2455),
.A2(n_2249),
.B(n_2253),
.C(n_2242),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2325),
.B(n_2172),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2474),
.B(n_2173),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_2505),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_2326),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2406),
.B(n_1429),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2415),
.B(n_2141),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2446),
.B(n_2181),
.Y(n_2791)
);

OR2x6_ASAP7_75t_L g2792 ( 
.A(n_2362),
.B(n_1730),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2562),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_2371),
.B(n_1429),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2562),
.Y(n_2795)
);

OAI221xp5_ASAP7_75t_L g2796 ( 
.A1(n_2411),
.A2(n_2159),
.B1(n_2255),
.B2(n_2254),
.C(n_2238),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2363),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2369),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2465),
.B(n_2184),
.Y(n_2799)
);

OR2x6_ASAP7_75t_L g2800 ( 
.A(n_2362),
.B(n_1995),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2373),
.Y(n_2801)
);

A2O1A1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2666),
.A2(n_2159),
.B(n_2186),
.C(n_2185),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_SL g2803 ( 
.A(n_2514),
.B(n_2471),
.Y(n_2803)
);

INVx2_ASAP7_75t_SL g2804 ( 
.A(n_2434),
.Y(n_2804)
);

NOR3xp33_ASAP7_75t_L g2805 ( 
.A(n_2376),
.B(n_1901),
.C(n_1620),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2548),
.B(n_2221),
.Y(n_2806)
);

INVx2_ASAP7_75t_SL g2807 ( 
.A(n_2397),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2543),
.B(n_2280),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2336),
.B(n_1430),
.Y(n_2809)
);

BUFx5_ASAP7_75t_L g2810 ( 
.A(n_2472),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2374),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2344),
.A2(n_2267),
.B1(n_2268),
.B2(n_2265),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2415),
.B(n_1989),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2336),
.B(n_2460),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2460),
.B(n_1430),
.Y(n_2815)
);

BUFx5_ASAP7_75t_L g2816 ( 
.A(n_2472),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2410),
.B(n_1443),
.Y(n_2817)
);

NAND3xp33_ASAP7_75t_L g2818 ( 
.A(n_2581),
.B(n_1852),
.C(n_1808),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2547),
.B(n_2294),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2651),
.B(n_1443),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2343),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2515),
.B(n_2243),
.Y(n_2822)
);

NAND2xp33_ASAP7_75t_L g2823 ( 
.A(n_2565),
.B(n_2136),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2651),
.B(n_1444),
.Y(n_2824)
);

INVxp67_ASAP7_75t_L g2825 ( 
.A(n_2573),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2380),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2568),
.B(n_2085),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2547),
.B(n_2294),
.Y(n_2828)
);

NOR2xp33_ASAP7_75t_L g2829 ( 
.A(n_2453),
.B(n_1444),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2453),
.B(n_1453),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2320),
.B(n_2297),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2420),
.B(n_1453),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2420),
.B(n_1456),
.Y(n_2833)
);

OR2x2_ASAP7_75t_L g2834 ( 
.A(n_2629),
.B(n_2251),
.Y(n_2834)
);

NOR3xp33_ASAP7_75t_L g2835 ( 
.A(n_2647),
.B(n_2256),
.C(n_2252),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2647),
.B(n_1456),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2381),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2384),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2399),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_SL g2840 ( 
.A(n_2586),
.B(n_2617),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2466),
.B(n_2271),
.Y(n_2841)
);

INVx2_ASAP7_75t_SL g2842 ( 
.A(n_2536),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2476),
.B(n_2297),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2344),
.B(n_2256),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2447),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2591),
.B(n_1474),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2479),
.B(n_2299),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2408),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2344),
.B(n_2591),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2484),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2486),
.Y(n_2851)
);

BUFx2_ASAP7_75t_R g2852 ( 
.A(n_2615),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2617),
.B(n_1147),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2439),
.B(n_2085),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2496),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2500),
.B(n_2504),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2596),
.B(n_1474),
.Y(n_2857)
);

NAND2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2333),
.B(n_2308),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2536),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2516),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2353),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2518),
.B(n_2528),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2539),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2541),
.B(n_2549),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2554),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2320),
.B(n_2299),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2328),
.B(n_2304),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2558),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2360),
.Y(n_2869)
);

BUFx4_ASAP7_75t_L g2870 ( 
.A(n_2403),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2626),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2328),
.B(n_2304),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2368),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2667),
.B(n_2088),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2448),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2560),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2497),
.B(n_2314),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2497),
.B(n_2314),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2501),
.B(n_2281),
.Y(n_2879)
);

NAND3xp33_ASAP7_75t_L g2880 ( 
.A(n_2649),
.B(n_1852),
.C(n_1808),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2454),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_R g2882 ( 
.A(n_2362),
.B(n_1484),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2456),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2458),
.Y(n_2884)
);

INVx2_ASAP7_75t_SL g2885 ( 
.A(n_2536),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2561),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2667),
.B(n_1151),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2606),
.B(n_1484),
.Y(n_2888)
);

AOI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2398),
.A2(n_2284),
.B1(n_2312),
.B2(n_2282),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2501),
.B(n_2512),
.Y(n_2890)
);

BUFx6f_ASAP7_75t_SL g2891 ( 
.A(n_2370),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2530),
.B(n_2088),
.Y(n_2892)
);

AOI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2398),
.A2(n_2316),
.B1(n_2317),
.B2(n_2315),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2468),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2563),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2627),
.B(n_1496),
.Y(n_2896)
);

BUFx6f_ASAP7_75t_L g2897 ( 
.A(n_2626),
.Y(n_2897)
);

BUFx6f_ASAP7_75t_L g2898 ( 
.A(n_2332),
.Y(n_2898)
);

NAND2xp33_ASAP7_75t_L g2899 ( 
.A(n_2565),
.B(n_2169),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2512),
.B(n_2070),
.Y(n_2900)
);

AND2x4_ASAP7_75t_SL g2901 ( 
.A(n_2618),
.B(n_1811),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_SL g2902 ( 
.A(n_2530),
.B(n_2088),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_2427),
.B(n_2088),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2566),
.B(n_2152),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2567),
.B(n_2152),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2570),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2469),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2493),
.B(n_2152),
.Y(n_2908)
);

NOR2x1p5_ASAP7_75t_L g2909 ( 
.A(n_2393),
.B(n_1882),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2669),
.B(n_1496),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2576),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_SL g2912 ( 
.A(n_2665),
.B(n_1899),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2669),
.B(n_1503),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_2577),
.B(n_1503),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2480),
.Y(n_2915)
);

AND2x4_ASAP7_75t_L g2916 ( 
.A(n_2351),
.B(n_2216),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2585),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2593),
.B(n_2152),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2597),
.B(n_2160),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2498),
.B(n_2160),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2482),
.Y(n_2921)
);

INVx3_ASAP7_75t_L g2922 ( 
.A(n_2366),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2319),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_2331),
.B(n_1521),
.Y(n_2924)
);

NOR3xp33_ASAP7_75t_L g2925 ( 
.A(n_2394),
.B(n_1528),
.C(n_1521),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2605),
.B(n_2160),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2608),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2503),
.B(n_2160),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2612),
.Y(n_2929)
);

OR2x6_ASAP7_75t_L g2930 ( 
.A(n_2393),
.B(n_1995),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_SL g2931 ( 
.A(n_2428),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2614),
.B(n_2177),
.Y(n_2932)
);

INVx3_ASAP7_75t_L g2933 ( 
.A(n_2366),
.Y(n_2933)
);

NOR2xp67_ASAP7_75t_L g2934 ( 
.A(n_2623),
.B(n_2216),
.Y(n_2934)
);

INVx2_ASAP7_75t_SL g2935 ( 
.A(n_2319),
.Y(n_2935)
);

NAND2xp33_ASAP7_75t_L g2936 ( 
.A(n_2565),
.B(n_2169),
.Y(n_2936)
);

INVx3_ASAP7_75t_L g2937 ( 
.A(n_2425),
.Y(n_2937)
);

HB1xp67_ASAP7_75t_L g2938 ( 
.A(n_2611),
.Y(n_2938)
);

CKINVDCx5p33_ASAP7_75t_R g2939 ( 
.A(n_2508),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_SL g2940 ( 
.A(n_2519),
.B(n_2177),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2385),
.B(n_2169),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2598),
.B(n_2177),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2425),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2331),
.B(n_1528),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2499),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2602),
.B(n_2177),
.Y(n_2946)
);

NOR2xp67_ASAP7_75t_L g2947 ( 
.A(n_2632),
.B(n_2220),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2634),
.Y(n_2948)
);

AO21x2_ASAP7_75t_L g2949 ( 
.A1(n_2329),
.A2(n_2301),
.B(n_2261),
.Y(n_2949)
);

INVx3_ASAP7_75t_L g2950 ( 
.A(n_2432),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2385),
.B(n_2169),
.Y(n_2951)
);

AO21x2_ASAP7_75t_L g2952 ( 
.A1(n_2329),
.A2(n_2250),
.B(n_2226),
.Y(n_2952)
);

BUFx2_ASAP7_75t_R g2953 ( 
.A(n_2428),
.Y(n_2953)
);

INVxp67_ASAP7_75t_SL g2954 ( 
.A(n_2569),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2386),
.B(n_2169),
.Y(n_2955)
);

BUFx5_ASAP7_75t_L g2956 ( 
.A(n_2472),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2386),
.B(n_2171),
.Y(n_2957)
);

AND2x4_ASAP7_75t_L g2958 ( 
.A(n_2351),
.B(n_2220),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2358),
.B(n_1536),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2624),
.B(n_1151),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2387),
.B(n_2171),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2635),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2636),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2358),
.B(n_1536),
.Y(n_2964)
);

NAND2xp33_ASAP7_75t_SL g2965 ( 
.A(n_2611),
.B(n_1967),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2707),
.B(n_2659),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2733),
.B(n_2711),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2700),
.B(n_1546),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2715),
.B(n_2637),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2674),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2688),
.A2(n_2582),
.B1(n_2654),
.B2(n_2652),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2850),
.Y(n_2972)
);

NAND2xp33_ASAP7_75t_L g2973 ( 
.A(n_2781),
.B(n_2565),
.Y(n_2973)
);

O2A1O1Ixp33_ASAP7_75t_L g2974 ( 
.A1(n_2790),
.A2(n_2724),
.B(n_2727),
.C(n_2725),
.Y(n_2974)
);

NAND2xp33_ASAP7_75t_L g2975 ( 
.A(n_2738),
.B(n_2565),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2703),
.B(n_2387),
.Y(n_2976)
);

INVx2_ASAP7_75t_SL g2977 ( 
.A(n_2698),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2851),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_SL g2979 ( 
.A(n_2803),
.B(n_2618),
.Y(n_2979)
);

INVx5_ASAP7_75t_L g2980 ( 
.A(n_2739),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2703),
.B(n_2388),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2769),
.B(n_2388),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2696),
.B(n_2390),
.Y(n_2983)
);

BUFx3_ASAP7_75t_L g2984 ( 
.A(n_2804),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2678),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2684),
.Y(n_2986)
);

INVx2_ASAP7_75t_SL g2987 ( 
.A(n_2807),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2713),
.B(n_2638),
.Y(n_2988)
);

AND2x4_ASAP7_75t_L g2989 ( 
.A(n_2842),
.B(n_2859),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2753),
.A2(n_2925),
.B1(n_2844),
.B2(n_2694),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2741),
.B(n_1546),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_2682),
.B(n_1552),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2855),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2860),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2697),
.B(n_1552),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2689),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2722),
.B(n_2643),
.Y(n_2997)
);

CKINVDCx20_ASAP7_75t_R g2998 ( 
.A(n_2695),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_SL g2999 ( 
.A(n_2803),
.B(n_2661),
.Y(n_2999)
);

AND2x4_ASAP7_75t_L g3000 ( 
.A(n_2885),
.B(n_2499),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2863),
.Y(n_3001)
);

INVx4_ASAP7_75t_L g3002 ( 
.A(n_2717),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2717),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2748),
.B(n_2661),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2696),
.B(n_2639),
.Y(n_3005)
);

INVxp67_ASAP7_75t_L g3006 ( 
.A(n_2759),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2857),
.B(n_2642),
.Y(n_3007)
);

O2A1O1Ixp33_ASAP7_75t_L g3008 ( 
.A1(n_2676),
.A2(n_2394),
.B(n_2522),
.C(n_2372),
.Y(n_3008)
);

INVx8_ASAP7_75t_L g3009 ( 
.A(n_2792),
.Y(n_3009)
);

INVx2_ASAP7_75t_SL g3010 ( 
.A(n_2763),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2730),
.B(n_2660),
.Y(n_3011)
);

O2A1O1Ixp33_ASAP7_75t_L g3012 ( 
.A1(n_2677),
.A2(n_2339),
.B(n_2396),
.C(n_2378),
.Y(n_3012)
);

OR2x6_ASAP7_75t_L g3013 ( 
.A(n_2792),
.B(n_2478),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2693),
.Y(n_3014)
);

AOI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2761),
.A2(n_2768),
.B1(n_2789),
.B2(n_2780),
.Y(n_3015)
);

AOI22xp5_ASAP7_75t_L g3016 ( 
.A1(n_2829),
.A2(n_1563),
.B1(n_1571),
.B2(n_1566),
.Y(n_3016)
);

AND2x4_ASAP7_75t_SL g3017 ( 
.A(n_2792),
.B(n_2508),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2777),
.B(n_1563),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_2705),
.B(n_2559),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2706),
.Y(n_3020)
);

INVxp67_ASAP7_75t_L g3021 ( 
.A(n_2914),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2712),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2736),
.B(n_2663),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2681),
.B(n_2664),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2849),
.A2(n_2582),
.B1(n_2433),
.B2(n_2659),
.Y(n_3025)
);

INVx2_ASAP7_75t_SL g3026 ( 
.A(n_2718),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2782),
.B(n_2582),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2888),
.B(n_2478),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2830),
.A2(n_1566),
.B1(n_1576),
.B2(n_1571),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2785),
.B(n_2646),
.Y(n_3030)
);

INVx2_ASAP7_75t_SL g3031 ( 
.A(n_2734),
.Y(n_3031)
);

A2O1A1Ixp33_ASAP7_75t_L g3032 ( 
.A1(n_2737),
.A2(n_2481),
.B(n_2422),
.C(n_2633),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2744),
.B(n_2646),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2806),
.B(n_2668),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2832),
.B(n_1576),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2756),
.B(n_2619),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2786),
.B(n_2619),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2833),
.B(n_1582),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_SL g3039 ( 
.A1(n_2836),
.A2(n_1582),
.B1(n_1967),
.B2(n_1656),
.Y(n_3039)
);

NAND3xp33_ASAP7_75t_SL g3040 ( 
.A(n_2774),
.B(n_1663),
.C(n_1622),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_2896),
.B(n_2382),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2719),
.Y(n_3042)
);

BUFx3_ASAP7_75t_L g3043 ( 
.A(n_2673),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2679),
.B(n_2390),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2835),
.B(n_2856),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2862),
.B(n_2633),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2864),
.B(n_2433),
.Y(n_3047)
);

OAI22xp5_ASAP7_75t_L g3048 ( 
.A1(n_2679),
.A2(n_2422),
.B1(n_2477),
.B2(n_2462),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2817),
.B(n_2820),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2924),
.A2(n_2433),
.B1(n_2659),
.B2(n_2649),
.Y(n_3050)
);

AOI22xp5_ASAP7_75t_L g3051 ( 
.A1(n_2757),
.A2(n_1995),
.B1(n_1663),
.B2(n_1656),
.Y(n_3051)
);

AOI22xp33_ASAP7_75t_L g3052 ( 
.A1(n_2944),
.A2(n_2417),
.B1(n_2429),
.B2(n_2416),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2865),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2824),
.B(n_1622),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2793),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2751),
.B(n_2382),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2771),
.B(n_2525),
.Y(n_3057)
);

INVx3_ASAP7_75t_L g3058 ( 
.A(n_2685),
.Y(n_3058)
);

INVxp67_ASAP7_75t_SL g3059 ( 
.A(n_2729),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2795),
.Y(n_3060)
);

A2O1A1Ixp33_ASAP7_75t_L g3061 ( 
.A1(n_2784),
.A2(n_2587),
.B(n_2443),
.C(n_2459),
.Y(n_3061)
);

O2A1O1Ixp33_ASAP7_75t_L g3062 ( 
.A1(n_2796),
.A2(n_2402),
.B(n_2424),
.C(n_2414),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2720),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2868),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_SL g3065 ( 
.A(n_2764),
.B(n_2788),
.Y(n_3065)
);

INVx3_ASAP7_75t_L g3066 ( 
.A(n_2685),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2959),
.B(n_2527),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2735),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2876),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2778),
.B(n_2525),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2755),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2954),
.B(n_2527),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2767),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2886),
.B(n_2450),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2794),
.B(n_1625),
.Y(n_3075)
);

AOI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_2846),
.A2(n_1751),
.B1(n_2414),
.B2(n_2402),
.Y(n_3076)
);

OAI22xp5_ASAP7_75t_SL g3077 ( 
.A1(n_2818),
.A2(n_1627),
.B1(n_1625),
.B2(n_749),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2964),
.B(n_2640),
.Y(n_3078)
);

INVx2_ASAP7_75t_SL g3079 ( 
.A(n_2901),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2709),
.B(n_2825),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2895),
.B(n_2644),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2906),
.B(n_2650),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2910),
.B(n_1627),
.Y(n_3083)
);

A2O1A1Ixp33_ASAP7_75t_L g3084 ( 
.A1(n_2704),
.A2(n_2599),
.B(n_2357),
.C(n_2444),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2911),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2917),
.B(n_2648),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2927),
.B(n_2440),
.Y(n_3087)
);

AOI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2913),
.A2(n_2444),
.B1(n_2467),
.B2(n_2424),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2776),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2783),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2929),
.B(n_2440),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_2758),
.A2(n_2765),
.B1(n_2766),
.B2(n_2840),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2948),
.B(n_2441),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_SL g3094 ( 
.A(n_2822),
.B(n_2665),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2962),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_SL g3096 ( 
.A(n_2912),
.B(n_2665),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2963),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2749),
.B(n_2441),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2809),
.B(n_2467),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2686),
.Y(n_3100)
);

OAI22xp5_ASAP7_75t_L g3101 ( 
.A1(n_2680),
.A2(n_2477),
.B1(n_2517),
.B2(n_2462),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_2813),
.A2(n_2475),
.B1(n_2529),
.B2(n_2511),
.Y(n_3102)
);

AOI22xp33_ASAP7_75t_L g3103 ( 
.A1(n_2742),
.A2(n_2475),
.B1(n_2529),
.B2(n_2511),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_2815),
.B(n_2834),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2887),
.B(n_2574),
.Y(n_3105)
);

NAND3xp33_ASAP7_75t_SL g3106 ( 
.A(n_2805),
.B(n_2571),
.C(n_914),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2701),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2912),
.B(n_2332),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2965),
.A2(n_2579),
.B1(n_2583),
.B2(n_2535),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2821),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2853),
.B(n_2332),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_2953),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2749),
.B(n_2442),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2747),
.B(n_2442),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2708),
.B(n_2535),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2702),
.Y(n_3116)
);

INVxp67_ASAP7_75t_L g3117 ( 
.A(n_2938),
.Y(n_3117)
);

INVx1_ASAP7_75t_SL g3118 ( 
.A(n_2882),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2680),
.B(n_2412),
.Y(n_3119)
);

AND2x6_ASAP7_75t_SL g3120 ( 
.A(n_2814),
.B(n_1987),
.Y(n_3120)
);

NAND2x1p5_ASAP7_75t_L g3121 ( 
.A(n_2699),
.B(n_2432),
.Y(n_3121)
);

AND2x4_ASAP7_75t_L g3122 ( 
.A(n_2923),
.B(n_2583),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2747),
.B(n_2412),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2683),
.B(n_2413),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2683),
.B(n_2413),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_2714),
.A2(n_2675),
.B1(n_2812),
.B2(n_2731),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2861),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2728),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2799),
.B(n_2841),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2726),
.B(n_2880),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2869),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2710),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2916),
.B(n_2513),
.Y(n_3133)
);

AND3x1_ASAP7_75t_L g3134 ( 
.A(n_2960),
.B(n_2802),
.C(n_2935),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_SL g3135 ( 
.A(n_2750),
.B(n_2332),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2916),
.A2(n_2584),
.B1(n_2594),
.B2(n_2579),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2958),
.B(n_2574),
.Y(n_3137)
);

OAI22xp5_ASAP7_75t_L g3138 ( 
.A1(n_2690),
.A2(n_2517),
.B1(n_2542),
.B2(n_2421),
.Y(n_3138)
);

AND2x6_ASAP7_75t_SL g3139 ( 
.A(n_2930),
.B(n_2800),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_SL g3140 ( 
.A(n_2754),
.B(n_2495),
.Y(n_3140)
);

A2O1A1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_2791),
.A2(n_2594),
.B(n_2584),
.C(n_2533),
.Y(n_3141)
);

AOI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_2732),
.A2(n_1731),
.B1(n_2592),
.B2(n_2492),
.Y(n_3142)
);

BUFx6f_ASAP7_75t_L g3143 ( 
.A(n_2717),
.Y(n_3143)
);

AND2x4_ASAP7_75t_L g3144 ( 
.A(n_2945),
.B(n_2485),
.Y(n_3144)
);

AND2x6_ASAP7_75t_SL g3145 ( 
.A(n_2930),
.B(n_1987),
.Y(n_3145)
);

INVxp67_ASAP7_75t_L g3146 ( 
.A(n_2852),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2716),
.B(n_1731),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_2728),
.Y(n_3148)
);

INVx5_ASAP7_75t_L g3149 ( 
.A(n_2739),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2958),
.B(n_2495),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2800),
.B(n_2487),
.Y(n_3151)
);

AND2x6_ASAP7_75t_SL g3152 ( 
.A(n_2930),
.B(n_1370),
.Y(n_3152)
);

O2A1O1Ixp33_ASAP7_75t_L g3153 ( 
.A1(n_2854),
.A2(n_2631),
.B(n_2641),
.C(n_2630),
.Y(n_3153)
);

AOI22xp33_ASAP7_75t_L g3154 ( 
.A1(n_2827),
.A2(n_2875),
.B1(n_2883),
.B2(n_2881),
.Y(n_3154)
);

BUFx8_ASAP7_75t_L g3155 ( 
.A(n_2743),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2740),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_2723),
.A2(n_2592),
.B1(n_2472),
.B2(n_2492),
.Y(n_3157)
);

O2A1O1Ixp5_ASAP7_75t_L g3158 ( 
.A1(n_2770),
.A2(n_2655),
.B(n_2533),
.C(n_2551),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_2884),
.A2(n_2492),
.B1(n_2575),
.B2(n_2494),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2873),
.Y(n_3160)
);

O2A1O1Ixp33_ASAP7_75t_L g3161 ( 
.A1(n_2892),
.A2(n_2653),
.B(n_2207),
.C(n_2257),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2752),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2894),
.A2(n_2492),
.B1(n_2580),
.B2(n_2578),
.Y(n_3163)
);

OAI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_2800),
.A2(n_2939),
.B1(n_2845),
.B2(n_2905),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2690),
.B(n_2513),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2691),
.B(n_2521),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2762),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2907),
.B(n_2589),
.Y(n_3168)
);

NOR2x2_ASAP7_75t_L g3169 ( 
.A(n_2915),
.B(n_2656),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_2922),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2772),
.Y(n_3171)
);

NAND2x1p5_ASAP7_75t_L g3172 ( 
.A(n_2739),
.B(n_2922),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2691),
.B(n_2521),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2773),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2692),
.B(n_2532),
.Y(n_3175)
);

INVx2_ASAP7_75t_SL g3176 ( 
.A(n_2870),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2692),
.B(n_2532),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2775),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_2933),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2843),
.B(n_2538),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2847),
.B(n_2538),
.Y(n_3181)
);

AOI22xp33_ASAP7_75t_L g3182 ( 
.A1(n_2921),
.A2(n_2492),
.B1(n_2592),
.B2(n_2545),
.Y(n_3182)
);

NAND2x1p5_ASAP7_75t_L g3183 ( 
.A(n_2739),
.B(n_2435),
.Y(n_3183)
);

AOI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_2909),
.A2(n_2592),
.B1(n_2613),
.B2(n_2306),
.Y(n_3184)
);

AND2x2_ASAP7_75t_SL g3185 ( 
.A(n_2823),
.B(n_2502),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2890),
.B(n_2418),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2779),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2797),
.A2(n_2542),
.B1(n_2421),
.B2(n_2426),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_2687),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2967),
.B(n_2798),
.Y(n_3190)
);

HB1xp67_ASAP7_75t_L g3191 ( 
.A(n_3010),
.Y(n_3191)
);

AOI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_3032),
.A2(n_2936),
.B(n_2899),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_3141),
.A2(n_2770),
.B(n_2551),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_3138),
.A2(n_2502),
.B(n_2902),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_3162),
.Y(n_3195)
);

INVx3_ASAP7_75t_L g3196 ( 
.A(n_2980),
.Y(n_3196)
);

O2A1O1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_3028),
.A2(n_2874),
.B(n_2942),
.C(n_2940),
.Y(n_3197)
);

OAI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_3015),
.A2(n_2947),
.B(n_2934),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_L g3199 ( 
.A(n_2992),
.B(n_2745),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3138),
.A2(n_2900),
.B(n_2858),
.Y(n_3200)
);

BUFx4f_ASAP7_75t_L g3201 ( 
.A(n_3009),
.Y(n_3201)
);

BUFx6f_ASAP7_75t_L g3202 ( 
.A(n_3009),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3129),
.B(n_3049),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2997),
.B(n_2801),
.Y(n_3204)
);

OAI321xp33_ASAP7_75t_L g3205 ( 
.A1(n_3050),
.A2(n_2926),
.A3(n_2918),
.B1(n_2932),
.B2(n_2919),
.C(n_2904),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_3171),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_3110),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3078),
.B(n_2811),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_2973),
.A2(n_2900),
.B(n_2531),
.Y(n_3209)
);

A2O1A1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2974),
.A2(n_2893),
.B(n_2889),
.C(n_2837),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2975),
.A2(n_2531),
.B(n_2550),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3127),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_3045),
.B(n_2826),
.Y(n_3213)
);

AOI21x1_ASAP7_75t_L g3214 ( 
.A1(n_3004),
.A2(n_2553),
.B(n_2552),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2976),
.A2(n_2550),
.B(n_2534),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_SL g3216 ( 
.A(n_3104),
.B(n_2838),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_2995),
.B(n_2787),
.Y(n_3217)
);

AOI21xp5_ASAP7_75t_L g3218 ( 
.A1(n_2976),
.A2(n_2534),
.B(n_2352),
.Y(n_3218)
);

O2A1O1Ixp5_ASAP7_75t_L g3219 ( 
.A1(n_3108),
.A2(n_2908),
.B(n_2920),
.C(n_2903),
.Y(n_3219)
);

NOR3xp33_ASAP7_75t_L g3220 ( 
.A(n_3106),
.B(n_2946),
.C(n_2928),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2981),
.A2(n_2590),
.B(n_2352),
.Y(n_3221)
);

BUFx12f_ASAP7_75t_L g3222 ( 
.A(n_3155),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2988),
.B(n_2839),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_2968),
.B(n_2848),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_3035),
.B(n_2743),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2969),
.B(n_2890),
.Y(n_3226)
);

HB1xp67_ASAP7_75t_L g3227 ( 
.A(n_3006),
.Y(n_3227)
);

NOR2xp33_ASAP7_75t_L g3228 ( 
.A(n_3038),
.B(n_2891),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3099),
.B(n_2879),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2991),
.B(n_2891),
.Y(n_3230)
);

AND2x2_ASAP7_75t_L g3231 ( 
.A(n_3067),
.B(n_1151),
.Y(n_3231)
);

BUFx3_ASAP7_75t_L g3232 ( 
.A(n_2984),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_2981),
.A2(n_2590),
.B(n_2352),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_3185),
.A2(n_2590),
.B(n_2941),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_3008),
.A2(n_2951),
.B(n_2941),
.Y(n_3235)
);

O2A1O1Ixp5_ASAP7_75t_L g3236 ( 
.A1(n_3130),
.A2(n_2879),
.B(n_2955),
.C(n_2951),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2972),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3124),
.A2(n_2957),
.B(n_2955),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3124),
.A2(n_2961),
.B(n_2957),
.Y(n_3239)
);

INVx4_ASAP7_75t_L g3240 ( 
.A(n_2980),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3057),
.B(n_2760),
.Y(n_3241)
);

HB1xp67_ASAP7_75t_L g3242 ( 
.A(n_2987),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_3125),
.A2(n_2961),
.B(n_2247),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3070),
.B(n_2760),
.Y(n_3244)
);

OAI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2990),
.A2(n_2931),
.B1(n_2937),
.B2(n_2933),
.Y(n_3245)
);

BUFx12f_ASAP7_75t_L g3246 ( 
.A(n_3155),
.Y(n_3246)
);

O2A1O1Ixp33_ASAP7_75t_L g3247 ( 
.A1(n_3041),
.A2(n_1380),
.B(n_1382),
.C(n_1378),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3011),
.B(n_2808),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_3018),
.B(n_2810),
.Y(n_3249)
);

NOR2xp33_ASAP7_75t_L g3250 ( 
.A(n_3016),
.B(n_2931),
.Y(n_3250)
);

INVx11_ASAP7_75t_L g3251 ( 
.A(n_3169),
.Y(n_3251)
);

NAND2x1p5_ASAP7_75t_L g3252 ( 
.A(n_2980),
.B(n_2937),
.Y(n_3252)
);

AOI22xp33_ASAP7_75t_L g3253 ( 
.A1(n_3040),
.A2(n_2592),
.B1(n_2545),
.B2(n_2613),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3023),
.B(n_3036),
.Y(n_3254)
);

OAI21xp33_ASAP7_75t_L g3255 ( 
.A1(n_3052),
.A2(n_916),
.B(n_828),
.Y(n_3255)
);

HB1xp67_ASAP7_75t_L g3256 ( 
.A(n_3034),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_SL g3257 ( 
.A(n_3092),
.B(n_2956),
.Y(n_3257)
);

OAI321xp33_ASAP7_75t_L g3258 ( 
.A1(n_3077),
.A2(n_2819),
.A3(n_2828),
.B1(n_2866),
.B2(n_2831),
.C(n_2808),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3037),
.B(n_2819),
.Y(n_3259)
);

AO21x1_ASAP7_75t_L g3260 ( 
.A1(n_3115),
.A2(n_2831),
.B(n_2828),
.Y(n_3260)
);

AOI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3125),
.A2(n_2247),
.B(n_2171),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2978),
.Y(n_3262)
);

AOI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_3075),
.A2(n_3054),
.B1(n_3083),
.B2(n_3056),
.Y(n_3263)
);

OAI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_3012),
.A2(n_3061),
.B(n_3084),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_3076),
.A2(n_2943),
.B1(n_2950),
.B2(n_2306),
.Y(n_3265)
);

A2O1A1Ixp33_ASAP7_75t_L g3266 ( 
.A1(n_3062),
.A2(n_2950),
.B(n_2943),
.C(n_2359),
.Y(n_3266)
);

A2O1A1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_3030),
.A2(n_2359),
.B(n_2400),
.C(n_2346),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3033),
.B(n_2866),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_3043),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_2966),
.B(n_2746),
.Y(n_3270)
);

INVxp67_ASAP7_75t_L g3271 ( 
.A(n_3080),
.Y(n_3271)
);

BUFx6f_ASAP7_75t_L g3272 ( 
.A(n_3009),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_3029),
.B(n_2721),
.Y(n_3273)
);

OAI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_3153),
.A2(n_2872),
.B(n_2867),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3131),
.Y(n_3275)
);

OAI21xp33_ASAP7_75t_L g3276 ( 
.A1(n_3147),
.A2(n_3007),
.B(n_3024),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_3003),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_SL g3278 ( 
.A(n_3164),
.B(n_2810),
.Y(n_3278)
);

OAI22xp33_ASAP7_75t_L g3279 ( 
.A1(n_3051),
.A2(n_3118),
.B1(n_3142),
.B2(n_3019),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_SL g3280 ( 
.A(n_3118),
.B(n_2810),
.Y(n_3280)
);

INVx3_ASAP7_75t_L g3281 ( 
.A(n_2980),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3026),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_3039),
.B(n_2979),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3021),
.B(n_2867),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2993),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3005),
.B(n_2872),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_2983),
.A2(n_2247),
.B(n_2171),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3059),
.B(n_2877),
.Y(n_3288)
);

INVxp67_ASAP7_75t_L g3289 ( 
.A(n_3065),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3074),
.B(n_2877),
.Y(n_3290)
);

INVx2_ASAP7_75t_SL g3291 ( 
.A(n_3017),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_2983),
.A2(n_2247),
.B(n_2171),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3151),
.B(n_2746),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3165),
.A2(n_2278),
.B(n_2247),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_3003),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2999),
.B(n_2746),
.Y(n_3296)
);

A2O1A1Ixp33_ASAP7_75t_L g3297 ( 
.A1(n_3088),
.A2(n_3046),
.B(n_3158),
.C(n_3027),
.Y(n_3297)
);

AOI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_3166),
.A2(n_2278),
.B(n_2183),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3105),
.B(n_2878),
.Y(n_3299)
);

OR2x6_ASAP7_75t_L g3300 ( 
.A(n_3013),
.B(n_3096),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3173),
.A2(n_2278),
.B(n_2183),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2994),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3175),
.A2(n_2278),
.B(n_2183),
.Y(n_3303)
);

NOR2xp67_ASAP7_75t_L g3304 ( 
.A(n_2977),
.B(n_3031),
.Y(n_3304)
);

INVxp67_ASAP7_75t_L g3305 ( 
.A(n_2989),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3001),
.Y(n_3306)
);

INVx11_ASAP7_75t_L g3307 ( 
.A(n_3003),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_3111),
.B(n_3122),
.Y(n_3308)
);

NAND2x1p5_ASAP7_75t_L g3309 ( 
.A(n_3149),
.B(n_2435),
.Y(n_3309)
);

AOI21xp33_ASAP7_75t_L g3310 ( 
.A1(n_2971),
.A2(n_2949),
.B(n_2952),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3168),
.B(n_2878),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3081),
.B(n_2418),
.Y(n_3312)
);

O2A1O1Ixp33_ASAP7_75t_L g3313 ( 
.A1(n_3117),
.A2(n_1387),
.B(n_2207),
.C(n_2165),
.Y(n_3313)
);

INVx3_ASAP7_75t_L g3314 ( 
.A(n_3149),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3082),
.B(n_2426),
.Y(n_3315)
);

AOI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_3177),
.A2(n_2278),
.B(n_2183),
.Y(n_3316)
);

AOI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3079),
.A2(n_2613),
.B1(n_2306),
.B2(n_2182),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_2982),
.A2(n_2182),
.B(n_2431),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_3025),
.A2(n_2306),
.B1(n_2523),
.B2(n_2490),
.Y(n_3319)
);

INVx4_ASAP7_75t_L g3320 ( 
.A(n_3149),
.Y(n_3320)
);

AO21x1_ASAP7_75t_L g3321 ( 
.A1(n_3047),
.A2(n_2523),
.B(n_2490),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3160),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2982),
.B(n_3072),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_L g3324 ( 
.A(n_3112),
.B(n_2871),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3048),
.A2(n_2182),
.B(n_2431),
.Y(n_3325)
);

BUFx3_ASAP7_75t_L g3326 ( 
.A(n_2989),
.Y(n_3326)
);

AOI21xp33_ASAP7_75t_L g3327 ( 
.A1(n_3126),
.A2(n_2949),
.B(n_2952),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3053),
.B(n_2436),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2970),
.Y(n_3329)
);

AOI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_3048),
.A2(n_2182),
.B(n_2436),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3064),
.Y(n_3331)
);

AOI22x1_ASAP7_75t_L g3332 ( 
.A1(n_3069),
.A2(n_2557),
.B1(n_2546),
.B2(n_2346),
.Y(n_3332)
);

AOI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_3149),
.A2(n_2557),
.B(n_2546),
.Y(n_3333)
);

INVx3_ASAP7_75t_L g3334 ( 
.A(n_3172),
.Y(n_3334)
);

O2A1O1Ixp33_ASAP7_75t_L g3335 ( 
.A1(n_3094),
.A2(n_2165),
.B(n_2257),
.C(n_2211),
.Y(n_3335)
);

HB1xp67_ASAP7_75t_L g3336 ( 
.A(n_3000),
.Y(n_3336)
);

NAND2xp33_ASAP7_75t_L g3337 ( 
.A(n_3137),
.B(n_2613),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3085),
.B(n_3095),
.Y(n_3338)
);

AOI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3134),
.A2(n_2613),
.B1(n_916),
.B2(n_921),
.Y(n_3339)
);

OAI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3161),
.A2(n_2211),
.B(n_2205),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3122),
.B(n_2810),
.Y(n_3341)
);

INVx1_ASAP7_75t_SL g3342 ( 
.A(n_3000),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3134),
.B(n_3144),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_SL g3344 ( 
.A(n_3144),
.B(n_2810),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_3172),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3097),
.B(n_2871),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3086),
.B(n_2871),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2985),
.Y(n_3348)
);

O2A1O1Ixp5_ASAP7_75t_L g3349 ( 
.A1(n_3101),
.A2(n_2552),
.B(n_2555),
.C(n_2553),
.Y(n_3349)
);

BUFx2_ASAP7_75t_L g3350 ( 
.A(n_3013),
.Y(n_3350)
);

OAI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3101),
.A2(n_2555),
.B(n_2228),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3100),
.B(n_2897),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_3109),
.B(n_2816),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_3107),
.B(n_2897),
.Y(n_3354)
);

OAI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_3102),
.A2(n_2205),
.B(n_2228),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_3116),
.B(n_2816),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3188),
.A2(n_2621),
.B(n_2572),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3132),
.B(n_2897),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3156),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3167),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_3188),
.A2(n_3123),
.B(n_3113),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3123),
.A2(n_3098),
.B(n_3157),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3114),
.A2(n_2621),
.B(n_2572),
.Y(n_3363)
);

A2O1A1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_3184),
.A2(n_2404),
.B(n_2405),
.C(n_2400),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_2986),
.Y(n_3365)
);

HB1xp67_ASAP7_75t_L g3366 ( 
.A(n_3133),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_3013),
.B(n_2898),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_2996),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3174),
.Y(n_3369)
);

INVx4_ASAP7_75t_L g3370 ( 
.A(n_3143),
.Y(n_3370)
);

OAI21xp33_ASAP7_75t_L g3371 ( 
.A1(n_3154),
.A2(n_921),
.B(n_918),
.Y(n_3371)
);

OAI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3103),
.A2(n_2079),
.B(n_2056),
.Y(n_3372)
);

NOR2x1_ASAP7_75t_L g3373 ( 
.A(n_3058),
.B(n_2404),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3180),
.A2(n_2572),
.B(n_2495),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3181),
.A2(n_2572),
.B(n_2495),
.Y(n_3375)
);

A2O1A1Ixp33_ASAP7_75t_L g3376 ( 
.A1(n_3178),
.A2(n_2430),
.B(n_2449),
.C(n_2405),
.Y(n_3376)
);

AOI21xp5_ASAP7_75t_L g3377 ( 
.A1(n_3044),
.A2(n_3119),
.B(n_3186),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_3187),
.B(n_2816),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3014),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3044),
.A2(n_2621),
.B(n_2662),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_3119),
.A2(n_2621),
.B(n_2662),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_SL g3382 ( 
.A(n_3112),
.B(n_2816),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3186),
.A2(n_2604),
.B(n_2601),
.Y(n_3383)
);

OAI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3136),
.A2(n_2463),
.B1(n_2506),
.B2(n_2430),
.Y(n_3384)
);

BUFx6f_ASAP7_75t_L g3385 ( 
.A(n_3143),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_3182),
.A2(n_2604),
.B(n_2601),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_3121),
.A2(n_2609),
.B(n_2607),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3058),
.B(n_2816),
.Y(n_3388)
);

OAI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3159),
.A2(n_2079),
.B(n_2056),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_3121),
.A2(n_2609),
.B(n_2607),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_3066),
.B(n_2956),
.Y(n_3391)
);

INVx4_ASAP7_75t_L g3392 ( 
.A(n_3143),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3087),
.B(n_2898),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3135),
.A2(n_2616),
.B(n_2610),
.Y(n_3394)
);

CKINVDCx10_ASAP7_75t_R g3395 ( 
.A(n_2998),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3140),
.A2(n_2616),
.B(n_2610),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3020),
.B(n_2898),
.Y(n_3397)
);

AOI21xp5_ASAP7_75t_L g3398 ( 
.A1(n_3183),
.A2(n_2622),
.B(n_2620),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3091),
.B(n_918),
.Y(n_3399)
);

HB1xp67_ASAP7_75t_L g3400 ( 
.A(n_3022),
.Y(n_3400)
);

A2O1A1Ixp33_ASAP7_75t_L g3401 ( 
.A1(n_3163),
.A2(n_2463),
.B(n_2506),
.C(n_2449),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3042),
.Y(n_3402)
);

NOR2xp33_ASAP7_75t_L g3403 ( 
.A(n_3146),
.B(n_1786),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3237),
.Y(n_3404)
);

BUFx4f_ASAP7_75t_L g3405 ( 
.A(n_3222),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3254),
.B(n_3323),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3203),
.B(n_3055),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3229),
.B(n_3060),
.Y(n_3408)
);

BUFx2_ASAP7_75t_L g3409 ( 
.A(n_3256),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_3271),
.B(n_3189),
.Y(n_3410)
);

INVx3_ASAP7_75t_L g3411 ( 
.A(n_3202),
.Y(n_3411)
);

OAI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_3263),
.A2(n_3093),
.B1(n_923),
.B2(n_927),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3259),
.B(n_3063),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3270),
.B(n_3068),
.Y(n_3414)
);

AND2x4_ASAP7_75t_L g3415 ( 
.A(n_3350),
.B(n_3300),
.Y(n_3415)
);

CKINVDCx8_ASAP7_75t_R g3416 ( 
.A(n_3395),
.Y(n_3416)
);

HB1xp67_ASAP7_75t_L g3417 ( 
.A(n_3366),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_L g3418 ( 
.A(n_3232),
.Y(n_3418)
);

NAND2xp33_ASAP7_75t_L g3419 ( 
.A(n_3276),
.B(n_3176),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_L g3420 ( 
.A(n_3279),
.B(n_3120),
.Y(n_3420)
);

AOI22xp33_ASAP7_75t_L g3421 ( 
.A1(n_3283),
.A2(n_3150),
.B1(n_3073),
.B2(n_3089),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3198),
.B(n_3066),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_3269),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3245),
.B(n_3128),
.Y(n_3424)
);

INVx3_ASAP7_75t_L g3425 ( 
.A(n_3202),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3268),
.B(n_3071),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3262),
.Y(n_3427)
);

NAND2x1_ASAP7_75t_L g3428 ( 
.A(n_3240),
.B(n_3128),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3285),
.Y(n_3429)
);

INVxp67_ASAP7_75t_SL g3430 ( 
.A(n_3288),
.Y(n_3430)
);

BUFx3_ASAP7_75t_L g3431 ( 
.A(n_3291),
.Y(n_3431)
);

INVx3_ASAP7_75t_L g3432 ( 
.A(n_3202),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3272),
.Y(n_3433)
);

OR2x2_ASAP7_75t_L g3434 ( 
.A(n_3299),
.B(n_3090),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3302),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3377),
.B(n_3148),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_3195),
.Y(n_3437)
);

HB1xp67_ASAP7_75t_L g3438 ( 
.A(n_3336),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3190),
.B(n_3148),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3204),
.B(n_3170),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3223),
.B(n_3170),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3361),
.B(n_3179),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3206),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3306),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3226),
.B(n_3179),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3208),
.B(n_3152),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3207),
.Y(n_3447)
);

OAI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3264),
.A2(n_3183),
.B(n_2071),
.Y(n_3448)
);

BUFx12f_ASAP7_75t_L g3449 ( 
.A(n_3246),
.Y(n_3449)
);

AND3x1_ASAP7_75t_SL g3450 ( 
.A(n_3331),
.B(n_3145),
.C(n_926),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3212),
.Y(n_3451)
);

BUFx2_ASAP7_75t_L g3452 ( 
.A(n_3293),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3248),
.B(n_3286),
.Y(n_3453)
);

BUFx4f_ASAP7_75t_L g3454 ( 
.A(n_3272),
.Y(n_3454)
);

HB1xp67_ASAP7_75t_L g3455 ( 
.A(n_3400),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3275),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3297),
.B(n_2620),
.Y(n_3457)
);

BUFx12f_ASAP7_75t_L g3458 ( 
.A(n_3272),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3362),
.B(n_3241),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3322),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3329),
.Y(n_3461)
);

INVx3_ASAP7_75t_L g3462 ( 
.A(n_3201),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3348),
.Y(n_3463)
);

BUFx3_ASAP7_75t_L g3464 ( 
.A(n_3326),
.Y(n_3464)
);

AND2x4_ASAP7_75t_L g3465 ( 
.A(n_3300),
.B(n_3002),
.Y(n_3465)
);

BUFx2_ASAP7_75t_L g3466 ( 
.A(n_3367),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3244),
.B(n_2622),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3213),
.B(n_3284),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3290),
.B(n_2625),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3359),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3311),
.B(n_2625),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_R g3472 ( 
.A(n_3201),
.B(n_3139),
.Y(n_3472)
);

INVx2_ASAP7_75t_SL g3473 ( 
.A(n_3307),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3260),
.B(n_2628),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_3199),
.B(n_3002),
.Y(n_3475)
);

BUFx2_ASAP7_75t_L g3476 ( 
.A(n_3367),
.Y(n_3476)
);

INVx3_ASAP7_75t_L g3477 ( 
.A(n_3277),
.Y(n_3477)
);

INVxp67_ASAP7_75t_SL g3478 ( 
.A(n_3338),
.Y(n_3478)
);

BUFx6f_ASAP7_75t_L g3479 ( 
.A(n_3277),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3365),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3224),
.B(n_3216),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3360),
.Y(n_3482)
);

BUFx6f_ASAP7_75t_L g3483 ( 
.A(n_3277),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3369),
.Y(n_3484)
);

INVx4_ASAP7_75t_L g3485 ( 
.A(n_3295),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3368),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3342),
.B(n_2556),
.Y(n_3487)
);

INVx2_ASAP7_75t_SL g3488 ( 
.A(n_3251),
.Y(n_3488)
);

INVx3_ASAP7_75t_L g3489 ( 
.A(n_3295),
.Y(n_3489)
);

BUFx2_ASAP7_75t_L g3490 ( 
.A(n_3342),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3379),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3402),
.Y(n_3492)
);

A2O1A1Ixp33_ASAP7_75t_SL g3493 ( 
.A1(n_3258),
.A2(n_2556),
.B(n_2079),
.C(n_2082),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3339),
.A2(n_923),
.B1(n_927),
.B2(n_926),
.Y(n_3494)
);

INVx4_ASAP7_75t_L g3495 ( 
.A(n_3295),
.Y(n_3495)
);

BUFx3_ASAP7_75t_L g3496 ( 
.A(n_3282),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3354),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3227),
.B(n_934),
.Y(n_3498)
);

CKINVDCx5p33_ASAP7_75t_R g3499 ( 
.A(n_3191),
.Y(n_3499)
);

AND2x4_ASAP7_75t_L g3500 ( 
.A(n_3300),
.B(n_2628),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_3231),
.B(n_2956),
.Y(n_3501)
);

BUFx3_ASAP7_75t_L g3502 ( 
.A(n_3242),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3296),
.B(n_3399),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3385),
.Y(n_3504)
);

INVx4_ASAP7_75t_L g3505 ( 
.A(n_3385),
.Y(n_3505)
);

HB1xp67_ASAP7_75t_L g3506 ( 
.A(n_3346),
.Y(n_3506)
);

AND2x4_ASAP7_75t_L g3507 ( 
.A(n_3343),
.B(n_2658),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3214),
.Y(n_3508)
);

AND2x6_ASAP7_75t_L g3509 ( 
.A(n_3196),
.B(n_3281),
.Y(n_3509)
);

BUFx3_ASAP7_75t_L g3510 ( 
.A(n_3385),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3238),
.B(n_2658),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3217),
.B(n_934),
.Y(n_3512)
);

AND2x4_ASAP7_75t_L g3513 ( 
.A(n_3334),
.B(n_2056),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3328),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3397),
.Y(n_3515)
);

INVxp67_ASAP7_75t_L g3516 ( 
.A(n_3289),
.Y(n_3516)
);

HB1xp67_ASAP7_75t_L g3517 ( 
.A(n_3352),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3358),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3308),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3347),
.Y(n_3520)
);

CKINVDCx5p33_ASAP7_75t_R g3521 ( 
.A(n_3230),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3393),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3356),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3373),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3334),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3305),
.B(n_664),
.Y(n_3526)
);

OR2x6_ASAP7_75t_L g3527 ( 
.A(n_3193),
.B(n_2082),
.Y(n_3527)
);

AND2x4_ASAP7_75t_L g3528 ( 
.A(n_3345),
.B(n_2082),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3345),
.Y(n_3529)
);

AND2x4_ASAP7_75t_L g3530 ( 
.A(n_3341),
.B(n_3344),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3196),
.Y(n_3531)
);

INVx2_ASAP7_75t_SL g3532 ( 
.A(n_3370),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3378),
.Y(n_3533)
);

INVxp67_ASAP7_75t_L g3534 ( 
.A(n_3324),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3280),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3236),
.Y(n_3536)
);

BUFx6f_ASAP7_75t_L g3537 ( 
.A(n_3370),
.Y(n_3537)
);

BUFx4f_ASAP7_75t_L g3538 ( 
.A(n_3252),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3281),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3314),
.Y(n_3540)
);

AND2x2_ASAP7_75t_L g3541 ( 
.A(n_3225),
.B(n_665),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3349),
.Y(n_3542)
);

AND3x1_ASAP7_75t_SL g3543 ( 
.A(n_3273),
.B(n_940),
.C(n_937),
.Y(n_3543)
);

INVx3_ASAP7_75t_L g3544 ( 
.A(n_3392),
.Y(n_3544)
);

AOI221xp5_ASAP7_75t_L g3545 ( 
.A1(n_3255),
.A2(n_940),
.B1(n_942),
.B2(n_941),
.C(n_937),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3228),
.B(n_668),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3220),
.B(n_2956),
.Y(n_3547)
);

NOR2xp33_ASAP7_75t_L g3548 ( 
.A(n_3250),
.B(n_941),
.Y(n_3548)
);

AO22x1_ASAP7_75t_L g3549 ( 
.A1(n_3403),
.A2(n_1027),
.B1(n_946),
.B2(n_950),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3314),
.Y(n_3550)
);

AND2x6_ASAP7_75t_L g3551 ( 
.A(n_3317),
.B(n_2956),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3392),
.Y(n_3552)
);

AND3x2_ASAP7_75t_SL g3553 ( 
.A(n_3382),
.B(n_704),
.C(n_1062),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3239),
.B(n_3312),
.Y(n_3554)
);

AND2x4_ASAP7_75t_SL g3555 ( 
.A(n_3240),
.B(n_2303),
.Y(n_3555)
);

AOI22xp5_ASAP7_75t_SL g3556 ( 
.A1(n_3192),
.A2(n_946),
.B1(n_950),
.B2(n_942),
.Y(n_3556)
);

AND2x2_ASAP7_75t_L g3557 ( 
.A(n_3249),
.B(n_672),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3371),
.B(n_674),
.Y(n_3558)
);

AO22x1_ASAP7_75t_L g3559 ( 
.A1(n_3265),
.A2(n_962),
.B1(n_953),
.B2(n_957),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3315),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3252),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_SL g3562 ( 
.A(n_3382),
.B(n_3205),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3235),
.B(n_2097),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3215),
.B(n_2097),
.Y(n_3564)
);

INVx2_ASAP7_75t_SL g3565 ( 
.A(n_3309),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3383),
.B(n_2097),
.Y(n_3566)
);

CKINVDCx5p33_ASAP7_75t_R g3567 ( 
.A(n_3320),
.Y(n_3567)
);

INVx3_ASAP7_75t_L g3568 ( 
.A(n_3320),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3321),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3278),
.B(n_676),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3351),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_SL g3572 ( 
.A1(n_3253),
.A2(n_953),
.B1(n_957),
.B2(n_952),
.Y(n_3572)
);

INVxp67_ASAP7_75t_L g3573 ( 
.A(n_3304),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3243),
.B(n_2100),
.Y(n_3574)
);

OR2x6_ASAP7_75t_L g3575 ( 
.A(n_3221),
.B(n_2100),
.Y(n_3575)
);

BUFx6f_ASAP7_75t_L g3576 ( 
.A(n_3309),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3210),
.B(n_3247),
.Y(n_3577)
);

INVx3_ASAP7_75t_L g3578 ( 
.A(n_3337),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3332),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3257),
.B(n_677),
.Y(n_3580)
);

AND2x6_ASAP7_75t_SL g3581 ( 
.A(n_3258),
.B(n_952),
.Y(n_3581)
);

INVx3_ASAP7_75t_L g3582 ( 
.A(n_3388),
.Y(n_3582)
);

INVxp67_ASAP7_75t_SL g3583 ( 
.A(n_3380),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_3205),
.B(n_960),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3218),
.A2(n_2032),
.B(n_2029),
.Y(n_3585)
);

INVxp67_ASAP7_75t_L g3586 ( 
.A(n_3391),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3274),
.B(n_2100),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3219),
.Y(n_3588)
);

HB1xp67_ASAP7_75t_L g3589 ( 
.A(n_3355),
.Y(n_3589)
);

BUFx3_ASAP7_75t_L g3590 ( 
.A(n_3384),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3194),
.B(n_2109),
.Y(n_3591)
);

INVx1_ASAP7_75t_SL g3592 ( 
.A(n_3387),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_3364),
.B(n_2109),
.Y(n_3593)
);

INVx6_ASAP7_75t_L g3594 ( 
.A(n_3197),
.Y(n_3594)
);

AO22x1_ASAP7_75t_L g3595 ( 
.A1(n_3372),
.A2(n_1033),
.B1(n_962),
.B2(n_1024),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3353),
.Y(n_3596)
);

OAI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3234),
.A2(n_1024),
.B1(n_1027),
.B2(n_960),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3340),
.Y(n_3598)
);

OAI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3266),
.A2(n_1032),
.B1(n_1033),
.B2(n_1028),
.Y(n_3599)
);

BUFx2_ASAP7_75t_R g3600 ( 
.A(n_3327),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3200),
.B(n_2109),
.Y(n_3601)
);

INVx4_ASAP7_75t_L g3602 ( 
.A(n_3376),
.Y(n_3602)
);

AOI22x1_ASAP7_75t_L g3603 ( 
.A1(n_3233),
.A2(n_1032),
.B1(n_1028),
.B2(n_1786),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3351),
.Y(n_3604)
);

INVx3_ASAP7_75t_L g3605 ( 
.A(n_3267),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3381),
.Y(n_3606)
);

AND3x2_ASAP7_75t_SL g3607 ( 
.A(n_3313),
.B(n_4),
.C(n_5),
.Y(n_3607)
);

BUFx6f_ASAP7_75t_L g3608 ( 
.A(n_3363),
.Y(n_3608)
);

BUFx2_ASAP7_75t_L g3609 ( 
.A(n_3389),
.Y(n_3609)
);

OR2x2_ASAP7_75t_L g3610 ( 
.A(n_3310),
.B(n_2071),
.Y(n_3610)
);

NOR2xp33_ASAP7_75t_L g3611 ( 
.A(n_3319),
.B(n_678),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3209),
.B(n_1803),
.Y(n_3612)
);

BUFx6f_ASAP7_75t_L g3613 ( 
.A(n_3374),
.Y(n_3613)
);

NOR2xp33_ASAP7_75t_L g3614 ( 
.A(n_3375),
.B(n_679),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_3394),
.Y(n_3615)
);

A2O1A1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_3357),
.A2(n_2145),
.B(n_2150),
.C(n_2111),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3318),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3211),
.B(n_1803),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3396),
.Y(n_3619)
);

BUFx2_ASAP7_75t_L g3620 ( 
.A(n_3401),
.Y(n_3620)
);

AND3x1_ASAP7_75t_SL g3621 ( 
.A(n_3335),
.B(n_5),
.C(n_6),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3390),
.B(n_680),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3404),
.Y(n_3623)
);

BUFx2_ASAP7_75t_L g3624 ( 
.A(n_3409),
.Y(n_3624)
);

INVx2_ASAP7_75t_SL g3625 ( 
.A(n_3418),
.Y(n_3625)
);

INVx3_ASAP7_75t_L g3626 ( 
.A(n_3415),
.Y(n_3626)
);

CKINVDCx5p33_ASAP7_75t_R g3627 ( 
.A(n_3416),
.Y(n_3627)
);

BUFx6f_ASAP7_75t_L g3628 ( 
.A(n_3418),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3430),
.B(n_3287),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3427),
.Y(n_3630)
);

NOR4xp25_ASAP7_75t_SL g3631 ( 
.A(n_3562),
.B(n_3298),
.C(n_3303),
.D(n_3301),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_3406),
.B(n_3316),
.Y(n_3632)
);

OR2x6_ASAP7_75t_L g3633 ( 
.A(n_3594),
.B(n_3325),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3452),
.B(n_3292),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_SL g3635 ( 
.A(n_3406),
.B(n_3294),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3429),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3435),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3444),
.Y(n_3638)
);

AOI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_3420),
.A2(n_1803),
.B1(n_1826),
.B2(n_1804),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3470),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3482),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3484),
.Y(n_3642)
);

INVx3_ASAP7_75t_L g3643 ( 
.A(n_3415),
.Y(n_3643)
);

INVx2_ASAP7_75t_SL g3644 ( 
.A(n_3418),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3497),
.B(n_3261),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3417),
.Y(n_3646)
);

NAND2x1p5_ASAP7_75t_L g3647 ( 
.A(n_3538),
.B(n_3398),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3459),
.A2(n_3386),
.B(n_3330),
.Y(n_3648)
);

CKINVDCx11_ASAP7_75t_R g3649 ( 
.A(n_3449),
.Y(n_3649)
);

OAI22xp5_ASAP7_75t_SL g3650 ( 
.A1(n_3548),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_3650)
);

O2A1O1Ixp33_ASAP7_75t_L g3651 ( 
.A1(n_3494),
.A2(n_3333),
.B(n_2145),
.C(n_2150),
.Y(n_3651)
);

NOR2xp67_ASAP7_75t_L g3652 ( 
.A(n_3573),
.B(n_7),
.Y(n_3652)
);

OAI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3585),
.A2(n_2032),
.B(n_2029),
.Y(n_3653)
);

OR2x2_ASAP7_75t_L g3654 ( 
.A(n_3478),
.B(n_2071),
.Y(n_3654)
);

BUFx4f_ASAP7_75t_L g3655 ( 
.A(n_3462),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3453),
.B(n_8),
.Y(n_3656)
);

BUFx6f_ASAP7_75t_L g3657 ( 
.A(n_3479),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3536),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3455),
.Y(n_3659)
);

AND2x2_ASAP7_75t_L g3660 ( 
.A(n_3506),
.B(n_9),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3517),
.B(n_10),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3556),
.A2(n_2111),
.B(n_2150),
.C(n_2145),
.Y(n_3662)
);

O2A1O1Ixp33_ASAP7_75t_L g3663 ( 
.A1(n_3494),
.A2(n_2111),
.B(n_2188),
.C(n_2175),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3437),
.Y(n_3664)
);

INVx5_ASAP7_75t_L g3665 ( 
.A(n_3594),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3453),
.B(n_3520),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3535),
.Y(n_3667)
);

INVx2_ASAP7_75t_SL g3668 ( 
.A(n_3423),
.Y(n_3668)
);

O2A1O1Ixp33_ASAP7_75t_L g3669 ( 
.A1(n_3412),
.A2(n_2175),
.B(n_2210),
.C(n_2188),
.Y(n_3669)
);

INVx1_ASAP7_75t_SL g3670 ( 
.A(n_3499),
.Y(n_3670)
);

AND3x2_ASAP7_75t_L g3671 ( 
.A(n_3584),
.B(n_3475),
.C(n_3516),
.Y(n_3671)
);

O2A1O1Ixp33_ASAP7_75t_L g3672 ( 
.A1(n_3412),
.A2(n_2175),
.B(n_2210),
.C(n_2188),
.Y(n_3672)
);

HB1xp67_ASAP7_75t_L g3673 ( 
.A(n_3490),
.Y(n_3673)
);

BUFx6f_ASAP7_75t_L g3674 ( 
.A(n_3479),
.Y(n_3674)
);

INVx3_ASAP7_75t_L g3675 ( 
.A(n_3525),
.Y(n_3675)
);

INVx4_ASAP7_75t_L g3676 ( 
.A(n_3567),
.Y(n_3676)
);

INVxp67_ASAP7_75t_L g3677 ( 
.A(n_3496),
.Y(n_3677)
);

A2O1A1Ixp33_ASAP7_75t_SL g3678 ( 
.A1(n_3614),
.A2(n_2210),
.B(n_2229),
.C(n_2237),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_3459),
.A2(n_2229),
.B(n_2303),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3443),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3502),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3491),
.Y(n_3682)
);

NOR2x1_ASAP7_75t_L g3683 ( 
.A(n_3481),
.B(n_2229),
.Y(n_3683)
);

O2A1O1Ixp33_ASAP7_75t_L g3684 ( 
.A1(n_3419),
.A2(n_2237),
.B(n_2298),
.C(n_2032),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3522),
.B(n_10),
.Y(n_3685)
);

A2O1A1Ixp33_ASAP7_75t_SL g3686 ( 
.A1(n_3622),
.A2(n_2298),
.B(n_2237),
.C(n_13),
.Y(n_3686)
);

INVx3_ASAP7_75t_L g3687 ( 
.A(n_3537),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3447),
.Y(n_3688)
);

INVxp67_ASAP7_75t_SL g3689 ( 
.A(n_3436),
.Y(n_3689)
);

INVx2_ASAP7_75t_SL g3690 ( 
.A(n_3431),
.Y(n_3690)
);

AND3x1_ASAP7_75t_L g3691 ( 
.A(n_3512),
.B(n_11),
.C(n_12),
.Y(n_3691)
);

INVx4_ASAP7_75t_L g3692 ( 
.A(n_3462),
.Y(n_3692)
);

OAI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3556),
.A2(n_2298),
.B1(n_1803),
.B2(n_1826),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3451),
.Y(n_3694)
);

CKINVDCx5p33_ASAP7_75t_R g3695 ( 
.A(n_3521),
.Y(n_3695)
);

OAI22xp5_ASAP7_75t_SL g3696 ( 
.A1(n_3446),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3523),
.Y(n_3697)
);

BUFx3_ASAP7_75t_L g3698 ( 
.A(n_3464),
.Y(n_3698)
);

BUFx4f_ASAP7_75t_L g3699 ( 
.A(n_3458),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3456),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3468),
.B(n_14),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3460),
.Y(n_3702)
);

AND2x4_ASAP7_75t_L g3703 ( 
.A(n_3530),
.B(n_693),
.Y(n_3703)
);

BUFx12f_ASAP7_75t_L g3704 ( 
.A(n_3488),
.Y(n_3704)
);

AOI22xp33_ASAP7_75t_L g3705 ( 
.A1(n_3572),
.A2(n_1804),
.B1(n_1827),
.B2(n_1826),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3461),
.Y(n_3706)
);

INVx3_ASAP7_75t_L g3707 ( 
.A(n_3529),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3560),
.B(n_15),
.Y(n_3708)
);

O2A1O1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3577),
.A2(n_19),
.B(n_16),
.C(n_18),
.Y(n_3709)
);

OAI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_3503),
.A2(n_1804),
.B1(n_1827),
.B2(n_1826),
.Y(n_3710)
);

INVx5_ASAP7_75t_L g3711 ( 
.A(n_3613),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3518),
.B(n_18),
.Y(n_3712)
);

INVx5_ASAP7_75t_L g3713 ( 
.A(n_3613),
.Y(n_3713)
);

OAI21xp33_ASAP7_75t_L g3714 ( 
.A1(n_3545),
.A2(n_1827),
.B(n_1804),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3463),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_SL g3716 ( 
.A(n_3538),
.B(n_1827),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3533),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3440),
.B(n_19),
.Y(n_3718)
);

HB1xp67_ASAP7_75t_L g3719 ( 
.A(n_3438),
.Y(n_3719)
);

O2A1O1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3599),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3441),
.B(n_20),
.Y(n_3721)
);

A2O1A1Ixp33_ASAP7_75t_L g3722 ( 
.A1(n_3611),
.A2(n_1829),
.B(n_24),
.C(n_21),
.Y(n_3722)
);

AND2x4_ASAP7_75t_L g3723 ( 
.A(n_3530),
.B(n_681),
.Y(n_3723)
);

NOR2x1_ASAP7_75t_SL g3724 ( 
.A(n_3588),
.B(n_1223),
.Y(n_3724)
);

AND2x4_ASAP7_75t_SL g3725 ( 
.A(n_3414),
.B(n_2303),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3436),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3434),
.B(n_23),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3480),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3486),
.Y(n_3729)
);

BUFx6f_ASAP7_75t_L g3730 ( 
.A(n_3479),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_SL g3731 ( 
.A1(n_3572),
.A2(n_1829),
.B1(n_1223),
.B2(n_25),
.Y(n_3731)
);

INVx3_ASAP7_75t_L g3732 ( 
.A(n_3537),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3492),
.Y(n_3733)
);

INVx5_ASAP7_75t_L g3734 ( 
.A(n_3613),
.Y(n_3734)
);

BUFx12f_ASAP7_75t_L g3735 ( 
.A(n_3473),
.Y(n_3735)
);

INVx1_ASAP7_75t_SL g3736 ( 
.A(n_3510),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3445),
.B(n_23),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3515),
.Y(n_3738)
);

NOR3xp33_ASAP7_75t_L g3739 ( 
.A(n_3559),
.B(n_24),
.C(n_25),
.Y(n_3739)
);

INVx2_ASAP7_75t_SL g3740 ( 
.A(n_3483),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3442),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3514),
.B(n_27),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3407),
.B(n_27),
.Y(n_3743)
);

OAI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3534),
.A2(n_1829),
.B1(n_2310),
.B2(n_2309),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3554),
.A2(n_2310),
.B(n_2309),
.Y(n_3745)
);

HB1xp67_ASAP7_75t_L g3746 ( 
.A(n_3519),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3407),
.B(n_28),
.Y(n_3747)
);

NOR2xp33_ASAP7_75t_L g3748 ( 
.A(n_3410),
.B(n_3541),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3442),
.Y(n_3749)
);

OR2x6_ASAP7_75t_L g3750 ( 
.A(n_3578),
.B(n_1829),
.Y(n_3750)
);

A2O1A1Ixp33_ASAP7_75t_L g3751 ( 
.A1(n_3558),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3531),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3466),
.B(n_29),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3408),
.B(n_31),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3554),
.A2(n_2310),
.B(n_2309),
.Y(n_3755)
);

NOR2xp33_ASAP7_75t_L g3756 ( 
.A(n_3546),
.B(n_31),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3408),
.B(n_33),
.Y(n_3757)
);

BUFx2_ASAP7_75t_SL g3758 ( 
.A(n_3509),
.Y(n_3758)
);

INVx6_ASAP7_75t_L g3759 ( 
.A(n_3483),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3426),
.B(n_33),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_3498),
.B(n_34),
.Y(n_3761)
);

HB1xp67_ASAP7_75t_L g3762 ( 
.A(n_3596),
.Y(n_3762)
);

INVx3_ASAP7_75t_SL g3763 ( 
.A(n_3411),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3421),
.A2(n_2309),
.B1(n_2310),
.B2(n_1223),
.Y(n_3764)
);

AOI221xp5_ASAP7_75t_L g3765 ( 
.A1(n_3549),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_3765)
);

BUFx8_ASAP7_75t_L g3766 ( 
.A(n_3537),
.Y(n_3766)
);

INVx6_ASAP7_75t_L g3767 ( 
.A(n_3483),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3508),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3539),
.Y(n_3769)
);

HB1xp67_ASAP7_75t_L g3770 ( 
.A(n_3596),
.Y(n_3770)
);

BUFx4f_ASAP7_75t_SL g3771 ( 
.A(n_3477),
.Y(n_3771)
);

NOR2x1_ASAP7_75t_R g3772 ( 
.A(n_3405),
.B(n_37),
.Y(n_3772)
);

HB1xp67_ASAP7_75t_L g3773 ( 
.A(n_3596),
.Y(n_3773)
);

CKINVDCx5p33_ASAP7_75t_R g3774 ( 
.A(n_3405),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3426),
.B(n_35),
.Y(n_3775)
);

BUFx2_ASAP7_75t_L g3776 ( 
.A(n_3476),
.Y(n_3776)
);

OAI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3607),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3540),
.Y(n_3778)
);

OR2x6_ASAP7_75t_L g3779 ( 
.A(n_3578),
.B(n_1712),
.Y(n_3779)
);

AND2x4_ASAP7_75t_L g3780 ( 
.A(n_3465),
.B(n_689),
.Y(n_3780)
);

A2O1A1Ixp33_ASAP7_75t_L g3781 ( 
.A1(n_3599),
.A2(n_3493),
.B(n_3609),
.C(n_3570),
.Y(n_3781)
);

BUFx6f_ASAP7_75t_L g3782 ( 
.A(n_3454),
.Y(n_3782)
);

AO21x2_ASAP7_75t_L g3783 ( 
.A1(n_3564),
.A2(n_39),
.B(n_41),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3439),
.B(n_43),
.Y(n_3784)
);

BUFx4f_ASAP7_75t_SL g3785 ( 
.A(n_3477),
.Y(n_3785)
);

OR2x6_ASAP7_75t_L g3786 ( 
.A(n_3527),
.B(n_1712),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3583),
.A2(n_1740),
.B(n_1735),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3569),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3550),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3413),
.B(n_43),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3612),
.A2(n_1740),
.B(n_1735),
.Y(n_3791)
);

AOI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3563),
.A2(n_1740),
.B(n_1735),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3542),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3590),
.A2(n_1740),
.B1(n_1735),
.B2(n_46),
.Y(n_3794)
);

CKINVDCx11_ASAP7_75t_R g3795 ( 
.A(n_3552),
.Y(n_3795)
);

OR2x6_ASAP7_75t_L g3796 ( 
.A(n_3527),
.B(n_682),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3474),
.Y(n_3797)
);

AND3x1_ASAP7_75t_SL g3798 ( 
.A(n_3450),
.B(n_44),
.C(n_45),
.Y(n_3798)
);

NOR2xp33_ASAP7_75t_L g3799 ( 
.A(n_3501),
.B(n_46),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3524),
.Y(n_3800)
);

AOI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_3563),
.A2(n_684),
.B(n_683),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_R g3802 ( 
.A(n_3454),
.B(n_685),
.Y(n_3802)
);

A2O1A1Ixp33_ASAP7_75t_L g3803 ( 
.A1(n_3589),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_3803)
);

OAI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3620),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_3804)
);

OR2x2_ASAP7_75t_L g3805 ( 
.A(n_3571),
.B(n_53),
.Y(n_3805)
);

AOI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3592),
.A2(n_688),
.B(n_687),
.Y(n_3806)
);

OR2x2_ASAP7_75t_L g3807 ( 
.A(n_3610),
.B(n_53),
.Y(n_3807)
);

OR2x2_ASAP7_75t_L g3808 ( 
.A(n_3582),
.B(n_54),
.Y(n_3808)
);

AND2x4_ASAP7_75t_L g3809 ( 
.A(n_3465),
.B(n_697),
.Y(n_3809)
);

OAI22xp5_ASAP7_75t_L g3810 ( 
.A1(n_3600),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3526),
.B(n_58),
.Y(n_3811)
);

INVx3_ASAP7_75t_L g3812 ( 
.A(n_3485),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3474),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3606),
.Y(n_3814)
);

CKINVDCx5p33_ASAP7_75t_R g3815 ( 
.A(n_3472),
.Y(n_3815)
);

INVx3_ASAP7_75t_L g3816 ( 
.A(n_3485),
.Y(n_3816)
);

BUFx6f_ASAP7_75t_SL g3817 ( 
.A(n_3495),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3582),
.B(n_3487),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3500),
.Y(n_3819)
);

NAND2x2_ASAP7_75t_L g3820 ( 
.A(n_3565),
.B(n_60),
.Y(n_3820)
);

O2A1O1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3547),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3617),
.Y(n_3822)
);

BUFx2_ASAP7_75t_SL g3823 ( 
.A(n_3509),
.Y(n_3823)
);

BUFx2_ASAP7_75t_L g3824 ( 
.A(n_3509),
.Y(n_3824)
);

BUFx6f_ASAP7_75t_L g3825 ( 
.A(n_3489),
.Y(n_3825)
);

OR2x2_ASAP7_75t_L g3826 ( 
.A(n_3413),
.B(n_61),
.Y(n_3826)
);

INVxp67_ASAP7_75t_L g3827 ( 
.A(n_3489),
.Y(n_3827)
);

INVx3_ASAP7_75t_L g3828 ( 
.A(n_3495),
.Y(n_3828)
);

HB1xp67_ASAP7_75t_L g3829 ( 
.A(n_3586),
.Y(n_3829)
);

NOR2xp33_ASAP7_75t_L g3830 ( 
.A(n_3411),
.B(n_62),
.Y(n_3830)
);

OR2x6_ASAP7_75t_L g3831 ( 
.A(n_3527),
.B(n_695),
.Y(n_3831)
);

BUFx3_ASAP7_75t_L g3832 ( 
.A(n_3504),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3500),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3592),
.A2(n_698),
.B(n_63),
.Y(n_3834)
);

INVx4_ASAP7_75t_L g3835 ( 
.A(n_3576),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3511),
.Y(n_3836)
);

BUFx12f_ASAP7_75t_L g3837 ( 
.A(n_3505),
.Y(n_3837)
);

OR2x6_ASAP7_75t_L g3838 ( 
.A(n_3576),
.B(n_63),
.Y(n_3838)
);

AND2x4_ASAP7_75t_L g3839 ( 
.A(n_3561),
.B(n_64),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3507),
.B(n_64),
.Y(n_3840)
);

NOR2xp33_ASAP7_75t_SL g3841 ( 
.A(n_3505),
.B(n_65),
.Y(n_3841)
);

AOI22x1_ASAP7_75t_L g3842 ( 
.A1(n_3602),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3471),
.B(n_66),
.Y(n_3843)
);

A2O1A1Ixp33_ASAP7_75t_L g3844 ( 
.A1(n_3605),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_3844)
);

OR2x6_ASAP7_75t_L g3845 ( 
.A(n_3576),
.B(n_68),
.Y(n_3845)
);

A2O1A1Ixp33_ASAP7_75t_L g3846 ( 
.A1(n_3605),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3511),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_3425),
.B(n_72),
.Y(n_3848)
);

INVx3_ASAP7_75t_L g3849 ( 
.A(n_3504),
.Y(n_3849)
);

INVx3_ASAP7_75t_L g3850 ( 
.A(n_3425),
.Y(n_3850)
);

AND2x4_ASAP7_75t_L g3851 ( 
.A(n_3507),
.B(n_72),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3658),
.Y(n_3852)
);

AOI22xp33_ASAP7_75t_L g3853 ( 
.A1(n_3777),
.A2(n_3650),
.B1(n_3739),
.B2(n_3696),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3648),
.A2(n_3684),
.B(n_3686),
.Y(n_3854)
);

INVx1_ASAP7_75t_SL g3855 ( 
.A(n_3795),
.Y(n_3855)
);

AOI22xp5_ASAP7_75t_L g3856 ( 
.A1(n_3810),
.A2(n_3691),
.B1(n_3841),
.B2(n_3765),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3714),
.A2(n_3422),
.B(n_3595),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3671),
.A2(n_3621),
.B1(n_3597),
.B2(n_3424),
.Y(n_3858)
);

AOI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3635),
.A2(n_3618),
.B(n_3457),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3689),
.B(n_3587),
.Y(n_3860)
);

BUFx3_ASAP7_75t_L g3861 ( 
.A(n_3735),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3800),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3624),
.B(n_3432),
.Y(n_3863)
);

AOI22xp33_ASAP7_75t_L g3864 ( 
.A1(n_3842),
.A2(n_3603),
.B1(n_3602),
.B2(n_3580),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3667),
.B(n_3587),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3623),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3630),
.Y(n_3867)
);

CKINVDCx20_ASAP7_75t_R g3868 ( 
.A(n_3627),
.Y(n_3868)
);

BUFx6f_ASAP7_75t_L g3869 ( 
.A(n_3628),
.Y(n_3869)
);

CKINVDCx5p33_ASAP7_75t_R g3870 ( 
.A(n_3695),
.Y(n_3870)
);

O2A1O1Ixp33_ASAP7_75t_SL g3871 ( 
.A1(n_3751),
.A2(n_3532),
.B(n_3553),
.C(n_3432),
.Y(n_3871)
);

BUFx2_ASAP7_75t_L g3872 ( 
.A(n_3626),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3636),
.Y(n_3873)
);

AND2x4_ASAP7_75t_L g3874 ( 
.A(n_3626),
.B(n_3575),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3637),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3638),
.Y(n_3876)
);

OR2x6_ASAP7_75t_L g3877 ( 
.A(n_3758),
.B(n_3575),
.Y(n_3877)
);

BUFx8_ASAP7_75t_SL g3878 ( 
.A(n_3774),
.Y(n_3878)
);

NAND2x1_ASAP7_75t_L g3879 ( 
.A(n_3726),
.B(n_3575),
.Y(n_3879)
);

INVx1_ASAP7_75t_SL g3880 ( 
.A(n_3670),
.Y(n_3880)
);

AND2x4_ASAP7_75t_L g3881 ( 
.A(n_3643),
.B(n_3608),
.Y(n_3881)
);

AOI22xp33_ASAP7_75t_SL g3882 ( 
.A1(n_3665),
.A2(n_3557),
.B1(n_3608),
.B2(n_3551),
.Y(n_3882)
);

CKINVDCx5p33_ASAP7_75t_R g3883 ( 
.A(n_3649),
.Y(n_3883)
);

NOR2xp33_ASAP7_75t_L g3884 ( 
.A(n_3748),
.B(n_3433),
.Y(n_3884)
);

INVx3_ASAP7_75t_L g3885 ( 
.A(n_3628),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3640),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3642),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3646),
.B(n_3604),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3719),
.B(n_3457),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3641),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3673),
.B(n_3598),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3643),
.B(n_3433),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3776),
.B(n_3568),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3659),
.B(n_3818),
.Y(n_3894)
);

CKINVDCx11_ASAP7_75t_R g3895 ( 
.A(n_3704),
.Y(n_3895)
);

INVx2_ASAP7_75t_SL g3896 ( 
.A(n_3628),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_SL g3897 ( 
.A(n_3815),
.B(n_3509),
.Y(n_3897)
);

BUFx4f_ASAP7_75t_L g3898 ( 
.A(n_3782),
.Y(n_3898)
);

INVx3_ASAP7_75t_L g3899 ( 
.A(n_3698),
.Y(n_3899)
);

BUFx8_ASAP7_75t_L g3900 ( 
.A(n_3817),
.Y(n_3900)
);

BUFx2_ASAP7_75t_L g3901 ( 
.A(n_3762),
.Y(n_3901)
);

CKINVDCx11_ASAP7_75t_R g3902 ( 
.A(n_3837),
.Y(n_3902)
);

INVx4_ASAP7_75t_SL g3903 ( 
.A(n_3838),
.Y(n_3903)
);

NAND3xp33_ASAP7_75t_L g3904 ( 
.A(n_3709),
.B(n_3608),
.C(n_3591),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3819),
.B(n_3568),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3741),
.B(n_3564),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3749),
.B(n_3601),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3746),
.B(n_3697),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3793),
.Y(n_3909)
);

HB1xp67_ASAP7_75t_L g3910 ( 
.A(n_3645),
.Y(n_3910)
);

OR2x2_ASAP7_75t_L g3911 ( 
.A(n_3797),
.B(n_3574),
.Y(n_3911)
);

BUFx4f_ASAP7_75t_SL g3912 ( 
.A(n_3766),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3717),
.Y(n_3913)
);

AND2x4_ASAP7_75t_L g3914 ( 
.A(n_3833),
.B(n_3591),
.Y(n_3914)
);

OAI221xp5_ASAP7_75t_L g3915 ( 
.A1(n_3731),
.A2(n_3543),
.B1(n_3544),
.B2(n_3428),
.C(n_3601),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3814),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3632),
.A2(n_3448),
.B(n_3574),
.Y(n_3917)
);

INVx3_ASAP7_75t_L g3918 ( 
.A(n_3825),
.Y(n_3918)
);

INVx5_ASAP7_75t_L g3919 ( 
.A(n_3633),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3682),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3788),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3770),
.B(n_3448),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3666),
.B(n_3471),
.Y(n_3923)
);

AOI22xp5_ASAP7_75t_L g3924 ( 
.A1(n_3665),
.A2(n_3551),
.B1(n_3513),
.B2(n_3528),
.Y(n_3924)
);

AOI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3796),
.A2(n_3616),
.B(n_3566),
.Y(n_3925)
);

CKINVDCx8_ASAP7_75t_R g3926 ( 
.A(n_3665),
.Y(n_3926)
);

CKINVDCx5p33_ASAP7_75t_R g3927 ( 
.A(n_3766),
.Y(n_3927)
);

NOR2xp33_ASAP7_75t_L g3928 ( 
.A(n_3676),
.B(n_3677),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3768),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3822),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3829),
.B(n_3615),
.Y(n_3931)
);

INVx4_ASAP7_75t_L g3932 ( 
.A(n_3676),
.Y(n_3932)
);

O2A1O1Ixp33_ASAP7_75t_L g3933 ( 
.A1(n_3803),
.A2(n_3579),
.B(n_3544),
.C(n_3566),
.Y(n_3933)
);

OAI22xp5_ASAP7_75t_L g3934 ( 
.A1(n_3722),
.A2(n_3593),
.B1(n_3528),
.B2(n_3513),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3773),
.B(n_3619),
.Y(n_3935)
);

INVxp67_ASAP7_75t_SL g3936 ( 
.A(n_3813),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3752),
.Y(n_3937)
);

BUFx2_ASAP7_75t_L g3938 ( 
.A(n_3824),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3733),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3664),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3836),
.B(n_3467),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3796),
.A2(n_3467),
.B(n_3469),
.Y(n_3942)
);

INVx4_ASAP7_75t_L g3943 ( 
.A(n_3657),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3847),
.B(n_3469),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3680),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3681),
.B(n_3593),
.Y(n_3946)
);

INVx3_ASAP7_75t_L g3947 ( 
.A(n_3825),
.Y(n_3947)
);

BUFx3_ASAP7_75t_L g3948 ( 
.A(n_3625),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3820),
.A2(n_3551),
.B1(n_3581),
.B2(n_3555),
.Y(n_3949)
);

NOR2xp33_ASAP7_75t_L g3950 ( 
.A(n_3756),
.B(n_73),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3831),
.A2(n_3629),
.B(n_3678),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_3718),
.B(n_73),
.Y(n_3952)
);

INVx3_ASAP7_75t_L g3953 ( 
.A(n_3825),
.Y(n_3953)
);

BUFx6f_ASAP7_75t_L g3954 ( 
.A(n_3657),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3831),
.A2(n_3581),
.B(n_3551),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3634),
.B(n_74),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3807),
.B(n_74),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3688),
.B(n_75),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3711),
.A2(n_75),
.B(n_76),
.Y(n_3959)
);

OAI21xp33_ASAP7_75t_L g3960 ( 
.A1(n_3844),
.A2(n_76),
.B(n_77),
.Y(n_3960)
);

BUFx10_ASAP7_75t_L g3961 ( 
.A(n_3838),
.Y(n_3961)
);

OR2x6_ASAP7_75t_L g3962 ( 
.A(n_3758),
.B(n_78),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3694),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_3711),
.B(n_78),
.Y(n_3964)
);

CKINVDCx5p33_ASAP7_75t_R g3965 ( 
.A(n_3644),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_SL g3966 ( 
.A(n_3711),
.B(n_79),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3769),
.Y(n_3967)
);

AND2x4_ASAP7_75t_L g3968 ( 
.A(n_3835),
.B(n_79),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3668),
.B(n_641),
.Y(n_3969)
);

AOI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3761),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3736),
.B(n_642),
.Y(n_3971)
);

OAI22xp5_ASAP7_75t_L g3972 ( 
.A1(n_3846),
.A2(n_83),
.B1(n_80),
.B2(n_81),
.Y(n_3972)
);

INVx2_ASAP7_75t_SL g3973 ( 
.A(n_3759),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3713),
.A2(n_83),
.B(n_84),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3700),
.Y(n_3975)
);

OR2x6_ASAP7_75t_SL g3976 ( 
.A(n_3805),
.B(n_84),
.Y(n_3976)
);

AND2x4_ASAP7_75t_L g3977 ( 
.A(n_3835),
.B(n_3778),
.Y(n_3977)
);

CKINVDCx5p33_ASAP7_75t_R g3978 ( 
.A(n_3771),
.Y(n_3978)
);

AOI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3713),
.A2(n_3734),
.B(n_3631),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3789),
.Y(n_3980)
);

OR2x2_ASAP7_75t_L g3981 ( 
.A(n_3738),
.B(n_85),
.Y(n_3981)
);

INVx1_ASAP7_75t_SL g3982 ( 
.A(n_3690),
.Y(n_3982)
);

INVx3_ASAP7_75t_L g3983 ( 
.A(n_3832),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3702),
.Y(n_3984)
);

INVx4_ASAP7_75t_L g3985 ( 
.A(n_3657),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3675),
.Y(n_3986)
);

NAND3xp33_ASAP7_75t_L g3987 ( 
.A(n_3834),
.B(n_85),
.C(n_86),
.Y(n_3987)
);

CKINVDCx5p33_ASAP7_75t_R g3988 ( 
.A(n_3785),
.Y(n_3988)
);

CKINVDCx20_ASAP7_75t_R g3989 ( 
.A(n_3699),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3706),
.Y(n_3990)
);

AOI22xp5_ASAP7_75t_L g3991 ( 
.A1(n_3799),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3633),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3715),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3763),
.B(n_652),
.Y(n_3994)
);

CKINVDCx20_ASAP7_75t_R g3995 ( 
.A(n_3655),
.Y(n_3995)
);

BUFx6f_ASAP7_75t_L g3996 ( 
.A(n_3674),
.Y(n_3996)
);

BUFx6f_ASAP7_75t_L g3997 ( 
.A(n_3674),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3675),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3707),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3728),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3729),
.Y(n_4001)
);

AOI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3798),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_4002)
);

NAND3xp33_ASAP7_75t_L g4003 ( 
.A(n_3720),
.B(n_93),
.C(n_94),
.Y(n_4003)
);

INVx2_ASAP7_75t_SL g4004 ( 
.A(n_3759),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3713),
.B(n_3734),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3707),
.Y(n_4006)
);

NOR2xp33_ASAP7_75t_L g4007 ( 
.A(n_3721),
.B(n_95),
.Y(n_4007)
);

BUFx6f_ASAP7_75t_L g4008 ( 
.A(n_3674),
.Y(n_4008)
);

AND2x4_ASAP7_75t_L g4009 ( 
.A(n_3827),
.B(n_95),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3705),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4010)
);

AND2x4_ASAP7_75t_L g4011 ( 
.A(n_3692),
.B(n_96),
.Y(n_4011)
);

OR2x6_ASAP7_75t_L g4012 ( 
.A(n_3823),
.B(n_97),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3849),
.Y(n_4013)
);

INVx3_ASAP7_75t_L g4014 ( 
.A(n_3767),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3660),
.B(n_644),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3737),
.B(n_100),
.Y(n_4016)
);

AOI22xp33_ASAP7_75t_L g4017 ( 
.A1(n_3811),
.A2(n_104),
.B1(n_101),
.B2(n_103),
.Y(n_4017)
);

NOR2x1_ASAP7_75t_L g4018 ( 
.A(n_3783),
.B(n_101),
.Y(n_4018)
);

AOI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_3804),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_4019)
);

INVx5_ASAP7_75t_L g4020 ( 
.A(n_3845),
.Y(n_4020)
);

AO32x2_ASAP7_75t_L g4021 ( 
.A1(n_3740),
.A2(n_108),
.A3(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_4021)
);

AND2x4_ASAP7_75t_SL g4022 ( 
.A(n_3782),
.B(n_107),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3826),
.B(n_108),
.Y(n_4023)
);

INVx3_ASAP7_75t_L g4024 ( 
.A(n_3767),
.Y(n_4024)
);

O2A1O1Ixp33_ASAP7_75t_L g4025 ( 
.A1(n_3821),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_3734),
.A2(n_112),
.B(n_113),
.Y(n_4026)
);

OR2x6_ASAP7_75t_L g4027 ( 
.A(n_3823),
.B(n_112),
.Y(n_4027)
);

BUFx2_ASAP7_75t_SL g4028 ( 
.A(n_3652),
.Y(n_4028)
);

BUFx2_ASAP7_75t_L g4029 ( 
.A(n_3692),
.Y(n_4029)
);

AOI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3794),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3808),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3840),
.A2(n_3851),
.B1(n_3845),
.B2(n_3703),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3654),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_L g4034 ( 
.A1(n_3853),
.A2(n_3987),
.B1(n_3960),
.B2(n_4003),
.Y(n_4034)
);

OAI21x1_ASAP7_75t_L g4035 ( 
.A1(n_3917),
.A2(n_3755),
.B(n_3745),
.Y(n_4035)
);

AND2x4_ASAP7_75t_L g4036 ( 
.A(n_3938),
.B(n_3786),
.Y(n_4036)
);

OAI21x1_ASAP7_75t_L g4037 ( 
.A1(n_3859),
.A2(n_3792),
.B(n_3679),
.Y(n_4037)
);

AO21x2_ASAP7_75t_L g4038 ( 
.A1(n_3979),
.A2(n_3854),
.B(n_3906),
.Y(n_4038)
);

BUFx8_ASAP7_75t_L g4039 ( 
.A(n_3971),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3936),
.B(n_3843),
.Y(n_4040)
);

O2A1O1Ixp33_ASAP7_75t_SL g4041 ( 
.A1(n_3964),
.A2(n_3781),
.B(n_3662),
.C(n_3656),
.Y(n_4041)
);

OAI21x1_ASAP7_75t_L g4042 ( 
.A1(n_3951),
.A2(n_3787),
.B(n_3653),
.Y(n_4042)
);

OAI21x1_ASAP7_75t_L g4043 ( 
.A1(n_3925),
.A2(n_3791),
.B(n_3647),
.Y(n_4043)
);

BUFx3_ASAP7_75t_L g4044 ( 
.A(n_3878),
.Y(n_4044)
);

OAI21x1_ASAP7_75t_L g4045 ( 
.A1(n_3879),
.A2(n_3801),
.B(n_3683),
.Y(n_4045)
);

O2A1O1Ixp33_ASAP7_75t_L g4046 ( 
.A1(n_4025),
.A2(n_3693),
.B(n_3701),
.C(n_3784),
.Y(n_4046)
);

CKINVDCx11_ASAP7_75t_R g4047 ( 
.A(n_3868),
.Y(n_4047)
);

AOI22xp5_ASAP7_75t_L g4048 ( 
.A1(n_3856),
.A2(n_3851),
.B1(n_3840),
.B2(n_3703),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_3870),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3852),
.Y(n_4050)
);

OAI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3904),
.A2(n_3806),
.B(n_3639),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3909),
.Y(n_4052)
);

OAI21x1_ASAP7_75t_L g4053 ( 
.A1(n_3933),
.A2(n_3710),
.B(n_3744),
.Y(n_4053)
);

OAI21x1_ASAP7_75t_L g4054 ( 
.A1(n_3942),
.A2(n_3651),
.B(n_3672),
.Y(n_4054)
);

INVx4_ASAP7_75t_L g4055 ( 
.A(n_3912),
.Y(n_4055)
);

AOI21xp5_ASAP7_75t_R g4056 ( 
.A1(n_3972),
.A2(n_3839),
.B(n_3723),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_4002),
.A2(n_3747),
.B1(n_3743),
.B2(n_3754),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_3932),
.B(n_3727),
.Y(n_4058)
);

BUFx6f_ASAP7_75t_L g4059 ( 
.A(n_3926),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3910),
.B(n_3757),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3921),
.Y(n_4061)
);

AO21x2_ASAP7_75t_L g4062 ( 
.A1(n_3860),
.A2(n_3724),
.B(n_3760),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_4029),
.B(n_3786),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_L g4064 ( 
.A1(n_3950),
.A2(n_3723),
.B1(n_3802),
.B2(n_3780),
.Y(n_4064)
);

AND2x4_ASAP7_75t_L g4065 ( 
.A(n_3901),
.B(n_3687),
.Y(n_4065)
);

OAI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_3976),
.A2(n_3790),
.B1(n_3775),
.B2(n_3708),
.Y(n_4066)
);

O2A1O1Ixp33_ASAP7_75t_SL g4067 ( 
.A1(n_3966),
.A2(n_3712),
.B(n_3742),
.C(n_3716),
.Y(n_4067)
);

OA21x2_ASAP7_75t_L g4068 ( 
.A1(n_3929),
.A2(n_3930),
.B(n_3916),
.Y(n_4068)
);

CKINVDCx14_ASAP7_75t_R g4069 ( 
.A(n_3883),
.Y(n_4069)
);

AND2x4_ASAP7_75t_L g4070 ( 
.A(n_3977),
.B(n_3874),
.Y(n_4070)
);

INVx3_ASAP7_75t_SL g4071 ( 
.A(n_3927),
.Y(n_4071)
);

OAI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_4020),
.A2(n_3839),
.B1(n_3685),
.B2(n_3764),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_L g4073 ( 
.A1(n_3955),
.A2(n_3669),
.B(n_3812),
.Y(n_4073)
);

OAI21x1_ASAP7_75t_L g4074 ( 
.A1(n_3907),
.A2(n_3828),
.B(n_3816),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3872),
.B(n_3894),
.Y(n_4075)
);

AND2x4_ASAP7_75t_L g4076 ( 
.A(n_3977),
.B(n_3732),
.Y(n_4076)
);

OAI21x1_ASAP7_75t_L g4077 ( 
.A1(n_4005),
.A2(n_3663),
.B(n_3850),
.Y(n_4077)
);

OA21x2_ASAP7_75t_L g4078 ( 
.A1(n_3908),
.A2(n_3661),
.B(n_3830),
.Y(n_4078)
);

NOR2x1_ASAP7_75t_SL g4079 ( 
.A(n_3877),
.B(n_3779),
.Y(n_4079)
);

INVx3_ASAP7_75t_L g4080 ( 
.A(n_3932),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3866),
.Y(n_4081)
);

AOI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_3857),
.A2(n_3750),
.B(n_3780),
.Y(n_4082)
);

BUFx2_ASAP7_75t_L g4083 ( 
.A(n_3983),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3913),
.B(n_3730),
.Y(n_4084)
);

OAI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_4020),
.A2(n_3750),
.B1(n_3779),
.B2(n_3782),
.Y(n_4085)
);

NOR2x1_ASAP7_75t_R g4086 ( 
.A(n_3895),
.B(n_3772),
.Y(n_4086)
);

OAI21x1_ASAP7_75t_L g4087 ( 
.A1(n_3931),
.A2(n_3848),
.B(n_3753),
.Y(n_4087)
);

BUFx6f_ASAP7_75t_L g4088 ( 
.A(n_3902),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3867),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3873),
.Y(n_4090)
);

NOR2x1_ASAP7_75t_SL g4091 ( 
.A(n_3877),
.B(n_3730),
.Y(n_4091)
);

OAI21x1_ASAP7_75t_L g4092 ( 
.A1(n_4018),
.A2(n_3725),
.B(n_3730),
.Y(n_4092)
);

OAI21x1_ASAP7_75t_L g4093 ( 
.A1(n_3865),
.A2(n_3809),
.B(n_116),
.Y(n_4093)
);

OAI21x1_ASAP7_75t_L g4094 ( 
.A1(n_3935),
.A2(n_3809),
.B(n_117),
.Y(n_4094)
);

O2A1O1Ixp33_ASAP7_75t_SL g4095 ( 
.A1(n_3855),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_4095)
);

NAND2x1p5_ASAP7_75t_L g4096 ( 
.A(n_3919),
.B(n_119),
.Y(n_4096)
);

OA21x2_ASAP7_75t_L g4097 ( 
.A1(n_3875),
.A2(n_3890),
.B(n_3886),
.Y(n_4097)
);

INVx2_ASAP7_75t_SL g4098 ( 
.A(n_3899),
.Y(n_4098)
);

AOI21xp5_ASAP7_75t_L g4099 ( 
.A1(n_3871),
.A2(n_121),
.B(n_122),
.Y(n_4099)
);

OAI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_4020),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_4100)
);

OA21x2_ASAP7_75t_L g4101 ( 
.A1(n_3889),
.A2(n_124),
.B(n_125),
.Y(n_4101)
);

AO21x2_ASAP7_75t_L g4102 ( 
.A1(n_3891),
.A2(n_125),
.B(n_126),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_3919),
.A2(n_126),
.B(n_127),
.Y(n_4103)
);

O2A1O1Ixp5_ASAP7_75t_L g4104 ( 
.A1(n_3959),
.A2(n_130),
.B(n_127),
.C(n_128),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3911),
.A2(n_3888),
.B(n_3924),
.Y(n_4105)
);

BUFx3_ASAP7_75t_L g4106 ( 
.A(n_3861),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3862),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_L g4108 ( 
.A1(n_3934),
.A2(n_128),
.B(n_130),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3858),
.A2(n_132),
.B(n_134),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3939),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3986),
.Y(n_4111)
);

OA21x2_ASAP7_75t_L g4112 ( 
.A1(n_3956),
.A2(n_4006),
.B(n_3944),
.Y(n_4112)
);

AND2x4_ASAP7_75t_L g4113 ( 
.A(n_3874),
.B(n_136),
.Y(n_4113)
);

NAND2x1p5_ASAP7_75t_L g4114 ( 
.A(n_3919),
.B(n_137),
.Y(n_4114)
);

O2A1O1Ixp33_ASAP7_75t_L g4115 ( 
.A1(n_4010),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3876),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_3970),
.A2(n_142),
.B1(n_139),
.B2(n_141),
.Y(n_4117)
);

BUFx3_ASAP7_75t_L g4118 ( 
.A(n_3900),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_L g4119 ( 
.A(n_3928),
.B(n_142),
.Y(n_4119)
);

OR2x6_ASAP7_75t_L g4120 ( 
.A(n_3962),
.B(n_143),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_3978),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3940),
.B(n_143),
.Y(n_4122)
);

OAI21x1_ASAP7_75t_L g4123 ( 
.A1(n_3922),
.A2(n_144),
.B(n_145),
.Y(n_4123)
);

CKINVDCx6p67_ASAP7_75t_R g4124 ( 
.A(n_3989),
.Y(n_4124)
);

OAI21x1_ASAP7_75t_L g4125 ( 
.A1(n_3941),
.A2(n_144),
.B(n_145),
.Y(n_4125)
);

BUFx3_ASAP7_75t_L g4126 ( 
.A(n_3900),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3887),
.Y(n_4127)
);

OAI21x1_ASAP7_75t_L g4128 ( 
.A1(n_4033),
.A2(n_146),
.B(n_147),
.Y(n_4128)
);

OAI21x1_ASAP7_75t_L g4129 ( 
.A1(n_3974),
.A2(n_146),
.B(n_148),
.Y(n_4129)
);

OAI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_4026),
.A2(n_148),
.B(n_149),
.Y(n_4130)
);

OAI21x1_ASAP7_75t_L g4131 ( 
.A1(n_3918),
.A2(n_150),
.B(n_151),
.Y(n_4131)
);

AOI21x1_ASAP7_75t_L g4132 ( 
.A1(n_3958),
.A2(n_150),
.B(n_151),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_3998),
.Y(n_4133)
);

BUFx3_ASAP7_75t_L g4134 ( 
.A(n_3988),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3863),
.B(n_3893),
.Y(n_4135)
);

OAI21x1_ASAP7_75t_L g4136 ( 
.A1(n_3947),
.A2(n_152),
.B(n_153),
.Y(n_4136)
);

OAI21x1_ASAP7_75t_L g4137 ( 
.A1(n_3953),
.A2(n_4013),
.B(n_3885),
.Y(n_4137)
);

HB1xp67_ASAP7_75t_L g4138 ( 
.A(n_4031),
.Y(n_4138)
);

AOI22xp33_ASAP7_75t_SL g4139 ( 
.A1(n_4028),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4139)
);

NOR2xp67_ASAP7_75t_L g4140 ( 
.A(n_3943),
.B(n_154),
.Y(n_4140)
);

OAI21x1_ASAP7_75t_L g4141 ( 
.A1(n_3937),
.A2(n_155),
.B(n_156),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_3948),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3999),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3920),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3945),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3963),
.Y(n_4146)
);

OA21x2_ASAP7_75t_L g4147 ( 
.A1(n_3975),
.A2(n_157),
.B(n_158),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_3967),
.Y(n_4148)
);

AND2x4_ASAP7_75t_L g4149 ( 
.A(n_3881),
.B(n_157),
.Y(n_4149)
);

INVx2_ASAP7_75t_SL g4150 ( 
.A(n_3965),
.Y(n_4150)
);

BUFx3_ASAP7_75t_L g4151 ( 
.A(n_3995),
.Y(n_4151)
);

AOI22xp33_ASAP7_75t_L g4152 ( 
.A1(n_3952),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_4152)
);

NOR2xp67_ASAP7_75t_L g4153 ( 
.A(n_3943),
.B(n_159),
.Y(n_4153)
);

AO21x2_ASAP7_75t_L g4154 ( 
.A1(n_3984),
.A2(n_160),
.B(n_161),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3980),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3990),
.B(n_3993),
.Y(n_4156)
);

AOI21x1_ASAP7_75t_L g4157 ( 
.A1(n_4023),
.A2(n_161),
.B(n_162),
.Y(n_4157)
);

AOI22xp33_ASAP7_75t_L g4158 ( 
.A1(n_4007),
.A2(n_4017),
.B1(n_3962),
.B2(n_4012),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4000),
.Y(n_4159)
);

AO32x2_ASAP7_75t_L g4160 ( 
.A1(n_3896),
.A2(n_164),
.A3(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_4160)
);

OAI21x1_ASAP7_75t_L g4161 ( 
.A1(n_3949),
.A2(n_163),
.B(n_164),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4001),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3914),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3914),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_3864),
.A2(n_165),
.B(n_166),
.Y(n_4165)
);

CKINVDCx5p33_ASAP7_75t_R g4166 ( 
.A(n_3880),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3892),
.Y(n_4167)
);

OAI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_3991),
.A2(n_166),
.B(n_167),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3981),
.Y(n_4169)
);

OAI21x1_ASAP7_75t_L g4170 ( 
.A1(n_4014),
.A2(n_167),
.B(n_168),
.Y(n_4170)
);

NOR2xp33_ASAP7_75t_L g4171 ( 
.A(n_3884),
.B(n_168),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_3946),
.B(n_169),
.Y(n_4172)
);

OAI21x1_ASAP7_75t_L g4173 ( 
.A1(n_4024),
.A2(n_169),
.B(n_170),
.Y(n_4173)
);

BUFx2_ASAP7_75t_SL g4174 ( 
.A(n_3961),
.Y(n_4174)
);

BUFx4f_ASAP7_75t_SL g4175 ( 
.A(n_3982),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_3905),
.Y(n_4176)
);

NAND2x1p5_ASAP7_75t_L g4177 ( 
.A(n_3881),
.B(n_171),
.Y(n_4177)
);

NAND2x1p5_ASAP7_75t_L g4178 ( 
.A(n_3985),
.B(n_171),
.Y(n_4178)
);

AO31x2_ASAP7_75t_L g4179 ( 
.A1(n_3985),
.A2(n_174),
.A3(n_172),
.B(n_173),
.Y(n_4179)
);

NAND2x1p5_ASAP7_75t_L g4180 ( 
.A(n_3898),
.B(n_174),
.Y(n_4180)
);

OAI21x1_ASAP7_75t_L g4181 ( 
.A1(n_3923),
.A2(n_3957),
.B(n_4032),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_3869),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_4016),
.B(n_175),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3869),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3869),
.Y(n_4185)
);

OAI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_4030),
.A2(n_177),
.B(n_179),
.Y(n_4186)
);

OAI21x1_ASAP7_75t_SL g4187 ( 
.A1(n_3973),
.A2(n_180),
.B(n_181),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_4070),
.B(n_4004),
.Y(n_4188)
);

OAI21xp5_ASAP7_75t_L g4189 ( 
.A1(n_4099),
.A2(n_4027),
.B(n_4012),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4068),
.Y(n_4190)
);

CKINVDCx5p33_ASAP7_75t_R g4191 ( 
.A(n_4047),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4068),
.Y(n_4192)
);

AO21x2_ASAP7_75t_L g4193 ( 
.A1(n_4099),
.A2(n_3994),
.B(n_4011),
.Y(n_4193)
);

OR2x2_ASAP7_75t_L g4194 ( 
.A(n_4060),
.B(n_4015),
.Y(n_4194)
);

AOI22xp33_ASAP7_75t_L g4195 ( 
.A1(n_4109),
.A2(n_3882),
.B1(n_4027),
.B2(n_3992),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_4079),
.B(n_4091),
.Y(n_4196)
);

BUFx3_ASAP7_75t_L g4197 ( 
.A(n_4088),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4097),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_4112),
.Y(n_4199)
);

INVx6_ASAP7_75t_L g4200 ( 
.A(n_4088),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4097),
.Y(n_4201)
);

INVx1_ASAP7_75t_SL g4202 ( 
.A(n_4112),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4156),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4137),
.Y(n_4204)
);

AOI22xp33_ASAP7_75t_L g4205 ( 
.A1(n_4109),
.A2(n_3915),
.B1(n_4019),
.B2(n_3961),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_4088),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_4078),
.B(n_4040),
.Y(n_4207)
);

OAI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_4034),
.A2(n_4009),
.B1(n_4021),
.B2(n_4011),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4156),
.Y(n_4209)
);

BUFx3_ASAP7_75t_L g4210 ( 
.A(n_4044),
.Y(n_4210)
);

OA21x2_ASAP7_75t_L g4211 ( 
.A1(n_4105),
.A2(n_4074),
.B(n_4181),
.Y(n_4211)
);

OAI22xp33_ASAP7_75t_L g4212 ( 
.A1(n_4051),
.A2(n_3897),
.B1(n_3996),
.B2(n_3954),
.Y(n_4212)
);

AOI22xp33_ASAP7_75t_L g4213 ( 
.A1(n_4168),
.A2(n_3903),
.B1(n_3968),
.B2(n_4022),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4070),
.B(n_3903),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_4081),
.Y(n_4215)
);

NAND2x1p5_ASAP7_75t_L g4216 ( 
.A(n_4078),
.B(n_3968),
.Y(n_4216)
);

BUFx2_ASAP7_75t_SL g4217 ( 
.A(n_4118),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4050),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4138),
.Y(n_4219)
);

INVx4_ASAP7_75t_L g4220 ( 
.A(n_4055),
.Y(n_4220)
);

INVx4_ASAP7_75t_L g4221 ( 
.A(n_4055),
.Y(n_4221)
);

AOI22xp33_ASAP7_75t_SL g4222 ( 
.A1(n_4066),
.A2(n_4021),
.B1(n_4009),
.B2(n_3969),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_4071),
.B(n_3954),
.Y(n_4223)
);

AOI22xp33_ASAP7_75t_SL g4224 ( 
.A1(n_4066),
.A2(n_4021),
.B1(n_3996),
.B2(n_3997),
.Y(n_4224)
);

INVx2_ASAP7_75t_SL g4225 ( 
.A(n_4175),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4052),
.Y(n_4226)
);

INVx3_ASAP7_75t_L g4227 ( 
.A(n_4080),
.Y(n_4227)
);

CKINVDCx20_ASAP7_75t_R g4228 ( 
.A(n_4124),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4061),
.Y(n_4229)
);

AOI21x1_ASAP7_75t_L g4230 ( 
.A1(n_4122),
.A2(n_3996),
.B(n_3954),
.Y(n_4230)
);

AOI21x1_ASAP7_75t_L g4231 ( 
.A1(n_4122),
.A2(n_4008),
.B(n_3997),
.Y(n_4231)
);

INVxp67_ASAP7_75t_L g4232 ( 
.A(n_4101),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_4090),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_4163),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4089),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4110),
.Y(n_4236)
);

INVx2_ASAP7_75t_SL g4237 ( 
.A(n_4142),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4135),
.B(n_3997),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4145),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4164),
.Y(n_4240)
);

INVx1_ASAP7_75t_SL g4241 ( 
.A(n_4174),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4146),
.Y(n_4242)
);

AOI22xp33_ASAP7_75t_SL g4243 ( 
.A1(n_4168),
.A2(n_4008),
.B1(n_182),
.B2(n_180),
.Y(n_4243)
);

INVx3_ASAP7_75t_L g4244 ( 
.A(n_4080),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_4159),
.Y(n_4245)
);

AND2x4_ASAP7_75t_L g4246 ( 
.A(n_4076),
.B(n_4008),
.Y(n_4246)
);

INVx2_ASAP7_75t_L g4247 ( 
.A(n_4162),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4116),
.Y(n_4248)
);

INVx3_ASAP7_75t_L g4249 ( 
.A(n_4059),
.Y(n_4249)
);

AOI22xp33_ASAP7_75t_SL g4250 ( 
.A1(n_4186),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_4111),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_4133),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_4143),
.Y(n_4253)
);

INVx6_ASAP7_75t_L g4254 ( 
.A(n_4059),
.Y(n_4254)
);

INVx1_ASAP7_75t_SL g4255 ( 
.A(n_4101),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4107),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_4075),
.B(n_4083),
.Y(n_4257)
);

OR2x6_ASAP7_75t_L g4258 ( 
.A(n_4096),
.B(n_183),
.Y(n_4258)
);

BUFx2_ASAP7_75t_R g4259 ( 
.A(n_4126),
.Y(n_4259)
);

AND2x4_ASAP7_75t_L g4260 ( 
.A(n_4076),
.B(n_184),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4127),
.Y(n_4261)
);

OAI22xp33_ASAP7_75t_L g4262 ( 
.A1(n_4051),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_4262)
);

AOI22xp33_ASAP7_75t_SL g4263 ( 
.A1(n_4186),
.A2(n_4100),
.B1(n_4120),
.B2(n_4057),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4040),
.B(n_186),
.Y(n_4264)
);

BUFx2_ASAP7_75t_R g4265 ( 
.A(n_4049),
.Y(n_4265)
);

HB1xp67_ASAP7_75t_L g4266 ( 
.A(n_4038),
.Y(n_4266)
);

AOI22xp33_ASAP7_75t_SL g4267 ( 
.A1(n_4100),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_4267)
);

OAI21x1_ASAP7_75t_L g4268 ( 
.A1(n_4035),
.A2(n_188),
.B(n_189),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4144),
.Y(n_4269)
);

AOI21x1_ASAP7_75t_L g4270 ( 
.A1(n_4140),
.A2(n_190),
.B(n_191),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4169),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4060),
.B(n_192),
.Y(n_4272)
);

AOI22xp33_ASAP7_75t_L g4273 ( 
.A1(n_4165),
.A2(n_651),
.B1(n_196),
.B2(n_194),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4148),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4155),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4084),
.Y(n_4276)
);

BUFx10_ASAP7_75t_L g4277 ( 
.A(n_4059),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4184),
.Y(n_4278)
);

HB1xp67_ASAP7_75t_L g4279 ( 
.A(n_4038),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4084),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4102),
.B(n_195),
.Y(n_4281)
);

BUFx2_ASAP7_75t_L g4282 ( 
.A(n_4065),
.Y(n_4282)
);

BUFx12f_ASAP7_75t_L g4283 ( 
.A(n_4121),
.Y(n_4283)
);

CKINVDCx20_ASAP7_75t_R g4284 ( 
.A(n_4069),
.Y(n_4284)
);

OAI21x1_ASAP7_75t_L g4285 ( 
.A1(n_4037),
.A2(n_195),
.B(n_196),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4185),
.Y(n_4286)
);

OA21x2_ASAP7_75t_L g4287 ( 
.A1(n_4087),
.A2(n_197),
.B(n_198),
.Y(n_4287)
);

CKINVDCx20_ASAP7_75t_R g4288 ( 
.A(n_4151),
.Y(n_4288)
);

OAI21x1_ASAP7_75t_L g4289 ( 
.A1(n_4042),
.A2(n_199),
.B(n_200),
.Y(n_4289)
);

AO21x2_ASAP7_75t_L g4290 ( 
.A1(n_4103),
.A2(n_199),
.B(n_201),
.Y(n_4290)
);

NAND2x1p5_ASAP7_75t_L g4291 ( 
.A(n_4043),
.B(n_201),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4167),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4065),
.B(n_202),
.Y(n_4293)
);

AOI22xp33_ASAP7_75t_L g4294 ( 
.A1(n_4165),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4147),
.Y(n_4295)
);

AOI21x1_ASAP7_75t_L g4296 ( 
.A1(n_4140),
.A2(n_204),
.B(n_205),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4147),
.Y(n_4297)
);

INVxp67_ASAP7_75t_L g4298 ( 
.A(n_4102),
.Y(n_4298)
);

INVx6_ASAP7_75t_L g4299 ( 
.A(n_4039),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4176),
.Y(n_4300)
);

AOI22xp33_ASAP7_75t_L g4301 ( 
.A1(n_4130),
.A2(n_4119),
.B1(n_4057),
.B2(n_4171),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4154),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4098),
.B(n_206),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4182),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_4096),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4182),
.Y(n_4306)
);

OAI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_4103),
.A2(n_206),
.B(n_207),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4154),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4179),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4182),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4179),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4179),
.Y(n_4312)
);

BUFx6f_ASAP7_75t_L g4313 ( 
.A(n_4178),
.Y(n_4313)
);

NAND2x1p5_ASAP7_75t_L g4314 ( 
.A(n_4045),
.B(n_208),
.Y(n_4314)
);

AOI22xp33_ASAP7_75t_L g4315 ( 
.A1(n_4130),
.A2(n_651),
.B1(n_210),
.B2(n_208),
.Y(n_4315)
);

OA21x2_ASAP7_75t_L g4316 ( 
.A1(n_4077),
.A2(n_209),
.B(n_211),
.Y(n_4316)
);

OAI21x1_ASAP7_75t_L g4317 ( 
.A1(n_4073),
.A2(n_211),
.B(n_212),
.Y(n_4317)
);

BUFx8_ASAP7_75t_SL g4318 ( 
.A(n_4134),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4063),
.Y(n_4319)
);

AO21x2_ASAP7_75t_L g4320 ( 
.A1(n_4153),
.A2(n_212),
.B(n_213),
.Y(n_4320)
);

AOI22xp33_ASAP7_75t_SL g4321 ( 
.A1(n_4120),
.A2(n_216),
.B1(n_213),
.B2(n_215),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_4166),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4063),
.Y(n_4323)
);

AOI21x1_ASAP7_75t_L g4324 ( 
.A1(n_4153),
.A2(n_215),
.B(n_217),
.Y(n_4324)
);

HB1xp67_ASAP7_75t_L g4325 ( 
.A(n_4062),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4036),
.Y(n_4326)
);

AOI222xp33_ASAP7_75t_L g4327 ( 
.A1(n_4086),
.A2(n_4152),
.B1(n_4158),
.B2(n_4117),
.C1(n_4183),
.C2(n_4072),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4092),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4036),
.Y(n_4329)
);

AOI22xp33_ASAP7_75t_L g4330 ( 
.A1(n_4058),
.A2(n_220),
.B1(n_217),
.B2(n_218),
.Y(n_4330)
);

OAI22xp33_ASAP7_75t_L g4331 ( 
.A1(n_4120),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_4331)
);

INVx3_ASAP7_75t_L g4332 ( 
.A(n_4106),
.Y(n_4332)
);

AO21x2_ASAP7_75t_L g4333 ( 
.A1(n_4157),
.A2(n_222),
.B(n_223),
.Y(n_4333)
);

CKINVDCx20_ASAP7_75t_R g4334 ( 
.A(n_4039),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4062),
.B(n_223),
.Y(n_4335)
);

HB1xp67_ASAP7_75t_L g4336 ( 
.A(n_4128),
.Y(n_4336)
);

INVx2_ASAP7_75t_SL g4337 ( 
.A(n_4150),
.Y(n_4337)
);

AOI21x1_ASAP7_75t_L g4338 ( 
.A1(n_4132),
.A2(n_224),
.B(n_225),
.Y(n_4338)
);

AND2x4_ASAP7_75t_L g4339 ( 
.A(n_4113),
.B(n_224),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4160),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4160),
.Y(n_4341)
);

BUFx2_ASAP7_75t_L g4342 ( 
.A(n_4113),
.Y(n_4342)
);

INVx2_ASAP7_75t_SL g4343 ( 
.A(n_4149),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4094),
.Y(n_4344)
);

AOI21x1_ASAP7_75t_L g4345 ( 
.A1(n_4082),
.A2(n_225),
.B(n_226),
.Y(n_4345)
);

AOI22xp5_ASAP7_75t_SL g4346 ( 
.A1(n_4180),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_4346)
);

BUFx8_ASAP7_75t_L g4347 ( 
.A(n_4149),
.Y(n_4347)
);

INVx1_ASAP7_75t_SL g4348 ( 
.A(n_4178),
.Y(n_4348)
);

BUFx3_ASAP7_75t_L g4349 ( 
.A(n_4172),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4160),
.Y(n_4350)
);

BUFx2_ASAP7_75t_L g4351 ( 
.A(n_4114),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4125),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4352),
.B(n_4082),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4198),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4190),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4192),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4201),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_4216),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4216),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4239),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_4230),
.Y(n_4361)
);

OAI21x1_ASAP7_75t_L g4362 ( 
.A1(n_4295),
.A2(n_4054),
.B(n_4123),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4214),
.B(n_4093),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4242),
.Y(n_4364)
);

HB1xp67_ASAP7_75t_L g4365 ( 
.A(n_4199),
.Y(n_4365)
);

OAI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_4263),
.A2(n_4104),
.B(n_4115),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4218),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_4231),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4226),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_4265),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4245),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4229),
.Y(n_4372)
);

OR2x2_ASAP7_75t_L g4373 ( 
.A(n_4207),
.B(n_4183),
.Y(n_4373)
);

INVx4_ASAP7_75t_L g4374 ( 
.A(n_4200),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_4241),
.B(n_4048),
.Y(n_4375)
);

AND2x4_ASAP7_75t_L g4376 ( 
.A(n_4196),
.B(n_4048),
.Y(n_4376)
);

INVx3_ASAP7_75t_L g4377 ( 
.A(n_4277),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4247),
.Y(n_4378)
);

OAI21x1_ASAP7_75t_L g4379 ( 
.A1(n_4297),
.A2(n_4053),
.B(n_4141),
.Y(n_4379)
);

INVxp67_ASAP7_75t_SL g4380 ( 
.A(n_4232),
.Y(n_4380)
);

BUFx3_ASAP7_75t_L g4381 ( 
.A(n_4299),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4235),
.Y(n_4382)
);

AO21x2_ASAP7_75t_L g4383 ( 
.A1(n_4266),
.A2(n_4095),
.B(n_4187),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4278),
.Y(n_4384)
);

INVx3_ASAP7_75t_L g4385 ( 
.A(n_4277),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4236),
.Y(n_4386)
);

INVxp67_ASAP7_75t_L g4387 ( 
.A(n_4336),
.Y(n_4387)
);

AOI22xp33_ASAP7_75t_L g4388 ( 
.A1(n_4263),
.A2(n_4139),
.B1(n_4108),
.B2(n_4129),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4248),
.Y(n_4389)
);

AO21x2_ASAP7_75t_L g4390 ( 
.A1(n_4279),
.A2(n_4085),
.B(n_4131),
.Y(n_4390)
);

BUFx6f_ASAP7_75t_L g4391 ( 
.A(n_4200),
.Y(n_4391)
);

INVx2_ASAP7_75t_SL g4392 ( 
.A(n_4299),
.Y(n_4392)
);

INVx3_ASAP7_75t_SL g4393 ( 
.A(n_4258),
.Y(n_4393)
);

INVx2_ASAP7_75t_L g4394 ( 
.A(n_4316),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4316),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4261),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4269),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4271),
.Y(n_4398)
);

INVx2_ASAP7_75t_SL g4399 ( 
.A(n_4197),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_4215),
.Y(n_4400)
);

OA21x2_ASAP7_75t_L g4401 ( 
.A1(n_4232),
.A2(n_4161),
.B(n_4136),
.Y(n_4401)
);

INVx2_ASAP7_75t_L g4402 ( 
.A(n_4233),
.Y(n_4402)
);

INVxp67_ASAP7_75t_SL g4403 ( 
.A(n_4298),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4241),
.B(n_4177),
.Y(n_4404)
);

OR2x2_ASAP7_75t_L g4405 ( 
.A(n_4207),
.B(n_4072),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4203),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4202),
.Y(n_4407)
);

INVx2_ASAP7_75t_SL g4408 ( 
.A(n_4206),
.Y(n_4408)
);

BUFx2_ASAP7_75t_L g4409 ( 
.A(n_4196),
.Y(n_4409)
);

BUFx2_ASAP7_75t_L g4410 ( 
.A(n_4282),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4209),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4222),
.B(n_4046),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4309),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4319),
.B(n_4064),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4202),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4311),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4276),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4280),
.Y(n_4418)
);

BUFx3_ASAP7_75t_L g4419 ( 
.A(n_4334),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_4251),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4312),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4252),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4253),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4335),
.Y(n_4424)
);

BUFx3_ASAP7_75t_L g4425 ( 
.A(n_4318),
.Y(n_4425)
);

OAI21x1_ASAP7_75t_L g4426 ( 
.A1(n_4204),
.A2(n_4308),
.B(n_4302),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4335),
.Y(n_4427)
);

NOR2xp67_ASAP7_75t_SL g4428 ( 
.A(n_4217),
.B(n_4086),
.Y(n_4428)
);

HB1xp67_ASAP7_75t_L g4429 ( 
.A(n_4255),
.Y(n_4429)
);

OR2x2_ASAP7_75t_L g4430 ( 
.A(n_4194),
.B(n_4219),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4256),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4275),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4274),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_4193),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_4193),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4287),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4344),
.Y(n_4437)
);

AOI21xp33_ASAP7_75t_L g4438 ( 
.A1(n_4327),
.A2(n_4224),
.B(n_4255),
.Y(n_4438)
);

OAI21x1_ASAP7_75t_L g4439 ( 
.A1(n_4328),
.A2(n_4173),
.B(n_4170),
.Y(n_4439)
);

INVx3_ASAP7_75t_L g4440 ( 
.A(n_4254),
.Y(n_4440)
);

INVxp67_ASAP7_75t_L g4441 ( 
.A(n_4259),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4287),
.Y(n_4442)
);

HB1xp67_ASAP7_75t_L g4443 ( 
.A(n_4325),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_4254),
.Y(n_4444)
);

OAI21x1_ASAP7_75t_L g4445 ( 
.A1(n_4211),
.A2(n_4180),
.B(n_4046),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4286),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4298),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_4227),
.A2(n_4244),
.B(n_4211),
.Y(n_4448)
);

INVx2_ASAP7_75t_L g4449 ( 
.A(n_4234),
.Y(n_4449)
);

INVx3_ASAP7_75t_L g4450 ( 
.A(n_4305),
.Y(n_4450)
);

A2O1A1Ixp33_ASAP7_75t_L g4451 ( 
.A1(n_4189),
.A2(n_4115),
.B(n_4056),
.C(n_4041),
.Y(n_4451)
);

AO21x2_ASAP7_75t_L g4452 ( 
.A1(n_4281),
.A2(n_4067),
.B(n_4056),
.Y(n_4452)
);

AO21x1_ASAP7_75t_L g4453 ( 
.A1(n_4340),
.A2(n_227),
.B(n_228),
.Y(n_4453)
);

BUFx6f_ASAP7_75t_L g4454 ( 
.A(n_4220),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4281),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4240),
.Y(n_4456)
);

BUFx2_ASAP7_75t_L g4457 ( 
.A(n_4305),
.Y(n_4457)
);

OA21x2_ASAP7_75t_L g4458 ( 
.A1(n_4341),
.A2(n_229),
.B(n_231),
.Y(n_4458)
);

BUFx2_ASAP7_75t_L g4459 ( 
.A(n_4305),
.Y(n_4459)
);

INVx2_ASAP7_75t_SL g4460 ( 
.A(n_4249),
.Y(n_4460)
);

OAI21x1_ASAP7_75t_L g4461 ( 
.A1(n_4227),
.A2(n_229),
.B(n_232),
.Y(n_4461)
);

INVx4_ASAP7_75t_L g4462 ( 
.A(n_4220),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4350),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_4323),
.B(n_232),
.Y(n_4464)
);

HB1xp67_ASAP7_75t_L g4465 ( 
.A(n_4333),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4300),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4292),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4317),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4264),
.Y(n_4469)
);

INVx1_ASAP7_75t_SL g4470 ( 
.A(n_4259),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4264),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_4313),
.Y(n_4472)
);

INVx3_ASAP7_75t_L g4473 ( 
.A(n_4221),
.Y(n_4473)
);

CKINVDCx10_ASAP7_75t_R g4474 ( 
.A(n_4258),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4342),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4304),
.Y(n_4476)
);

INVx3_ASAP7_75t_L g4477 ( 
.A(n_4221),
.Y(n_4477)
);

OAI21x1_ASAP7_75t_L g4478 ( 
.A1(n_4244),
.A2(n_234),
.B(n_235),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4313),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4306),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4310),
.Y(n_4481)
);

OR2x6_ASAP7_75t_L g4482 ( 
.A(n_4314),
.B(n_234),
.Y(n_4482)
);

NOR2x1_ASAP7_75t_SL g4483 ( 
.A(n_4313),
.B(n_237),
.Y(n_4483)
);

CKINVDCx20_ASAP7_75t_R g4484 ( 
.A(n_4284),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4272),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4320),
.Y(n_4486)
);

OR2x2_ASAP7_75t_L g4487 ( 
.A(n_4237),
.B(n_238),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4326),
.B(n_4329),
.Y(n_4488)
);

CKINVDCx5p33_ASAP7_75t_R g4489 ( 
.A(n_4265),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4272),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4268),
.Y(n_4491)
);

AND2x4_ASAP7_75t_SL g4492 ( 
.A(n_4249),
.B(n_238),
.Y(n_4492)
);

AOI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_4224),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4246),
.B(n_240),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4257),
.Y(n_4495)
);

AND2x4_ASAP7_75t_L g4496 ( 
.A(n_4246),
.B(n_241),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4188),
.B(n_242),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4208),
.Y(n_4498)
);

NOR2xp33_ASAP7_75t_L g4499 ( 
.A(n_4332),
.B(n_243),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4208),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4333),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_4320),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4314),
.Y(n_4503)
);

BUFx3_ASAP7_75t_L g4504 ( 
.A(n_4322),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4270),
.Y(n_4505)
);

INVx1_ASAP7_75t_SL g4506 ( 
.A(n_4228),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4285),
.Y(n_4507)
);

BUFx2_ASAP7_75t_L g4508 ( 
.A(n_4189),
.Y(n_4508)
);

HB1xp67_ASAP7_75t_L g4509 ( 
.A(n_4290),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4345),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4409),
.B(n_4332),
.Y(n_4511)
);

AOI221xp5_ASAP7_75t_L g4512 ( 
.A1(n_4438),
.A2(n_4262),
.B1(n_4301),
.B2(n_4331),
.C(n_4222),
.Y(n_4512)
);

BUFx2_ASAP7_75t_L g4513 ( 
.A(n_4504),
.Y(n_4513)
);

AOI22xp33_ASAP7_75t_L g4514 ( 
.A1(n_4508),
.A2(n_4412),
.B1(n_4366),
.B2(n_4498),
.Y(n_4514)
);

AOI22xp33_ASAP7_75t_L g4515 ( 
.A1(n_4500),
.A2(n_4327),
.B1(n_4243),
.B2(n_4250),
.Y(n_4515)
);

NOR2x1_ASAP7_75t_SL g4516 ( 
.A(n_4452),
.B(n_4258),
.Y(n_4516)
);

AOI22xp33_ASAP7_75t_L g4517 ( 
.A1(n_4376),
.A2(n_4243),
.B1(n_4250),
.B2(n_4195),
.Y(n_4517)
);

AOI22xp33_ASAP7_75t_L g4518 ( 
.A1(n_4376),
.A2(n_4307),
.B1(n_4205),
.B2(n_4290),
.Y(n_4518)
);

HB1xp67_ASAP7_75t_L g4519 ( 
.A(n_4429),
.Y(n_4519)
);

OR2x2_ASAP7_75t_L g4520 ( 
.A(n_4430),
.B(n_4348),
.Y(n_4520)
);

AOI21xp5_ASAP7_75t_L g4521 ( 
.A1(n_4451),
.A2(n_4307),
.B(n_4346),
.Y(n_4521)
);

OAI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_4451),
.A2(n_4388),
.B1(n_4493),
.B2(n_4393),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_4441),
.A2(n_4346),
.B(n_4191),
.Y(n_4523)
);

NOR2x1_ASAP7_75t_R g4524 ( 
.A(n_4370),
.B(n_4283),
.Y(n_4524)
);

INVx3_ASAP7_75t_L g4525 ( 
.A(n_4381),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4504),
.B(n_4351),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_SL g4527 ( 
.A1(n_4483),
.A2(n_4291),
.B(n_4339),
.Y(n_4527)
);

AOI22xp33_ASAP7_75t_SL g4528 ( 
.A1(n_4509),
.A2(n_4348),
.B1(n_4347),
.B2(n_4291),
.Y(n_4528)
);

AOI22x1_ASAP7_75t_L g4529 ( 
.A1(n_4370),
.A2(n_4225),
.B1(n_4260),
.B2(n_4339),
.Y(n_4529)
);

A2O1A1Ixp33_ASAP7_75t_L g4530 ( 
.A1(n_4441),
.A2(n_4388),
.B(n_4445),
.C(n_4489),
.Y(n_4530)
);

OAI33xp33_ASAP7_75t_L g4531 ( 
.A1(n_4463),
.A2(n_4212),
.A3(n_4321),
.B1(n_4267),
.B2(n_4338),
.B3(n_4315),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4429),
.Y(n_4532)
);

OAI21x1_ASAP7_75t_L g4533 ( 
.A1(n_4448),
.A2(n_4324),
.B(n_4296),
.Y(n_4533)
);

OAI221xp5_ASAP7_75t_L g4534 ( 
.A1(n_4509),
.A2(n_4321),
.B1(n_4213),
.B2(n_4267),
.C(n_4294),
.Y(n_4534)
);

INVx4_ASAP7_75t_L g4535 ( 
.A(n_4425),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4413),
.Y(n_4536)
);

OAI22xp5_ASAP7_75t_L g4537 ( 
.A1(n_4393),
.A2(n_4273),
.B1(n_4343),
.B2(n_4337),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4416),
.Y(n_4538)
);

AND2x4_ASAP7_75t_L g4539 ( 
.A(n_4377),
.B(n_4260),
.Y(n_4539)
);

BUFx6f_ASAP7_75t_L g4540 ( 
.A(n_4425),
.Y(n_4540)
);

AOI33xp33_ASAP7_75t_L g4541 ( 
.A1(n_4455),
.A2(n_4330),
.A3(n_4303),
.B1(n_4293),
.B2(n_4238),
.B3(n_4347),
.Y(n_4541)
);

CKINVDCx5p33_ASAP7_75t_R g4542 ( 
.A(n_4489),
.Y(n_4542)
);

AOI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_4376),
.A2(n_4349),
.B1(n_4223),
.B2(n_4210),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4470),
.A2(n_4288),
.B1(n_4289),
.B2(n_245),
.Y(n_4544)
);

AOI222xp33_ASAP7_75t_L g4545 ( 
.A1(n_4428),
.A2(n_246),
.B1(n_249),
.B2(n_243),
.C1(n_244),
.C2(n_248),
.Y(n_4545)
);

OAI22xp5_ASAP7_75t_L g4546 ( 
.A1(n_4465),
.A2(n_249),
.B1(n_244),
.B2(n_248),
.Y(n_4546)
);

AOI322xp5_ASAP7_75t_L g4547 ( 
.A1(n_4465),
.A2(n_255),
.A3(n_254),
.B1(n_252),
.B2(n_250),
.C1(n_251),
.C2(n_253),
.Y(n_4547)
);

A2O1A1Ixp33_ASAP7_75t_L g4548 ( 
.A1(n_4445),
.A2(n_254),
.B(n_250),
.C(n_253),
.Y(n_4548)
);

BUFx12f_ASAP7_75t_L g4549 ( 
.A(n_4392),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4440),
.B(n_4444),
.Y(n_4550)
);

OAI22xp33_ASAP7_75t_L g4551 ( 
.A1(n_4410),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_4551)
);

OAI21x1_ASAP7_75t_L g4552 ( 
.A1(n_4426),
.A2(n_257),
.B(n_259),
.Y(n_4552)
);

AOI221xp5_ASAP7_75t_L g4553 ( 
.A1(n_4380),
.A2(n_263),
.B1(n_259),
.B2(n_260),
.C(n_264),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4440),
.B(n_263),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4444),
.B(n_265),
.Y(n_4555)
);

NAND3xp33_ASAP7_75t_L g4556 ( 
.A(n_4380),
.B(n_4501),
.C(n_4510),
.Y(n_4556)
);

AOI22xp33_ASAP7_75t_L g4557 ( 
.A1(n_4363),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_4557)
);

AOI22xp33_ASAP7_75t_SL g4558 ( 
.A1(n_4452),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_4375),
.B(n_4457),
.Y(n_4559)
);

AOI21xp33_ASAP7_75t_L g4560 ( 
.A1(n_4405),
.A2(n_269),
.B(n_270),
.Y(n_4560)
);

INVx3_ASAP7_75t_L g4561 ( 
.A(n_4381),
.Y(n_4561)
);

OR2x2_ASAP7_75t_L g4562 ( 
.A(n_4373),
.B(n_269),
.Y(n_4562)
);

AOI22xp33_ASAP7_75t_L g4563 ( 
.A1(n_4424),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_4563)
);

OAI22xp5_ASAP7_75t_L g4564 ( 
.A1(n_4495),
.A2(n_4482),
.B1(n_4385),
.B2(n_4377),
.Y(n_4564)
);

AOI22xp33_ASAP7_75t_L g4565 ( 
.A1(n_4427),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_4565)
);

AOI22xp33_ASAP7_75t_L g4566 ( 
.A1(n_4475),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_4566)
);

AOI22xp5_ASAP7_75t_L g4567 ( 
.A1(n_4374),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.Y(n_4567)
);

AOI22xp33_ASAP7_75t_SL g4568 ( 
.A1(n_4383),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_4568)
);

A2O1A1Ixp33_ASAP7_75t_L g4569 ( 
.A1(n_4486),
.A2(n_283),
.B(n_279),
.C(n_282),
.Y(n_4569)
);

AO21x2_ASAP7_75t_L g4570 ( 
.A1(n_4403),
.A2(n_282),
.B(n_283),
.Y(n_4570)
);

OAI221xp5_ASAP7_75t_L g4571 ( 
.A1(n_4353),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.C(n_287),
.Y(n_4571)
);

INVxp67_ASAP7_75t_SL g4572 ( 
.A(n_4391),
.Y(n_4572)
);

O2A1O1Ixp33_ASAP7_75t_L g4573 ( 
.A1(n_4486),
.A2(n_4502),
.B(n_4482),
.C(n_4453),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4485),
.B(n_287),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4421),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4459),
.B(n_288),
.Y(n_4576)
);

OAI221xp5_ASAP7_75t_L g4577 ( 
.A1(n_4502),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4360),
.Y(n_4578)
);

AOI222xp33_ASAP7_75t_L g4579 ( 
.A1(n_4490),
.A2(n_291),
.B1(n_293),
.B2(n_289),
.C1(n_290),
.C2(n_292),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4482),
.A2(n_297),
.B1(n_292),
.B2(n_294),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4404),
.B(n_294),
.Y(n_4581)
);

OAI22xp5_ASAP7_75t_L g4582 ( 
.A1(n_4385),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_4582)
);

AOI22xp33_ASAP7_75t_L g4583 ( 
.A1(n_4414),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4364),
.Y(n_4584)
);

AOI22xp33_ASAP7_75t_L g4585 ( 
.A1(n_4390),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4367),
.Y(n_4586)
);

BUFx2_ASAP7_75t_L g4587 ( 
.A(n_4374),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4369),
.Y(n_4588)
);

AOI22xp33_ASAP7_75t_L g4589 ( 
.A1(n_4390),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_4589)
);

AOI22xp33_ASAP7_75t_L g4590 ( 
.A1(n_4454),
.A2(n_306),
.B1(n_303),
.B2(n_304),
.Y(n_4590)
);

AOI221xp5_ASAP7_75t_L g4591 ( 
.A1(n_4436),
.A2(n_308),
.B1(n_304),
.B2(n_307),
.C(n_309),
.Y(n_4591)
);

OAI22xp5_ASAP7_75t_L g4592 ( 
.A1(n_4458),
.A2(n_310),
.B1(n_307),
.B2(n_308),
.Y(n_4592)
);

INVxp67_ASAP7_75t_SL g4593 ( 
.A(n_4391),
.Y(n_4593)
);

HB1xp67_ASAP7_75t_L g4594 ( 
.A(n_4365),
.Y(n_4594)
);

AOI22xp33_ASAP7_75t_L g4595 ( 
.A1(n_4454),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_4595)
);

OAI21x1_ASAP7_75t_L g4596 ( 
.A1(n_4426),
.A2(n_312),
.B(n_313),
.Y(n_4596)
);

OAI221xp5_ASAP7_75t_L g4597 ( 
.A1(n_4473),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.C(n_316),
.Y(n_4597)
);

BUFx6f_ASAP7_75t_L g4598 ( 
.A(n_4419),
.Y(n_4598)
);

AOI22xp33_ASAP7_75t_L g4599 ( 
.A1(n_4454),
.A2(n_317),
.B1(n_314),
.B2(n_316),
.Y(n_4599)
);

BUFx6f_ASAP7_75t_L g4600 ( 
.A(n_4419),
.Y(n_4600)
);

AOI222xp33_ASAP7_75t_L g4601 ( 
.A1(n_4469),
.A2(n_320),
.B1(n_322),
.B2(n_318),
.C1(n_319),
.C2(n_321),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4391),
.Y(n_4602)
);

OAI211xp5_ASAP7_75t_L g4603 ( 
.A1(n_4434),
.A2(n_322),
.B(n_318),
.C(n_320),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4488),
.B(n_323),
.Y(n_4604)
);

CKINVDCx5p33_ASAP7_75t_R g4605 ( 
.A(n_4484),
.Y(n_4605)
);

AOI21xp33_ASAP7_75t_L g4606 ( 
.A1(n_4442),
.A2(n_324),
.B(n_325),
.Y(n_4606)
);

OAI211xp5_ASAP7_75t_L g4607 ( 
.A1(n_4434),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_4607)
);

BUFx4f_ASAP7_75t_SL g4608 ( 
.A(n_4484),
.Y(n_4608)
);

AOI221xp5_ASAP7_75t_L g4609 ( 
.A1(n_4387),
.A2(n_4435),
.B1(n_4395),
.B2(n_4394),
.C(n_4403),
.Y(n_4609)
);

AOI21xp5_ASAP7_75t_L g4610 ( 
.A1(n_4383),
.A2(n_326),
.B(n_327),
.Y(n_4610)
);

AOI22xp33_ASAP7_75t_L g4611 ( 
.A1(n_4454),
.A2(n_331),
.B1(n_328),
.B2(n_329),
.Y(n_4611)
);

BUFx3_ASAP7_75t_L g4612 ( 
.A(n_4391),
.Y(n_4612)
);

AOI22xp33_ASAP7_75t_L g4613 ( 
.A1(n_4471),
.A2(n_331),
.B1(n_328),
.B2(n_329),
.Y(n_4613)
);

AOI22xp33_ASAP7_75t_L g4614 ( 
.A1(n_4468),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_4614)
);

A2O1A1Ixp33_ASAP7_75t_L g4615 ( 
.A1(n_4435),
.A2(n_336),
.B(n_333),
.C(n_335),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4460),
.B(n_336),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4450),
.B(n_338),
.Y(n_4617)
);

AOI22xp33_ASAP7_75t_L g4618 ( 
.A1(n_4468),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4450),
.B(n_339),
.Y(n_4619)
);

INVx4_ASAP7_75t_L g4620 ( 
.A(n_4496),
.Y(n_4620)
);

AO21x2_ASAP7_75t_L g4621 ( 
.A1(n_4365),
.A2(n_340),
.B(n_341),
.Y(n_4621)
);

AOI222xp33_ASAP7_75t_L g4622 ( 
.A1(n_4499),
.A2(n_341),
.B1(n_342),
.B2(n_344),
.C1(n_345),
.C2(n_346),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4372),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4472),
.B(n_342),
.Y(n_4624)
);

OAI22xp33_ASAP7_75t_L g4625 ( 
.A1(n_4458),
.A2(n_347),
.B1(n_344),
.B2(n_345),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4503),
.B(n_347),
.Y(n_4626)
);

AOI22xp33_ASAP7_75t_L g4627 ( 
.A1(n_4491),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_4627)
);

AOI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4507),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4473),
.Y(n_4629)
);

CKINVDCx5p33_ASAP7_75t_R g4630 ( 
.A(n_4474),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4477),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4472),
.B(n_351),
.Y(n_4632)
);

CKINVDCx5p33_ASAP7_75t_R g4633 ( 
.A(n_4506),
.Y(n_4633)
);

OAI211xp5_ASAP7_75t_SL g4634 ( 
.A1(n_4387),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_4634)
);

AOI21xp5_ASAP7_75t_L g4635 ( 
.A1(n_4458),
.A2(n_353),
.B(n_355),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4477),
.Y(n_4636)
);

AOI22xp33_ASAP7_75t_L g4637 ( 
.A1(n_4462),
.A2(n_4395),
.B1(n_4394),
.B2(n_4401),
.Y(n_4637)
);

AO221x2_ASAP7_75t_L g4638 ( 
.A1(n_4358),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.C(n_359),
.Y(n_4638)
);

OAI21xp33_ASAP7_75t_L g4639 ( 
.A1(n_4437),
.A2(n_359),
.B(n_360),
.Y(n_4639)
);

INVx3_ASAP7_75t_L g4640 ( 
.A(n_4462),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4479),
.B(n_360),
.Y(n_4641)
);

OAI21x1_ASAP7_75t_L g4642 ( 
.A1(n_4358),
.A2(n_361),
.B(n_362),
.Y(n_4642)
);

CKINVDCx5p33_ASAP7_75t_R g4643 ( 
.A(n_4492),
.Y(n_4643)
);

AOI322xp5_ASAP7_75t_L g4644 ( 
.A1(n_4499),
.A2(n_361),
.A3(n_363),
.B1(n_364),
.B2(n_365),
.C1(n_366),
.C2(n_367),
.Y(n_4644)
);

OAI21xp33_ASAP7_75t_L g4645 ( 
.A1(n_4437),
.A2(n_363),
.B(n_364),
.Y(n_4645)
);

AOI221xp5_ASAP7_75t_L g4646 ( 
.A1(n_4447),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.C(n_368),
.Y(n_4646)
);

AOI221xp5_ASAP7_75t_L g4647 ( 
.A1(n_4407),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.C(n_371),
.Y(n_4647)
);

OAI211xp5_ASAP7_75t_L g4648 ( 
.A1(n_4401),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_4492),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4407),
.Y(n_4650)
);

A2O1A1Ixp33_ASAP7_75t_L g4651 ( 
.A1(n_4362),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4479),
.B(n_4399),
.Y(n_4652)
);

OAI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4461),
.A2(n_4478),
.B(n_4362),
.Y(n_4653)
);

OAI21x1_ASAP7_75t_L g4654 ( 
.A1(n_4359),
.A2(n_374),
.B(n_375),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4594),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4519),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4598),
.Y(n_4657)
);

INVxp67_ASAP7_75t_SL g4658 ( 
.A(n_4573),
.Y(n_4658)
);

INVx2_ASAP7_75t_L g4659 ( 
.A(n_4598),
.Y(n_4659)
);

INVxp67_ASAP7_75t_L g4660 ( 
.A(n_4513),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4650),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4532),
.Y(n_4662)
);

INVxp67_ASAP7_75t_L g4663 ( 
.A(n_4621),
.Y(n_4663)
);

AND2x2_ASAP7_75t_L g4664 ( 
.A(n_4516),
.B(n_4359),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4598),
.Y(n_4665)
);

INVx2_ASAP7_75t_SL g4666 ( 
.A(n_4600),
.Y(n_4666)
);

OR2x2_ASAP7_75t_L g4667 ( 
.A(n_4520),
.B(n_4415),
.Y(n_4667)
);

BUFx2_ASAP7_75t_L g4668 ( 
.A(n_4549),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4536),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4538),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4600),
.Y(n_4671)
);

NOR2x1p5_ASAP7_75t_L g4672 ( 
.A(n_4535),
.B(n_4496),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4525),
.B(n_4408),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4525),
.B(n_4476),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4575),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4561),
.B(n_4480),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4600),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4578),
.Y(n_4678)
);

OR2x6_ASAP7_75t_L g4679 ( 
.A(n_4521),
.B(n_4496),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4620),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4561),
.B(n_4361),
.Y(n_4681)
);

BUFx2_ASAP7_75t_L g4682 ( 
.A(n_4572),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4515),
.B(n_4481),
.Y(n_4683)
);

OR2x2_ASAP7_75t_L g4684 ( 
.A(n_4562),
.B(n_4415),
.Y(n_4684)
);

AND2x2_ASAP7_75t_L g4685 ( 
.A(n_4559),
.B(n_4361),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4620),
.B(n_4368),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4511),
.B(n_4368),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4550),
.B(n_4446),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4584),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4512),
.B(n_4517),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4587),
.B(n_4446),
.Y(n_4691)
);

INVx2_ASAP7_75t_L g4692 ( 
.A(n_4612),
.Y(n_4692)
);

OR2x2_ASAP7_75t_L g4693 ( 
.A(n_4602),
.B(n_4505),
.Y(n_4693)
);

BUFx2_ASAP7_75t_L g4694 ( 
.A(n_4593),
.Y(n_4694)
);

INVx2_ASAP7_75t_L g4695 ( 
.A(n_4621),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4526),
.B(n_4384),
.Y(n_4696)
);

OR2x2_ASAP7_75t_L g4697 ( 
.A(n_4564),
.B(n_4505),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4586),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4652),
.B(n_4640),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4588),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4623),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4570),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4640),
.B(n_4355),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4539),
.B(n_4401),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4539),
.B(n_4543),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4570),
.Y(n_4706)
);

INVx2_ASAP7_75t_L g4707 ( 
.A(n_4540),
.Y(n_4707)
);

AND2x2_ASAP7_75t_L g4708 ( 
.A(n_4535),
.B(n_4494),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4514),
.B(n_4464),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4624),
.Y(n_4710)
);

BUFx2_ASAP7_75t_L g4711 ( 
.A(n_4542),
.Y(n_4711)
);

AND2x4_ASAP7_75t_L g4712 ( 
.A(n_4629),
.B(n_4355),
.Y(n_4712)
);

INVx5_ASAP7_75t_L g4713 ( 
.A(n_4540),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4632),
.Y(n_4714)
);

OR2x2_ASAP7_75t_L g4715 ( 
.A(n_4631),
.B(n_4420),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4641),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4574),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4636),
.B(n_4420),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4540),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4528),
.B(n_4497),
.Y(n_4720)
);

BUFx2_ASAP7_75t_L g4721 ( 
.A(n_4524),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4556),
.Y(n_4722)
);

OR2x2_ASAP7_75t_L g4723 ( 
.A(n_4626),
.B(n_4422),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4653),
.B(n_4384),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4556),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4610),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4529),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4533),
.Y(n_4728)
);

INVx2_ASAP7_75t_L g4729 ( 
.A(n_4552),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4653),
.B(n_4422),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4581),
.B(n_4439),
.Y(n_4731)
);

BUFx3_ASAP7_75t_L g4732 ( 
.A(n_4608),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4558),
.B(n_4398),
.Y(n_4733)
);

NOR2xp33_ASAP7_75t_L g4734 ( 
.A(n_4630),
.B(n_4487),
.Y(n_4734)
);

CKINVDCx10_ASAP7_75t_R g4735 ( 
.A(n_4605),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4637),
.B(n_4423),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4596),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4609),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4617),
.Y(n_4739)
);

AOI22xp33_ASAP7_75t_SL g4740 ( 
.A1(n_4522),
.A2(n_4461),
.B1(n_4379),
.B2(n_4443),
.Y(n_4740)
);

NOR2x1_ASAP7_75t_SL g4741 ( 
.A(n_4648),
.B(n_4522),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4619),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_4638),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4523),
.B(n_4439),
.Y(n_4744)
);

HB1xp67_ASAP7_75t_L g4745 ( 
.A(n_4638),
.Y(n_4745)
);

OR2x2_ASAP7_75t_L g4746 ( 
.A(n_4518),
.B(n_4423),
.Y(n_4746)
);

INVx2_ASAP7_75t_SL g4747 ( 
.A(n_4643),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4576),
.B(n_4449),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4568),
.B(n_4382),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4616),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4530),
.B(n_4431),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4554),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4604),
.B(n_4431),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4585),
.B(n_4386),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4555),
.B(n_4432),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4537),
.B(n_4432),
.Y(n_4756)
);

HB1xp67_ASAP7_75t_L g4757 ( 
.A(n_4592),
.Y(n_4757)
);

BUFx2_ASAP7_75t_L g4758 ( 
.A(n_4649),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4633),
.B(n_4449),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4625),
.Y(n_4760)
);

OR2x2_ASAP7_75t_L g4761 ( 
.A(n_4589),
.B(n_4456),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4527),
.B(n_4456),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4541),
.B(n_4467),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_4642),
.B(n_4467),
.Y(n_4764)
);

HB1xp67_ASAP7_75t_L g4765 ( 
.A(n_4635),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4654),
.B(n_4400),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4546),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4758),
.B(n_4417),
.Y(n_4768)
);

BUFx3_ASAP7_75t_L g4769 ( 
.A(n_4668),
.Y(n_4769)
);

AND2x2_ASAP7_75t_L g4770 ( 
.A(n_4747),
.B(n_4417),
.Y(n_4770)
);

OAI22xp5_ASAP7_75t_L g4771 ( 
.A1(n_4658),
.A2(n_4534),
.B1(n_4548),
.B2(n_4651),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4682),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4713),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4747),
.B(n_4418),
.Y(n_4774)
);

OR2x2_ASAP7_75t_L g4775 ( 
.A(n_4722),
.B(n_4418),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4713),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4743),
.B(n_4544),
.Y(n_4777)
);

INVx2_ASAP7_75t_L g4778 ( 
.A(n_4713),
.Y(n_4778)
);

INVx3_ASAP7_75t_L g4779 ( 
.A(n_4713),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4673),
.B(n_4400),
.Y(n_4780)
);

OR2x2_ASAP7_75t_L g4781 ( 
.A(n_4725),
.B(n_4356),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4732),
.Y(n_4782)
);

INVx2_ASAP7_75t_SL g4783 ( 
.A(n_4735),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4732),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4694),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4699),
.B(n_4402),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4743),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4699),
.B(n_4402),
.Y(n_4788)
);

BUFx2_ASAP7_75t_L g4789 ( 
.A(n_4745),
.Y(n_4789)
);

BUFx2_ASAP7_75t_L g4790 ( 
.A(n_4745),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4741),
.B(n_4560),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4658),
.B(n_4551),
.Y(n_4792)
);

INVx4_ASAP7_75t_L g4793 ( 
.A(n_4711),
.Y(n_4793)
);

OAI22xp5_ASAP7_75t_L g4794 ( 
.A1(n_4740),
.A2(n_4571),
.B1(n_4557),
.B2(n_4614),
.Y(n_4794)
);

INVx2_ASAP7_75t_L g4795 ( 
.A(n_4672),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4663),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4660),
.B(n_4545),
.Y(n_4797)
);

INVx2_ASAP7_75t_L g4798 ( 
.A(n_4666),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4663),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4666),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4695),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_4705),
.B(n_4707),
.Y(n_4802)
);

OR2x2_ASAP7_75t_L g4803 ( 
.A(n_4738),
.B(n_4356),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4686),
.Y(n_4804)
);

INVx2_ASAP7_75t_L g4805 ( 
.A(n_4686),
.Y(n_4805)
);

NOR2x1_ASAP7_75t_L g4806 ( 
.A(n_4695),
.B(n_4580),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4702),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4660),
.B(n_4545),
.Y(n_4808)
);

AOI22xp33_ASAP7_75t_L g4809 ( 
.A1(n_4690),
.A2(n_4531),
.B1(n_4553),
.B2(n_4591),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4707),
.B(n_4371),
.Y(n_4810)
);

BUFx2_ASAP7_75t_L g4811 ( 
.A(n_4679),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4726),
.B(n_4657),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4706),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_4686),
.Y(n_4814)
);

INVx2_ASAP7_75t_L g4815 ( 
.A(n_4703),
.Y(n_4815)
);

AND2x2_ASAP7_75t_L g4816 ( 
.A(n_4719),
.B(n_4371),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4703),
.Y(n_4817)
);

HB1xp67_ASAP7_75t_L g4818 ( 
.A(n_4679),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_4719),
.B(n_4378),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4703),
.Y(n_4820)
);

NOR2x1_ASAP7_75t_L g4821 ( 
.A(n_4679),
.B(n_4580),
.Y(n_4821)
);

INVx2_ASAP7_75t_L g4822 ( 
.A(n_4664),
.Y(n_4822)
);

OR2x2_ASAP7_75t_L g4823 ( 
.A(n_4738),
.B(n_4357),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_SL g4824 ( 
.A(n_4740),
.B(n_4622),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4661),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4656),
.Y(n_4826)
);

BUFx2_ASAP7_75t_L g4827 ( 
.A(n_4726),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4685),
.B(n_4378),
.Y(n_4828)
);

INVx1_ASAP7_75t_SL g4829 ( 
.A(n_4708),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4685),
.B(n_4657),
.Y(n_4830)
);

OR2x2_ASAP7_75t_L g4831 ( 
.A(n_4655),
.B(n_4357),
.Y(n_4831)
);

INVx3_ASAP7_75t_L g4832 ( 
.A(n_4712),
.Y(n_4832)
);

AND2x2_ASAP7_75t_L g4833 ( 
.A(n_4659),
.B(n_4406),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4659),
.B(n_4567),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4662),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4665),
.B(n_4547),
.Y(n_4836)
);

HB1xp67_ASAP7_75t_L g4837 ( 
.A(n_4665),
.Y(n_4837)
);

NOR2xp67_ASAP7_75t_L g4838 ( 
.A(n_4727),
.B(n_4443),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4765),
.Y(n_4839)
);

BUFx12f_ASAP7_75t_L g4840 ( 
.A(n_4721),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4769),
.B(n_4671),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4789),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4789),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4790),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4790),
.Y(n_4845)
);

OR2x2_ASAP7_75t_L g4846 ( 
.A(n_4785),
.B(n_4760),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4827),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4832),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4827),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4837),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4832),
.Y(n_4851)
);

INVx5_ASAP7_75t_SL g4852 ( 
.A(n_4773),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4824),
.B(n_4757),
.Y(n_4853)
);

NAND2x1_ASAP7_75t_L g4854 ( 
.A(n_4779),
.B(n_4664),
.Y(n_4854)
);

AND2x4_ASAP7_75t_L g4855 ( 
.A(n_4793),
.B(n_4671),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4832),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4772),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4769),
.B(n_4677),
.Y(n_4858)
);

OR2x2_ASAP7_75t_L g4859 ( 
.A(n_4785),
.B(n_4746),
.Y(n_4859)
);

AND2x2_ASAP7_75t_L g4860 ( 
.A(n_4802),
.B(n_4677),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4802),
.B(n_4759),
.Y(n_4861)
);

AOI22xp5_ASAP7_75t_L g4862 ( 
.A1(n_4771),
.A2(n_4794),
.B1(n_4809),
.B2(n_4791),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4779),
.Y(n_4863)
);

HB1xp67_ASAP7_75t_L g4864 ( 
.A(n_4806),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4779),
.Y(n_4865)
);

OR2x2_ASAP7_75t_L g4866 ( 
.A(n_4787),
.B(n_4684),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4782),
.B(n_4692),
.Y(n_4867)
);

AND2x2_ASAP7_75t_L g4868 ( 
.A(n_4782),
.B(n_4692),
.Y(n_4868)
);

AND2x2_ASAP7_75t_L g4869 ( 
.A(n_4784),
.B(n_4727),
.Y(n_4869)
);

HB1xp67_ASAP7_75t_L g4870 ( 
.A(n_4806),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4772),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4801),
.Y(n_4872)
);

HB1xp67_ASAP7_75t_L g4873 ( 
.A(n_4787),
.Y(n_4873)
);

INVx3_ASAP7_75t_L g4874 ( 
.A(n_4793),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4784),
.B(n_4720),
.Y(n_4875)
);

HB1xp67_ASAP7_75t_L g4876 ( 
.A(n_4839),
.Y(n_4876)
);

INVxp33_ASAP7_75t_SL g4877 ( 
.A(n_4818),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4793),
.Y(n_4878)
);

OR2x2_ASAP7_75t_L g4879 ( 
.A(n_4829),
.B(n_4757),
.Y(n_4879)
);

OAI321xp33_ASAP7_75t_L g4880 ( 
.A1(n_4792),
.A2(n_4777),
.A3(n_4808),
.B1(n_4797),
.B2(n_4751),
.C(n_4811),
.Y(n_4880)
);

AOI221xp5_ASAP7_75t_L g4881 ( 
.A1(n_4839),
.A2(n_4765),
.B1(n_4683),
.B2(n_4751),
.C(n_4767),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4783),
.B(n_4748),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4801),
.Y(n_4883)
);

INVx4_ASAP7_75t_L g4884 ( 
.A(n_4840),
.Y(n_4884)
);

OR2x2_ASAP7_75t_L g4885 ( 
.A(n_4829),
.B(n_4667),
.Y(n_4885)
);

AND2x4_ASAP7_75t_L g4886 ( 
.A(n_4804),
.B(n_4680),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4831),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4831),
.Y(n_4888)
);

AND2x2_ASAP7_75t_L g4889 ( 
.A(n_4783),
.B(n_4830),
.Y(n_4889)
);

INVx2_ASAP7_75t_SL g4890 ( 
.A(n_4815),
.Y(n_4890)
);

OR2x2_ASAP7_75t_L g4891 ( 
.A(n_4812),
.B(n_4710),
.Y(n_4891)
);

AOI22xp33_ASAP7_75t_L g4892 ( 
.A1(n_4821),
.A2(n_4763),
.B1(n_4744),
.B2(n_4756),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4796),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4796),
.Y(n_4894)
);

BUFx3_ASAP7_75t_L g4895 ( 
.A(n_4840),
.Y(n_4895)
);

AOI22xp5_ASAP7_75t_L g4896 ( 
.A1(n_4821),
.A2(n_4733),
.B1(n_4749),
.B2(n_4756),
.Y(n_4896)
);

INVx4_ASAP7_75t_L g4897 ( 
.A(n_4773),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4799),
.Y(n_4898)
);

OR2x2_ASAP7_75t_L g4899 ( 
.A(n_4836),
.B(n_4714),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4799),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4864),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4889),
.B(n_4830),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4864),
.Y(n_4903)
);

NAND4xp25_ASAP7_75t_L g4904 ( 
.A(n_4862),
.B(n_4795),
.C(n_4834),
.D(n_4811),
.Y(n_4904)
);

NOR2xp33_ASAP7_75t_L g4905 ( 
.A(n_4884),
.B(n_4795),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4860),
.B(n_4768),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4870),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4870),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4882),
.B(n_4768),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4895),
.B(n_4822),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4841),
.B(n_4798),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4895),
.B(n_4822),
.Y(n_4912)
);

OR2x2_ASAP7_75t_L g4913 ( 
.A(n_4879),
.B(n_4680),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4844),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4884),
.B(n_4798),
.Y(n_4915)
);

AND3x1_ASAP7_75t_L g4916 ( 
.A(n_4881),
.B(n_4774),
.C(n_4770),
.Y(n_4916)
);

AND2x4_ASAP7_75t_L g4917 ( 
.A(n_4844),
.B(n_4804),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4861),
.B(n_4800),
.Y(n_4918)
);

HB1xp67_ASAP7_75t_L g4919 ( 
.A(n_4873),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4876),
.Y(n_4920)
);

OR2x2_ASAP7_75t_L g4921 ( 
.A(n_4853),
.B(n_4803),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_4858),
.B(n_4800),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4875),
.B(n_4770),
.Y(n_4923)
);

AND2x2_ASAP7_75t_L g4924 ( 
.A(n_4867),
.B(n_4774),
.Y(n_4924)
);

AND2x4_ASAP7_75t_SL g4925 ( 
.A(n_4855),
.B(n_4776),
.Y(n_4925)
);

OR2x2_ASAP7_75t_L g4926 ( 
.A(n_4853),
.B(n_4803),
.Y(n_4926)
);

AND2x2_ASAP7_75t_L g4927 ( 
.A(n_4868),
.B(n_4780),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4869),
.B(n_4780),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4876),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4855),
.B(n_4691),
.Y(n_4930)
);

INVxp67_ASAP7_75t_SL g4931 ( 
.A(n_4874),
.Y(n_4931)
);

AND2x4_ASAP7_75t_L g4932 ( 
.A(n_4848),
.B(n_4805),
.Y(n_4932)
);

OR2x2_ASAP7_75t_L g4933 ( 
.A(n_4842),
.B(n_4823),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4854),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4873),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4874),
.B(n_4691),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4852),
.B(n_4762),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4877),
.B(n_4838),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4877),
.B(n_4838),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4852),
.B(n_4786),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4852),
.B(n_4786),
.Y(n_4941)
);

INVx3_ASAP7_75t_L g4942 ( 
.A(n_4897),
.Y(n_4942)
);

HB1xp67_ASAP7_75t_L g4943 ( 
.A(n_4843),
.Y(n_4943)
);

AND2x2_ASAP7_75t_SL g4944 ( 
.A(n_4881),
.B(n_4823),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4892),
.B(n_4752),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4845),
.Y(n_4946)
);

HB1xp67_ASAP7_75t_L g4947 ( 
.A(n_4848),
.Y(n_4947)
);

OR2x2_ASAP7_75t_L g4948 ( 
.A(n_4847),
.B(n_4781),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4851),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4886),
.B(n_4788),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4851),
.Y(n_4951)
);

AND2x2_ASAP7_75t_L g4952 ( 
.A(n_4886),
.B(n_4788),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4856),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4878),
.B(n_4696),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4856),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4863),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4919),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4947),
.Y(n_4958)
);

AND2x2_ASAP7_75t_L g4959 ( 
.A(n_4902),
.B(n_4739),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4902),
.B(n_4742),
.Y(n_4960)
);

OR2x2_ASAP7_75t_L g4961 ( 
.A(n_4906),
.B(n_4846),
.Y(n_4961)
);

AND2x2_ASAP7_75t_L g4962 ( 
.A(n_4909),
.B(n_4750),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4920),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4909),
.B(n_4716),
.Y(n_4964)
);

AND2x4_ASAP7_75t_L g4965 ( 
.A(n_4925),
.B(n_4878),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4944),
.B(n_4942),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4918),
.B(n_4927),
.Y(n_4967)
);

OR2x2_ASAP7_75t_L g4968 ( 
.A(n_4921),
.B(n_4885),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4929),
.Y(n_4969)
);

NAND2x1p5_ASAP7_75t_L g4970 ( 
.A(n_4942),
.B(n_4897),
.Y(n_4970)
);

OR2x2_ASAP7_75t_L g4971 ( 
.A(n_4921),
.B(n_4859),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4935),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4944),
.B(n_4849),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4932),
.Y(n_4974)
);

AND2x4_ASAP7_75t_L g4975 ( 
.A(n_4925),
.B(n_4890),
.Y(n_4975)
);

AOI22xp5_ASAP7_75t_L g4976 ( 
.A1(n_4916),
.A2(n_4896),
.B1(n_4892),
.B2(n_4709),
.Y(n_4976)
);

OR2x2_ASAP7_75t_L g4977 ( 
.A(n_4926),
.B(n_4866),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4942),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4918),
.B(n_4850),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4917),
.B(n_4863),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4932),
.Y(n_4981)
);

AND2x2_ASAP7_75t_L g4982 ( 
.A(n_4927),
.B(n_4734),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4928),
.B(n_4734),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4928),
.B(n_4755),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4924),
.B(n_4755),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4917),
.B(n_4865),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4917),
.B(n_4865),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4932),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4931),
.B(n_4887),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4924),
.B(n_4696),
.Y(n_4990)
);

AND2x2_ASAP7_75t_L g4991 ( 
.A(n_4930),
.B(n_4753),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4914),
.B(n_4888),
.Y(n_4992)
);

AND2x2_ASAP7_75t_L g4993 ( 
.A(n_4930),
.B(n_4753),
.Y(n_4993)
);

NAND2x1p5_ASAP7_75t_L g4994 ( 
.A(n_4915),
.B(n_4776),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4933),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4933),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4956),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4914),
.B(n_4857),
.Y(n_4998)
);

OR2x2_ASAP7_75t_L g4999 ( 
.A(n_4926),
.B(n_4899),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4937),
.B(n_4778),
.Y(n_5000)
);

OAI211xp5_ASAP7_75t_L g5001 ( 
.A1(n_4938),
.A2(n_4644),
.B(n_4622),
.C(n_4647),
.Y(n_5001)
);

AND2x4_ASAP7_75t_L g5002 ( 
.A(n_4940),
.B(n_4778),
.Y(n_5002)
);

OR2x2_ASAP7_75t_L g5003 ( 
.A(n_4913),
.B(n_4923),
.Y(n_5003)
);

OR2x2_ASAP7_75t_L g5004 ( 
.A(n_4911),
.B(n_4891),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4937),
.B(n_4717),
.Y(n_5005)
);

BUFx3_ASAP7_75t_L g5006 ( 
.A(n_4940),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4967),
.B(n_4950),
.Y(n_5007)
);

AND2x2_ASAP7_75t_L g5008 ( 
.A(n_4982),
.B(n_4950),
.Y(n_5008)
);

INVx2_ASAP7_75t_L g5009 ( 
.A(n_4994),
.Y(n_5009)
);

OAI22xp33_ASAP7_75t_L g5010 ( 
.A1(n_4976),
.A2(n_4880),
.B1(n_4939),
.B2(n_4697),
.Y(n_5010)
);

AND2x2_ASAP7_75t_L g5011 ( 
.A(n_4983),
.B(n_4952),
.Y(n_5011)
);

AND2x4_ASAP7_75t_L g5012 ( 
.A(n_4975),
.B(n_4934),
.Y(n_5012)
);

BUFx3_ASAP7_75t_L g5013 ( 
.A(n_4975),
.Y(n_5013)
);

OR2x2_ASAP7_75t_L g5014 ( 
.A(n_4971),
.B(n_4922),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4994),
.Y(n_5015)
);

NAND4xp75_ASAP7_75t_L g5016 ( 
.A(n_4973),
.B(n_4915),
.C(n_4910),
.D(n_4912),
.Y(n_5016)
);

HB1xp67_ASAP7_75t_L g5017 ( 
.A(n_4966),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4974),
.B(n_4981),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4988),
.Y(n_5019)
);

INVx2_ASAP7_75t_L g5020 ( 
.A(n_4970),
.Y(n_5020)
);

AND2x2_ASAP7_75t_L g5021 ( 
.A(n_4990),
.B(n_4952),
.Y(n_5021)
);

INVx2_ASAP7_75t_L g5022 ( 
.A(n_4970),
.Y(n_5022)
);

AND2x4_ASAP7_75t_SL g5023 ( 
.A(n_4991),
.B(n_4941),
.Y(n_5023)
);

INVx2_ASAP7_75t_SL g5024 ( 
.A(n_4965),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4976),
.B(n_4907),
.Y(n_5025)
);

OR2x2_ASAP7_75t_L g5026 ( 
.A(n_4977),
.B(n_4945),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4979),
.B(n_4907),
.Y(n_5027)
);

OR2x2_ASAP7_75t_L g5028 ( 
.A(n_4968),
.B(n_4973),
.Y(n_5028)
);

NAND2xp5_ASAP7_75t_L g5029 ( 
.A(n_4985),
.B(n_4908),
.Y(n_5029)
);

INVx2_ASAP7_75t_SL g5030 ( 
.A(n_4965),
.Y(n_5030)
);

AND2x2_ASAP7_75t_L g5031 ( 
.A(n_4993),
.B(n_4941),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4995),
.B(n_4908),
.Y(n_5032)
);

OR2x2_ASAP7_75t_L g5033 ( 
.A(n_4999),
.B(n_4948),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4980),
.Y(n_5034)
);

NAND3xp33_ASAP7_75t_SL g5035 ( 
.A(n_4966),
.B(n_4903),
.C(n_4901),
.Y(n_5035)
);

INVx2_ASAP7_75t_SL g5036 ( 
.A(n_5006),
.Y(n_5036)
);

HB1xp67_ASAP7_75t_L g5037 ( 
.A(n_4980),
.Y(n_5037)
);

BUFx2_ASAP7_75t_L g5038 ( 
.A(n_4996),
.Y(n_5038)
);

OAI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_5001),
.A2(n_4880),
.B(n_4904),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_4986),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4984),
.B(n_4954),
.Y(n_5041)
);

AND2x2_ASAP7_75t_L g5042 ( 
.A(n_4962),
.B(n_4910),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4959),
.B(n_4912),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4960),
.B(n_4936),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4986),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4964),
.B(n_4936),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4987),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4987),
.Y(n_5048)
);

INVx1_ASAP7_75t_SL g5049 ( 
.A(n_5000),
.Y(n_5049)
);

BUFx2_ASAP7_75t_L g5050 ( 
.A(n_5002),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_5002),
.Y(n_5051)
);

INVx1_ASAP7_75t_SL g5052 ( 
.A(n_4989),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4989),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4978),
.B(n_4954),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4992),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4958),
.B(n_4956),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_5005),
.B(n_4943),
.Y(n_5057)
);

AOI22xp5_ASAP7_75t_L g5058 ( 
.A1(n_4957),
.A2(n_4905),
.B1(n_4736),
.B2(n_4676),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4992),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_5024),
.B(n_4934),
.Y(n_5060)
);

AND2x2_ASAP7_75t_L g5061 ( 
.A(n_5007),
.B(n_5003),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5030),
.B(n_4871),
.Y(n_5062)
);

NOR3xp33_ASAP7_75t_SL g5063 ( 
.A(n_5010),
.B(n_4946),
.C(n_4998),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_5012),
.B(n_4949),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_5050),
.Y(n_5065)
);

AND2x2_ASAP7_75t_L g5066 ( 
.A(n_5008),
.B(n_4961),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_5012),
.B(n_4951),
.Y(n_5067)
);

HB1xp67_ASAP7_75t_L g5068 ( 
.A(n_5013),
.Y(n_5068)
);

AOI22xp5_ASAP7_75t_L g5069 ( 
.A1(n_5039),
.A2(n_5025),
.B1(n_5035),
.B2(n_5052),
.Y(n_5069)
);

NOR2x1_ASAP7_75t_L g5070 ( 
.A(n_5016),
.B(n_4998),
.Y(n_5070)
);

OAI322xp33_ASAP7_75t_L g5071 ( 
.A1(n_5025),
.A2(n_4826),
.A3(n_4948),
.B1(n_4825),
.B2(n_4900),
.C1(n_4893),
.C2(n_4894),
.Y(n_5071)
);

OA222x2_ASAP7_75t_L g5072 ( 
.A1(n_5028),
.A2(n_4898),
.B1(n_4997),
.B2(n_4963),
.C1(n_4972),
.C2(n_4969),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_5033),
.Y(n_5073)
);

AOI211xp5_ASAP7_75t_L g5074 ( 
.A1(n_5039),
.A2(n_5035),
.B(n_5052),
.C(n_5017),
.Y(n_5074)
);

AOI22xp5_ASAP7_75t_L g5075 ( 
.A1(n_5049),
.A2(n_4826),
.B1(n_4807),
.B2(n_4813),
.Y(n_5075)
);

A2O1A1Ixp33_ASAP7_75t_L g5076 ( 
.A1(n_5017),
.A2(n_4736),
.B(n_4781),
.C(n_4805),
.Y(n_5076)
);

AND2x2_ASAP7_75t_L g5077 ( 
.A(n_5011),
.B(n_5004),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_5049),
.B(n_4953),
.Y(n_5078)
);

INVx2_ASAP7_75t_L g5079 ( 
.A(n_5009),
.Y(n_5079)
);

NOR2xp33_ASAP7_75t_SL g5080 ( 
.A(n_5042),
.B(n_4814),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_5015),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_5043),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5044),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5046),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_5051),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_5027),
.Y(n_5086)
);

NAND2x1_ASAP7_75t_L g5087 ( 
.A(n_5038),
.B(n_4814),
.Y(n_5087)
);

HB1xp67_ASAP7_75t_L g5088 ( 
.A(n_5037),
.Y(n_5088)
);

NOR2xp33_ASAP7_75t_L g5089 ( 
.A(n_5023),
.B(n_4825),
.Y(n_5089)
);

NAND2x1_ASAP7_75t_L g5090 ( 
.A(n_5021),
.B(n_4815),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_5031),
.B(n_4955),
.Y(n_5091)
);

HB1xp67_ASAP7_75t_L g5092 ( 
.A(n_5057),
.Y(n_5092)
);

NAND2x1p5_ASAP7_75t_L g5093 ( 
.A(n_5036),
.B(n_4817),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_5027),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_5014),
.Y(n_5095)
);

NAND2xp5_ASAP7_75t_L g5096 ( 
.A(n_5058),
.B(n_4817),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5057),
.Y(n_5097)
);

INVx3_ASAP7_75t_SL g5098 ( 
.A(n_5020),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5041),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_5041),
.Y(n_5100)
);

INVx2_ASAP7_75t_SL g5101 ( 
.A(n_5022),
.Y(n_5101)
);

AO22x1_ASAP7_75t_L g5102 ( 
.A1(n_5019),
.A2(n_4872),
.B1(n_4883),
.B2(n_4820),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5029),
.Y(n_5103)
);

AOI211xp5_ASAP7_75t_L g5104 ( 
.A1(n_5026),
.A2(n_4813),
.B(n_4807),
.C(n_4606),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5029),
.Y(n_5105)
);

AND2x2_ASAP7_75t_L g5106 ( 
.A(n_5053),
.B(n_4674),
.Y(n_5106)
);

AND2x2_ASAP7_75t_L g5107 ( 
.A(n_5061),
.B(n_5054),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_5066),
.B(n_5054),
.Y(n_5108)
);

BUFx2_ASAP7_75t_L g5109 ( 
.A(n_5093),
.Y(n_5109)
);

AO21x2_ASAP7_75t_L g5110 ( 
.A1(n_5069),
.A2(n_5032),
.B(n_5056),
.Y(n_5110)
);

CKINVDCx16_ASAP7_75t_R g5111 ( 
.A(n_5077),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_5068),
.B(n_5034),
.Y(n_5112)
);

AND2x2_ASAP7_75t_L g5113 ( 
.A(n_5091),
.B(n_5082),
.Y(n_5113)
);

INVx4_ASAP7_75t_L g5114 ( 
.A(n_5098),
.Y(n_5114)
);

OR2x2_ASAP7_75t_L g5115 ( 
.A(n_5087),
.B(n_5018),
.Y(n_5115)
);

INVx2_ASAP7_75t_SL g5116 ( 
.A(n_5090),
.Y(n_5116)
);

OR2x2_ASAP7_75t_L g5117 ( 
.A(n_5060),
.B(n_5018),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5064),
.Y(n_5118)
);

INVx2_ASAP7_75t_L g5119 ( 
.A(n_5065),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_5067),
.Y(n_5120)
);

NAND3xp33_ASAP7_75t_L g5121 ( 
.A(n_5074),
.B(n_5032),
.C(n_5056),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_5069),
.Y(n_5122)
);

OR2x2_ASAP7_75t_L g5123 ( 
.A(n_5062),
.B(n_5040),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_5076),
.B(n_5045),
.Y(n_5124)
);

BUFx2_ASAP7_75t_L g5125 ( 
.A(n_5088),
.Y(n_5125)
);

OR2x2_ASAP7_75t_L g5126 ( 
.A(n_5073),
.B(n_5047),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_5083),
.B(n_5048),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_L g5128 ( 
.A(n_5080),
.B(n_5055),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_5074),
.Y(n_5129)
);

NAND4xp25_ASAP7_75t_L g5130 ( 
.A(n_5084),
.B(n_5059),
.C(n_4835),
.D(n_4820),
.Y(n_5130)
);

CKINVDCx5p33_ASAP7_75t_R g5131 ( 
.A(n_5063),
.Y(n_5131)
);

OR2x2_ASAP7_75t_L g5132 ( 
.A(n_5078),
.B(n_4775),
.Y(n_5132)
);

OAI22xp33_ASAP7_75t_L g5133 ( 
.A1(n_5096),
.A2(n_4693),
.B1(n_4728),
.B2(n_4775),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5070),
.Y(n_5134)
);

OR2x2_ASAP7_75t_L g5135 ( 
.A(n_5085),
.B(n_4835),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_5089),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_L g5137 ( 
.A(n_5102),
.B(n_4833),
.Y(n_5137)
);

AND2x2_ASAP7_75t_L g5138 ( 
.A(n_5106),
.B(n_4688),
.Y(n_5138)
);

AND2x4_ASAP7_75t_L g5139 ( 
.A(n_5095),
.B(n_4833),
.Y(n_5139)
);

HB1xp67_ASAP7_75t_L g5140 ( 
.A(n_5092),
.Y(n_5140)
);

AND2x2_ASAP7_75t_L g5141 ( 
.A(n_5101),
.B(n_4688),
.Y(n_5141)
);

AND2x4_ASAP7_75t_L g5142 ( 
.A(n_5079),
.B(n_4810),
.Y(n_5142)
);

AND2x2_ASAP7_75t_L g5143 ( 
.A(n_5081),
.B(n_4687),
.Y(n_5143)
);

NAND2xp5_ASAP7_75t_L g5144 ( 
.A(n_5103),
.B(n_4810),
.Y(n_5144)
);

OR2x2_ASAP7_75t_L g5145 ( 
.A(n_5105),
.B(n_5086),
.Y(n_5145)
);

BUFx3_ASAP7_75t_L g5146 ( 
.A(n_5109),
.Y(n_5146)
);

NOR2xp33_ASAP7_75t_L g5147 ( 
.A(n_5111),
.B(n_5094),
.Y(n_5147)
);

OAI221xp5_ASAP7_75t_L g5148 ( 
.A1(n_5122),
.A2(n_5104),
.B1(n_5097),
.B2(n_5100),
.C(n_5099),
.Y(n_5148)
);

INVx3_ASAP7_75t_L g5149 ( 
.A(n_5114),
.Y(n_5149)
);

INVx2_ASAP7_75t_L g5150 ( 
.A(n_5115),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_5116),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5137),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_5142),
.B(n_5104),
.Y(n_5153)
);

NOR2xp33_ASAP7_75t_SL g5154 ( 
.A(n_5114),
.B(n_5072),
.Y(n_5154)
);

INVx1_ASAP7_75t_SL g5155 ( 
.A(n_5110),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_5141),
.Y(n_5156)
);

INVx3_ASAP7_75t_SL g5157 ( 
.A(n_5126),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_5143),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_5108),
.B(n_5107),
.Y(n_5159)
);

HB1xp67_ASAP7_75t_L g5160 ( 
.A(n_5110),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5142),
.B(n_5139),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_5138),
.Y(n_5162)
);

INVx1_ASAP7_75t_SL g5163 ( 
.A(n_5125),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_5139),
.B(n_5075),
.Y(n_5164)
);

AOI21xp5_ASAP7_75t_L g5165 ( 
.A1(n_5121),
.A2(n_5071),
.B(n_5072),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5113),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_5140),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_5132),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_5112),
.B(n_4687),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_5134),
.B(n_5075),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_5117),
.Y(n_5171)
);

AND2x4_ASAP7_75t_L g5172 ( 
.A(n_5119),
.B(n_4816),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_5134),
.Y(n_5173)
);

AND2x2_ASAP7_75t_L g5174 ( 
.A(n_5127),
.B(n_4816),
.Y(n_5174)
);

INVx2_ASAP7_75t_SL g5175 ( 
.A(n_5135),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_5128),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_5145),
.Y(n_5177)
);

NOR2x1_ASAP7_75t_L g5178 ( 
.A(n_5122),
.B(n_4819),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5144),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5160),
.Y(n_5180)
);

NOR4xp25_ASAP7_75t_SL g5181 ( 
.A(n_5148),
.B(n_5131),
.C(n_5129),
.D(n_5136),
.Y(n_5181)
);

AO22x1_ASAP7_75t_L g5182 ( 
.A1(n_5155),
.A2(n_5129),
.B1(n_5136),
.B2(n_5118),
.Y(n_5182)
);

OAI221xp5_ASAP7_75t_L g5183 ( 
.A1(n_5154),
.A2(n_5130),
.B1(n_5124),
.B2(n_5120),
.C(n_5123),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_5169),
.B(n_5133),
.Y(n_5184)
);

OAI22xp5_ASAP7_75t_L g5185 ( 
.A1(n_5163),
.A2(n_4729),
.B1(n_4737),
.B2(n_4728),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5154),
.Y(n_5186)
);

NAND2xp5_ASAP7_75t_L g5187 ( 
.A(n_5172),
.B(n_4729),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_5174),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5178),
.Y(n_5189)
);

NOR2xp33_ASAP7_75t_L g5190 ( 
.A(n_5157),
.B(n_4819),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_SL g5191 ( 
.A(n_5163),
.B(n_4681),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_5172),
.Y(n_5192)
);

INVxp67_ASAP7_75t_L g5193 ( 
.A(n_5147),
.Y(n_5193)
);

AOI221xp5_ASAP7_75t_L g5194 ( 
.A1(n_5165),
.A2(n_5155),
.B1(n_5170),
.B2(n_5173),
.C(n_5167),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_5149),
.Y(n_5195)
);

OAI221xp5_ASAP7_75t_L g5196 ( 
.A1(n_5170),
.A2(n_4675),
.B1(n_4678),
.B2(n_4670),
.C(n_4669),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_5149),
.B(n_4737),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_SL g5198 ( 
.A(n_5150),
.B(n_4681),
.Y(n_5198)
);

NAND3xp33_ASAP7_75t_L g5199 ( 
.A(n_5164),
.B(n_4601),
.C(n_4579),
.Y(n_5199)
);

NOR2xp33_ASAP7_75t_L g5200 ( 
.A(n_5166),
.B(n_4723),
.Y(n_5200)
);

NOR2xp67_ASAP7_75t_SL g5201 ( 
.A(n_5146),
.B(n_4761),
.Y(n_5201)
);

NAND2xp5_ASAP7_75t_L g5202 ( 
.A(n_5159),
.B(n_4689),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_5151),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5161),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5164),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_5156),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5162),
.Y(n_5207)
);

OAI22xp33_ASAP7_75t_L g5208 ( 
.A1(n_5177),
.A2(n_4718),
.B1(n_4715),
.B2(n_4700),
.Y(n_5208)
);

NOR2x1_ASAP7_75t_L g5209 ( 
.A(n_5153),
.B(n_4698),
.Y(n_5209)
);

INVx1_ASAP7_75t_SL g5210 ( 
.A(n_5168),
.Y(n_5210)
);

OAI22xp33_ASAP7_75t_L g5211 ( 
.A1(n_5152),
.A2(n_4701),
.B1(n_4754),
.B2(n_4577),
.Y(n_5211)
);

OAI322xp33_ASAP7_75t_L g5212 ( 
.A1(n_5176),
.A2(n_4724),
.A3(n_4730),
.B1(n_4597),
.B2(n_4582),
.C1(n_4704),
.C2(n_4828),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_5158),
.B(n_4828),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_5171),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5179),
.B(n_4731),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_5175),
.B(n_4764),
.Y(n_5216)
);

INVx2_ASAP7_75t_L g5217 ( 
.A(n_5215),
.Y(n_5217)
);

OAI221xp5_ASAP7_75t_L g5218 ( 
.A1(n_5194),
.A2(n_4646),
.B1(n_4730),
.B2(n_4724),
.C(n_4569),
.Y(n_5218)
);

OAI22xp5_ASAP7_75t_L g5219 ( 
.A1(n_5199),
.A2(n_5186),
.B1(n_5210),
.B2(n_5193),
.Y(n_5219)
);

AOI221x1_ASAP7_75t_L g5220 ( 
.A1(n_5189),
.A2(n_4712),
.B1(n_4615),
.B2(n_4766),
.C(n_4634),
.Y(n_5220)
);

OAI22xp5_ASAP7_75t_L g5221 ( 
.A1(n_5199),
.A2(n_4712),
.B1(n_4354),
.B2(n_4566),
.Y(n_5221)
);

OAI211xp5_ASAP7_75t_L g5222 ( 
.A1(n_5191),
.A2(n_4601),
.B(n_4579),
.C(n_4603),
.Y(n_5222)
);

OAI21xp33_ASAP7_75t_L g5223 ( 
.A1(n_5190),
.A2(n_4583),
.B(n_4639),
.Y(n_5223)
);

NOR2x1_ASAP7_75t_L g5224 ( 
.A(n_5180),
.B(n_4607),
.Y(n_5224)
);

INVx1_ASAP7_75t_SL g5225 ( 
.A(n_5198),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5201),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5187),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5197),
.Y(n_5228)
);

NAND2xp5_ASAP7_75t_L g5229 ( 
.A(n_5192),
.B(n_5185),
.Y(n_5229)
);

HB1xp67_ASAP7_75t_L g5230 ( 
.A(n_5213),
.Y(n_5230)
);

CKINVDCx14_ASAP7_75t_R g5231 ( 
.A(n_5203),
.Y(n_5231)
);

INVx2_ASAP7_75t_L g5232 ( 
.A(n_5195),
.Y(n_5232)
);

OAI221xp5_ASAP7_75t_L g5233 ( 
.A1(n_5183),
.A2(n_4599),
.B1(n_4611),
.B2(n_4595),
.C(n_4590),
.Y(n_5233)
);

AOI21xp33_ASAP7_75t_SL g5234 ( 
.A1(n_5182),
.A2(n_5205),
.B(n_5216),
.Y(n_5234)
);

OAI22xp33_ASAP7_75t_L g5235 ( 
.A1(n_5207),
.A2(n_4354),
.B1(n_4411),
.B2(n_4396),
.Y(n_5235)
);

AND2x2_ASAP7_75t_L g5236 ( 
.A(n_5188),
.B(n_4389),
.Y(n_5236)
);

OAI22xp5_ASAP7_75t_L g5237 ( 
.A1(n_5206),
.A2(n_4618),
.B1(n_4628),
.B2(n_4627),
.Y(n_5237)
);

OAI22xp5_ASAP7_75t_L g5238 ( 
.A1(n_5214),
.A2(n_4565),
.B1(n_4563),
.B2(n_4613),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5184),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_5202),
.Y(n_5240)
);

OAI22xp5_ASAP7_75t_L g5241 ( 
.A1(n_5204),
.A2(n_4397),
.B1(n_4433),
.B2(n_4466),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_L g5242 ( 
.A(n_5208),
.B(n_4645),
.Y(n_5242)
);

AOI22xp5_ASAP7_75t_L g5243 ( 
.A1(n_5200),
.A2(n_4379),
.B1(n_377),
.B2(n_375),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_5209),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_SL g5245 ( 
.A(n_5211),
.B(n_650),
.Y(n_5245)
);

OAI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_5196),
.A2(n_5181),
.B(n_5212),
.Y(n_5246)
);

AND2x2_ASAP7_75t_L g5247 ( 
.A(n_5212),
.B(n_376),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5201),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5201),
.Y(n_5249)
);

OAI22xp33_ASAP7_75t_L g5250 ( 
.A1(n_5199),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_5201),
.Y(n_5251)
);

OAI21xp33_ASAP7_75t_L g5252 ( 
.A1(n_5210),
.A2(n_378),
.B(n_379),
.Y(n_5252)
);

XNOR2xp5_ASAP7_75t_L g5253 ( 
.A(n_5210),
.B(n_380),
.Y(n_5253)
);

OR2x2_ASAP7_75t_L g5254 ( 
.A(n_5191),
.B(n_381),
.Y(n_5254)
);

OAI321xp33_ASAP7_75t_L g5255 ( 
.A1(n_5183),
.A2(n_381),
.A3(n_382),
.B1(n_383),
.B2(n_385),
.C(n_386),
.Y(n_5255)
);

OAI22xp5_ASAP7_75t_L g5256 ( 
.A1(n_5199),
.A2(n_387),
.B1(n_382),
.B2(n_385),
.Y(n_5256)
);

AND2x2_ASAP7_75t_L g5257 ( 
.A(n_5215),
.B(n_387),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5201),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_5201),
.Y(n_5259)
);

INVx1_ASAP7_75t_SL g5260 ( 
.A(n_5191),
.Y(n_5260)
);

INVx3_ASAP7_75t_L g5261 ( 
.A(n_5192),
.Y(n_5261)
);

AND2x2_ASAP7_75t_L g5262 ( 
.A(n_5215),
.B(n_388),
.Y(n_5262)
);

AND2x2_ASAP7_75t_L g5263 ( 
.A(n_5261),
.B(n_389),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5253),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_5257),
.Y(n_5265)
);

NOR2xp33_ASAP7_75t_L g5266 ( 
.A(n_5261),
.B(n_389),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_5262),
.B(n_390),
.Y(n_5267)
);

AOI22xp33_ASAP7_75t_SL g5268 ( 
.A1(n_5231),
.A2(n_5218),
.B1(n_5248),
.B2(n_5226),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_5224),
.B(n_5247),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_5224),
.B(n_390),
.Y(n_5270)
);

AOI22xp5_ASAP7_75t_L g5271 ( 
.A1(n_5260),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_5271)
);

AOI22xp33_ASAP7_75t_L g5272 ( 
.A1(n_5249),
.A2(n_395),
.B1(n_391),
.B2(n_394),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_SL g5273 ( 
.A(n_5251),
.B(n_394),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_5223),
.B(n_396),
.Y(n_5274)
);

NOR2xp33_ASAP7_75t_L g5275 ( 
.A(n_5255),
.B(n_5258),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_5259),
.B(n_396),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_5219),
.Y(n_5277)
);

BUFx2_ASAP7_75t_L g5278 ( 
.A(n_5244),
.Y(n_5278)
);

AOI22xp5_ASAP7_75t_L g5279 ( 
.A1(n_5225),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_5254),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_5242),
.Y(n_5281)
);

HB1xp67_ASAP7_75t_L g5282 ( 
.A(n_5256),
.Y(n_5282)
);

OAI22xp5_ASAP7_75t_L g5283 ( 
.A1(n_5233),
.A2(n_401),
.B1(n_398),
.B2(n_399),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5229),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5217),
.Y(n_5285)
);

NOR2x1_ASAP7_75t_L g5286 ( 
.A(n_5246),
.B(n_401),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_5250),
.B(n_402),
.Y(n_5287)
);

INVx2_ASAP7_75t_L g5288 ( 
.A(n_5232),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5236),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_5230),
.Y(n_5290)
);

NAND2xp33_ASAP7_75t_SL g5291 ( 
.A(n_5245),
.B(n_403),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_5239),
.B(n_404),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5252),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5227),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5228),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5221),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_5222),
.B(n_404),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_5234),
.A2(n_405),
.B(n_406),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_5240),
.Y(n_5299)
);

INVx2_ASAP7_75t_SL g5300 ( 
.A(n_5241),
.Y(n_5300)
);

AND2x2_ASAP7_75t_L g5301 ( 
.A(n_5238),
.B(n_405),
.Y(n_5301)
);

NOR2xp33_ASAP7_75t_L g5302 ( 
.A(n_5237),
.B(n_406),
.Y(n_5302)
);

HB1xp67_ASAP7_75t_L g5303 ( 
.A(n_5243),
.Y(n_5303)
);

OR2x2_ASAP7_75t_L g5304 ( 
.A(n_5235),
.B(n_407),
.Y(n_5304)
);

INVx1_ASAP7_75t_SL g5305 ( 
.A(n_5220),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5257),
.B(n_407),
.Y(n_5306)
);

AND2x2_ASAP7_75t_L g5307 ( 
.A(n_5261),
.B(n_408),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_5261),
.B(n_408),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_L g5309 ( 
.A(n_5257),
.B(n_409),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5253),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_L g5311 ( 
.A(n_5257),
.B(n_410),
.Y(n_5311)
);

OR2x2_ASAP7_75t_L g5312 ( 
.A(n_5221),
.B(n_410),
.Y(n_5312)
);

NOR2xp33_ASAP7_75t_L g5313 ( 
.A(n_5261),
.B(n_411),
.Y(n_5313)
);

INVx1_ASAP7_75t_SL g5314 ( 
.A(n_5257),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5257),
.B(n_412),
.Y(n_5315)
);

OR2x2_ASAP7_75t_L g5316 ( 
.A(n_5221),
.B(n_413),
.Y(n_5316)
);

NAND2xp5_ASAP7_75t_L g5317 ( 
.A(n_5257),
.B(n_413),
.Y(n_5317)
);

OAI22xp5_ASAP7_75t_L g5318 ( 
.A1(n_5218),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5253),
.Y(n_5319)
);

AOI311xp33_ASAP7_75t_L g5320 ( 
.A1(n_5298),
.A2(n_414),
.A3(n_416),
.B(n_417),
.C(n_418),
.Y(n_5320)
);

INVxp67_ASAP7_75t_L g5321 ( 
.A(n_5266),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_SL g5322 ( 
.A(n_5305),
.B(n_417),
.Y(n_5322)
);

AOI22xp5_ASAP7_75t_L g5323 ( 
.A1(n_5277),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_5263),
.B(n_419),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_5307),
.B(n_420),
.Y(n_5325)
);

INVx1_ASAP7_75t_SL g5326 ( 
.A(n_5305),
.Y(n_5326)
);

NOR3xp33_ASAP7_75t_SL g5327 ( 
.A(n_5291),
.B(n_421),
.C(n_422),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_5308),
.B(n_421),
.Y(n_5328)
);

NOR2x1p5_ASAP7_75t_L g5329 ( 
.A(n_5297),
.B(n_422),
.Y(n_5329)
);

NOR2xp33_ASAP7_75t_L g5330 ( 
.A(n_5314),
.B(n_423),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_5292),
.B(n_424),
.Y(n_5331)
);

AOI321xp33_ASAP7_75t_L g5332 ( 
.A1(n_5286),
.A2(n_5275),
.A3(n_5285),
.B1(n_5296),
.B2(n_5284),
.C(n_5269),
.Y(n_5332)
);

AOI222xp33_ASAP7_75t_L g5333 ( 
.A1(n_5278),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.C1(n_427),
.C2(n_428),
.Y(n_5333)
);

INVx4_ASAP7_75t_L g5334 ( 
.A(n_5290),
.Y(n_5334)
);

INVx1_ASAP7_75t_SL g5335 ( 
.A(n_5270),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_5313),
.B(n_427),
.Y(n_5336)
);

A2O1A1Ixp33_ASAP7_75t_L g5337 ( 
.A1(n_5302),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5267),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_5314),
.B(n_429),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5306),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_5265),
.B(n_430),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5279),
.B(n_431),
.Y(n_5342)
);

INVxp67_ASAP7_75t_L g5343 ( 
.A(n_5309),
.Y(n_5343)
);

OAI21xp5_ASAP7_75t_L g5344 ( 
.A1(n_5268),
.A2(n_432),
.B(n_433),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_5271),
.B(n_432),
.Y(n_5345)
);

XNOR2xp5_ASAP7_75t_L g5346 ( 
.A(n_5283),
.B(n_434),
.Y(n_5346)
);

OAI21x1_ASAP7_75t_L g5347 ( 
.A1(n_5318),
.A2(n_435),
.B(n_436),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5311),
.Y(n_5348)
);

NAND2xp5_ASAP7_75t_L g5349 ( 
.A(n_5288),
.B(n_435),
.Y(n_5349)
);

AOI21xp33_ASAP7_75t_L g5350 ( 
.A1(n_5312),
.A2(n_437),
.B(n_438),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_5316),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5315),
.Y(n_5352)
);

NAND2xp5_ASAP7_75t_L g5353 ( 
.A(n_5272),
.B(n_5317),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_5301),
.B(n_437),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5276),
.Y(n_5355)
);

NOR2x1_ASAP7_75t_L g5356 ( 
.A(n_5273),
.B(n_5289),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5274),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5304),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_5287),
.Y(n_5359)
);

NOR2x1_ASAP7_75t_L g5360 ( 
.A(n_5280),
.B(n_439),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5282),
.Y(n_5361)
);

INVxp67_ASAP7_75t_SL g5362 ( 
.A(n_5303),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5294),
.Y(n_5363)
);

OR2x2_ASAP7_75t_L g5364 ( 
.A(n_5264),
.B(n_439),
.Y(n_5364)
);

AOI22x1_ASAP7_75t_L g5365 ( 
.A1(n_5334),
.A2(n_5300),
.B1(n_5295),
.B2(n_5299),
.Y(n_5365)
);

NOR3xp33_ASAP7_75t_L g5366 ( 
.A(n_5334),
.B(n_5319),
.C(n_5310),
.Y(n_5366)
);

AO22x2_ASAP7_75t_L g5367 ( 
.A1(n_5326),
.A2(n_5281),
.B1(n_5293),
.B2(n_442),
.Y(n_5367)
);

AO21x1_ASAP7_75t_L g5368 ( 
.A1(n_5322),
.A2(n_440),
.B(n_441),
.Y(n_5368)
);

NOR4xp25_ASAP7_75t_L g5369 ( 
.A(n_5344),
.B(n_443),
.C(n_440),
.D(n_442),
.Y(n_5369)
);

AOI211xp5_ASAP7_75t_L g5370 ( 
.A1(n_5350),
.A2(n_446),
.B(n_443),
.C(n_445),
.Y(n_5370)
);

AND2x2_ASAP7_75t_L g5371 ( 
.A(n_5362),
.B(n_5320),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_5360),
.Y(n_5372)
);

AOI21xp5_ASAP7_75t_L g5373 ( 
.A1(n_5339),
.A2(n_445),
.B(n_446),
.Y(n_5373)
);

NOR3xp33_ASAP7_75t_L g5374 ( 
.A(n_5361),
.B(n_447),
.C(n_448),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_SL g5375 ( 
.A(n_5332),
.B(n_448),
.Y(n_5375)
);

NOR2xp67_ASAP7_75t_L g5376 ( 
.A(n_5341),
.B(n_5330),
.Y(n_5376)
);

OAI21xp5_ASAP7_75t_L g5377 ( 
.A1(n_5356),
.A2(n_5346),
.B(n_5363),
.Y(n_5377)
);

AOI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_5335),
.A2(n_454),
.B1(n_450),
.B2(n_451),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5349),
.Y(n_5379)
);

NOR2xp67_ASAP7_75t_L g5380 ( 
.A(n_5323),
.B(n_451),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5364),
.Y(n_5381)
);

AOI21xp5_ASAP7_75t_L g5382 ( 
.A1(n_5354),
.A2(n_454),
.B(n_455),
.Y(n_5382)
);

OAI211xp5_ASAP7_75t_SL g5383 ( 
.A1(n_5327),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_5383)
);

OAI22xp5_ASAP7_75t_L g5384 ( 
.A1(n_5324),
.A2(n_459),
.B1(n_456),
.B2(n_458),
.Y(n_5384)
);

NAND3xp33_ASAP7_75t_L g5385 ( 
.A(n_5333),
.B(n_458),
.C(n_459),
.Y(n_5385)
);

AOI22x1_ASAP7_75t_L g5386 ( 
.A1(n_5329),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_5386)
);

NOR3x1_ASAP7_75t_L g5387 ( 
.A(n_5325),
.B(n_460),
.C(n_462),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_SL g5388 ( 
.A(n_5328),
.B(n_463),
.Y(n_5388)
);

AOI21xp5_ASAP7_75t_L g5389 ( 
.A1(n_5336),
.A2(n_464),
.B(n_465),
.Y(n_5389)
);

AND2x2_ASAP7_75t_L g5390 ( 
.A(n_5351),
.B(n_464),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_5337),
.B(n_465),
.Y(n_5391)
);

AOI211xp5_ASAP7_75t_L g5392 ( 
.A1(n_5342),
.A2(n_466),
.B(n_467),
.C(n_468),
.Y(n_5392)
);

AOI22xp5_ASAP7_75t_L g5393 ( 
.A1(n_5358),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.Y(n_5393)
);

NOR2x1_ASAP7_75t_L g5394 ( 
.A(n_5331),
.B(n_469),
.Y(n_5394)
);

NOR3x1_ASAP7_75t_L g5395 ( 
.A(n_5345),
.B(n_470),
.C(n_471),
.Y(n_5395)
);

HB1xp67_ASAP7_75t_L g5396 ( 
.A(n_5347),
.Y(n_5396)
);

AOI211xp5_ASAP7_75t_L g5397 ( 
.A1(n_5321),
.A2(n_470),
.B(n_471),
.C(n_472),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5353),
.Y(n_5398)
);

OAI22xp5_ASAP7_75t_L g5399 ( 
.A1(n_5343),
.A2(n_472),
.B1(n_473),
.B2(n_475),
.Y(n_5399)
);

AO22x1_ASAP7_75t_L g5400 ( 
.A1(n_5357),
.A2(n_473),
.B1(n_475),
.B2(n_476),
.Y(n_5400)
);

NAND2xp5_ASAP7_75t_L g5401 ( 
.A(n_5338),
.B(n_476),
.Y(n_5401)
);

NOR3x1_ASAP7_75t_L g5402 ( 
.A(n_5359),
.B(n_477),
.C(n_478),
.Y(n_5402)
);

AO22x2_ASAP7_75t_L g5403 ( 
.A1(n_5340),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_5403)
);

BUFx2_ASAP7_75t_L g5404 ( 
.A(n_5367),
.Y(n_5404)
);

OAI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_5385),
.A2(n_5375),
.B(n_5366),
.Y(n_5405)
);

AOI21xp5_ASAP7_75t_L g5406 ( 
.A1(n_5396),
.A2(n_5372),
.B(n_5388),
.Y(n_5406)
);

AOI21xp5_ASAP7_75t_L g5407 ( 
.A1(n_5377),
.A2(n_5352),
.B(n_5348),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_5365),
.Y(n_5408)
);

AOI22xp5_ASAP7_75t_L g5409 ( 
.A1(n_5371),
.A2(n_5355),
.B1(n_481),
.B2(n_483),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5367),
.Y(n_5410)
);

AOI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5369),
.A2(n_480),
.B1(n_481),
.B2(n_484),
.C(n_485),
.Y(n_5411)
);

AOI211xp5_ASAP7_75t_L g5412 ( 
.A1(n_5368),
.A2(n_485),
.B(n_486),
.C(n_487),
.Y(n_5412)
);

AOI21xp33_ASAP7_75t_L g5413 ( 
.A1(n_5394),
.A2(n_5398),
.B(n_5391),
.Y(n_5413)
);

AOI211xp5_ASAP7_75t_SL g5414 ( 
.A1(n_5376),
.A2(n_486),
.B(n_487),
.C(n_488),
.Y(n_5414)
);

AOI322xp5_ASAP7_75t_L g5415 ( 
.A1(n_5381),
.A2(n_488),
.A3(n_489),
.B1(n_490),
.B2(n_491),
.C1(n_492),
.C2(n_494),
.Y(n_5415)
);

AOI21xp33_ASAP7_75t_L g5416 ( 
.A1(n_5383),
.A2(n_489),
.B(n_491),
.Y(n_5416)
);

NOR2xp67_ASAP7_75t_L g5417 ( 
.A(n_5382),
.B(n_492),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5402),
.Y(n_5418)
);

OAI31xp33_ASAP7_75t_L g5419 ( 
.A1(n_5379),
.A2(n_650),
.A3(n_495),
.B(n_496),
.Y(n_5419)
);

O2A1O1Ixp33_ASAP7_75t_L g5420 ( 
.A1(n_5373),
.A2(n_494),
.B(n_495),
.C(n_497),
.Y(n_5420)
);

OAI221xp5_ASAP7_75t_SL g5421 ( 
.A1(n_5370),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.C(n_500),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5401),
.Y(n_5422)
);

AOI322xp5_ASAP7_75t_L g5423 ( 
.A1(n_5374),
.A2(n_5390),
.A3(n_5378),
.B1(n_5393),
.B2(n_5395),
.C1(n_5380),
.C2(n_5387),
.Y(n_5423)
);

OAI221xp5_ASAP7_75t_L g5424 ( 
.A1(n_5386),
.A2(n_498),
.B1(n_499),
.B2(n_501),
.C(n_502),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_L g5425 ( 
.A(n_5397),
.B(n_502),
.Y(n_5425)
);

AOI21xp33_ASAP7_75t_L g5426 ( 
.A1(n_5392),
.A2(n_503),
.B(n_504),
.Y(n_5426)
);

O2A1O1Ixp33_ASAP7_75t_SL g5427 ( 
.A1(n_5389),
.A2(n_503),
.B(n_504),
.C(n_505),
.Y(n_5427)
);

INVx2_ASAP7_75t_L g5428 ( 
.A(n_5403),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5403),
.Y(n_5429)
);

OAI221xp5_ASAP7_75t_L g5430 ( 
.A1(n_5384),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.C(n_508),
.Y(n_5430)
);

AOI22xp5_ASAP7_75t_L g5431 ( 
.A1(n_5399),
.A2(n_649),
.B1(n_508),
.B2(n_509),
.Y(n_5431)
);

OAI21xp33_ASAP7_75t_SL g5432 ( 
.A1(n_5400),
.A2(n_507),
.B(n_511),
.Y(n_5432)
);

OAI21xp5_ASAP7_75t_L g5433 ( 
.A1(n_5385),
.A2(n_511),
.B(n_512),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_5367),
.Y(n_5434)
);

OAI21xp33_ASAP7_75t_SL g5435 ( 
.A1(n_5429),
.A2(n_513),
.B(n_514),
.Y(n_5435)
);

AOI221xp5_ASAP7_75t_L g5436 ( 
.A1(n_5416),
.A2(n_513),
.B1(n_515),
.B2(n_516),
.C(n_517),
.Y(n_5436)
);

NAND2xp5_ASAP7_75t_L g5437 ( 
.A(n_5414),
.B(n_517),
.Y(n_5437)
);

O2A1O1Ixp5_ASAP7_75t_L g5438 ( 
.A1(n_5433),
.A2(n_518),
.B(n_519),
.C(n_520),
.Y(n_5438)
);

AOI211xp5_ASAP7_75t_SL g5439 ( 
.A1(n_5413),
.A2(n_518),
.B(n_520),
.C(n_521),
.Y(n_5439)
);

AOI221xp5_ASAP7_75t_L g5440 ( 
.A1(n_5426),
.A2(n_521),
.B1(n_522),
.B2(n_523),
.C(n_524),
.Y(n_5440)
);

AOI221xp5_ASAP7_75t_SL g5441 ( 
.A1(n_5406),
.A2(n_522),
.B1(n_524),
.B2(n_525),
.C(n_526),
.Y(n_5441)
);

OAI211xp5_ASAP7_75t_SL g5442 ( 
.A1(n_5423),
.A2(n_526),
.B(n_527),
.C(n_529),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_L g5443 ( 
.A(n_5411),
.B(n_530),
.Y(n_5443)
);

NAND4xp25_ASAP7_75t_L g5444 ( 
.A(n_5409),
.B(n_530),
.C(n_531),
.D(n_532),
.Y(n_5444)
);

NAND4xp75_ASAP7_75t_L g5445 ( 
.A(n_5405),
.B(n_531),
.C(n_533),
.D(n_534),
.Y(n_5445)
);

NOR3xp33_ASAP7_75t_L g5446 ( 
.A(n_5418),
.B(n_649),
.C(n_534),
.Y(n_5446)
);

AOI221xp5_ASAP7_75t_L g5447 ( 
.A1(n_5427),
.A2(n_533),
.B1(n_535),
.B2(n_536),
.C(n_537),
.Y(n_5447)
);

O2A1O1Ixp5_ASAP7_75t_L g5448 ( 
.A1(n_5428),
.A2(n_538),
.B(n_539),
.C(n_540),
.Y(n_5448)
);

A2O1A1Ixp33_ASAP7_75t_L g5449 ( 
.A1(n_5420),
.A2(n_538),
.B(n_541),
.C(n_542),
.Y(n_5449)
);

NAND2xp5_ASAP7_75t_L g5450 ( 
.A(n_5412),
.B(n_541),
.Y(n_5450)
);

NOR2xp67_ASAP7_75t_SL g5451 ( 
.A(n_5408),
.B(n_5410),
.Y(n_5451)
);

OAI21xp5_ASAP7_75t_SL g5452 ( 
.A1(n_5431),
.A2(n_648),
.B(n_543),
.Y(n_5452)
);

INVx1_ASAP7_75t_SL g5453 ( 
.A(n_5404),
.Y(n_5453)
);

NAND4xp25_ASAP7_75t_L g5454 ( 
.A(n_5407),
.B(n_542),
.C(n_543),
.D(n_544),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_5425),
.Y(n_5455)
);

HB1xp67_ASAP7_75t_L g5456 ( 
.A(n_5432),
.Y(n_5456)
);

NAND4xp25_ASAP7_75t_L g5457 ( 
.A(n_5421),
.B(n_544),
.C(n_545),
.D(n_546),
.Y(n_5457)
);

OAI221xp5_ASAP7_75t_L g5458 ( 
.A1(n_5424),
.A2(n_545),
.B1(n_546),
.B2(n_548),
.C(n_549),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5417),
.B(n_548),
.Y(n_5459)
);

NAND3xp33_ASAP7_75t_L g5460 ( 
.A(n_5419),
.B(n_549),
.C(n_550),
.Y(n_5460)
);

NOR2x1p5_ASAP7_75t_L g5461 ( 
.A(n_5434),
.B(n_550),
.Y(n_5461)
);

OAI21xp33_ASAP7_75t_SL g5462 ( 
.A1(n_5422),
.A2(n_551),
.B(n_552),
.Y(n_5462)
);

AOI21xp33_ASAP7_75t_L g5463 ( 
.A1(n_5430),
.A2(n_553),
.B(n_554),
.Y(n_5463)
);

NAND2xp5_ASAP7_75t_L g5464 ( 
.A(n_5461),
.B(n_5415),
.Y(n_5464)
);

NAND4xp25_ASAP7_75t_L g5465 ( 
.A(n_5436),
.B(n_553),
.C(n_554),
.D(n_555),
.Y(n_5465)
);

NAND2x1p5_ASAP7_75t_L g5466 ( 
.A(n_5453),
.B(n_556),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5437),
.Y(n_5467)
);

AND2x2_ASAP7_75t_L g5468 ( 
.A(n_5459),
.B(n_557),
.Y(n_5468)
);

NOR3xp33_ASAP7_75t_L g5469 ( 
.A(n_5456),
.B(n_648),
.C(n_558),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_5445),
.Y(n_5470)
);

AND2x4_ASAP7_75t_L g5471 ( 
.A(n_5460),
.B(n_557),
.Y(n_5471)
);

BUFx8_ASAP7_75t_SL g5472 ( 
.A(n_5455),
.Y(n_5472)
);

NOR3xp33_ASAP7_75t_L g5473 ( 
.A(n_5463),
.B(n_5458),
.C(n_5457),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5435),
.Y(n_5474)
);

NOR2xp33_ASAP7_75t_L g5475 ( 
.A(n_5444),
.B(n_559),
.Y(n_5475)
);

NOR3x1_ASAP7_75t_L g5476 ( 
.A(n_5452),
.B(n_647),
.C(n_561),
.Y(n_5476)
);

AND2x2_ASAP7_75t_L g5477 ( 
.A(n_5439),
.B(n_560),
.Y(n_5477)
);

XNOR2xp5_ASAP7_75t_L g5478 ( 
.A(n_5454),
.B(n_560),
.Y(n_5478)
);

NOR3xp33_ASAP7_75t_L g5479 ( 
.A(n_5450),
.B(n_562),
.C(n_563),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5438),
.Y(n_5480)
);

NOR2x1_ASAP7_75t_L g5481 ( 
.A(n_5442),
.B(n_562),
.Y(n_5481)
);

NOR2x1_ASAP7_75t_L g5482 ( 
.A(n_5449),
.B(n_565),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_5462),
.Y(n_5483)
);

NAND3x1_ASAP7_75t_L g5484 ( 
.A(n_5446),
.B(n_565),
.C(n_566),
.Y(n_5484)
);

NOR3xp33_ASAP7_75t_L g5485 ( 
.A(n_5440),
.B(n_646),
.C(n_567),
.Y(n_5485)
);

NAND4xp75_ASAP7_75t_L g5486 ( 
.A(n_5441),
.B(n_566),
.C(n_567),
.D(n_568),
.Y(n_5486)
);

NOR2x1_ASAP7_75t_L g5487 ( 
.A(n_5443),
.B(n_568),
.Y(n_5487)
);

NAND4xp75_ASAP7_75t_L g5488 ( 
.A(n_5447),
.B(n_569),
.C(n_570),
.D(n_572),
.Y(n_5488)
);

NOR2x1_ASAP7_75t_L g5489 ( 
.A(n_5448),
.B(n_569),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5451),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5461),
.Y(n_5491)
);

AND4x1_ASAP7_75t_L g5492 ( 
.A(n_5490),
.B(n_646),
.C(n_572),
.D(n_573),
.Y(n_5492)
);

AOI221xp5_ASAP7_75t_L g5493 ( 
.A1(n_5475),
.A2(n_570),
.B1(n_573),
.B2(n_574),
.C(n_575),
.Y(n_5493)
);

AND3x2_ASAP7_75t_L g5494 ( 
.A(n_5474),
.B(n_574),
.C(n_576),
.Y(n_5494)
);

NAND2xp5_ASAP7_75t_L g5495 ( 
.A(n_5468),
.B(n_576),
.Y(n_5495)
);

NOR4xp25_ASAP7_75t_L g5496 ( 
.A(n_5483),
.B(n_5480),
.C(n_5470),
.D(n_5491),
.Y(n_5496)
);

NAND4xp75_ASAP7_75t_L g5497 ( 
.A(n_5487),
.B(n_577),
.C(n_578),
.D(n_579),
.Y(n_5497)
);

AOI221x1_ASAP7_75t_SL g5498 ( 
.A1(n_5471),
.A2(n_577),
.B1(n_579),
.B2(n_580),
.C(n_581),
.Y(n_5498)
);

INVxp67_ASAP7_75t_L g5499 ( 
.A(n_5466),
.Y(n_5499)
);

NAND3xp33_ASAP7_75t_SL g5500 ( 
.A(n_5469),
.B(n_580),
.C(n_581),
.Y(n_5500)
);

OAI221xp5_ASAP7_75t_L g5501 ( 
.A1(n_5479),
.A2(n_582),
.B1(n_583),
.B2(n_584),
.C(n_585),
.Y(n_5501)
);

NAND4xp25_ASAP7_75t_SL g5502 ( 
.A(n_5481),
.B(n_5485),
.C(n_5489),
.D(n_5473),
.Y(n_5502)
);

NAND2xp5_ASAP7_75t_SL g5503 ( 
.A(n_5471),
.B(n_582),
.Y(n_5503)
);

NAND3xp33_ASAP7_75t_SL g5504 ( 
.A(n_5464),
.B(n_586),
.C(n_587),
.Y(n_5504)
);

NOR3xp33_ASAP7_75t_L g5505 ( 
.A(n_5467),
.B(n_586),
.C(n_588),
.Y(n_5505)
);

NAND4xp25_ASAP7_75t_L g5506 ( 
.A(n_5476),
.B(n_588),
.C(n_589),
.D(n_590),
.Y(n_5506)
);

NAND5xp2_ASAP7_75t_L g5507 ( 
.A(n_5477),
.B(n_589),
.C(n_591),
.D(n_592),
.E(n_593),
.Y(n_5507)
);

NAND3x2_ASAP7_75t_L g5508 ( 
.A(n_5484),
.B(n_593),
.C(n_594),
.Y(n_5508)
);

OAI21xp33_ASAP7_75t_L g5509 ( 
.A1(n_5465),
.A2(n_594),
.B(n_595),
.Y(n_5509)
);

AOI211xp5_ASAP7_75t_SL g5510 ( 
.A1(n_5472),
.A2(n_595),
.B(n_596),
.C(n_597),
.Y(n_5510)
);

NAND4xp75_ASAP7_75t_L g5511 ( 
.A(n_5482),
.B(n_5478),
.C(n_5488),
.D(n_5486),
.Y(n_5511)
);

NOR4xp25_ASAP7_75t_L g5512 ( 
.A(n_5490),
.B(n_597),
.C(n_598),
.D(n_599),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5494),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_L g5514 ( 
.A(n_5507),
.B(n_599),
.Y(n_5514)
);

AOI22xp5_ASAP7_75t_L g5515 ( 
.A1(n_5504),
.A2(n_5509),
.B1(n_5502),
.B2(n_5506),
.Y(n_5515)
);

NAND2xp5_ASAP7_75t_L g5516 ( 
.A(n_5498),
.B(n_5495),
.Y(n_5516)
);

XNOR2xp5_ASAP7_75t_L g5517 ( 
.A(n_5508),
.B(n_600),
.Y(n_5517)
);

NOR2x1_ASAP7_75t_L g5518 ( 
.A(n_5497),
.B(n_600),
.Y(n_5518)
);

INVx2_ASAP7_75t_L g5519 ( 
.A(n_5511),
.Y(n_5519)
);

NOR2x1_ASAP7_75t_L g5520 ( 
.A(n_5500),
.B(n_601),
.Y(n_5520)
);

OAI22xp5_ASAP7_75t_SL g5521 ( 
.A1(n_5499),
.A2(n_601),
.B1(n_602),
.B2(n_603),
.Y(n_5521)
);

NOR3xp33_ASAP7_75t_L g5522 ( 
.A(n_5503),
.B(n_603),
.C(n_604),
.Y(n_5522)
);

AND2x4_ASAP7_75t_L g5523 ( 
.A(n_5505),
.B(n_605),
.Y(n_5523)
);

NOR2xp33_ASAP7_75t_L g5524 ( 
.A(n_5501),
.B(n_605),
.Y(n_5524)
);

NOR3xp33_ASAP7_75t_L g5525 ( 
.A(n_5513),
.B(n_5496),
.C(n_5493),
.Y(n_5525)
);

NOR3xp33_ASAP7_75t_L g5526 ( 
.A(n_5519),
.B(n_5512),
.C(n_5510),
.Y(n_5526)
);

AOI211xp5_ASAP7_75t_L g5527 ( 
.A1(n_5522),
.A2(n_5492),
.B(n_607),
.C(n_609),
.Y(n_5527)
);

NOR2xp33_ASAP7_75t_L g5528 ( 
.A(n_5514),
.B(n_606),
.Y(n_5528)
);

OAI21xp33_ASAP7_75t_L g5529 ( 
.A1(n_5515),
.A2(n_606),
.B(n_607),
.Y(n_5529)
);

AOI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_5517),
.A2(n_610),
.B1(n_611),
.B2(n_612),
.Y(n_5530)
);

AOI221xp5_ASAP7_75t_SL g5531 ( 
.A1(n_5528),
.A2(n_5524),
.B1(n_5516),
.B2(n_5521),
.C(n_5518),
.Y(n_5531)
);

NAND3xp33_ASAP7_75t_SL g5532 ( 
.A(n_5526),
.B(n_5520),
.C(n_5523),
.Y(n_5532)
);

A2O1A1Ixp33_ASAP7_75t_L g5533 ( 
.A1(n_5527),
.A2(n_5523),
.B(n_611),
.C(n_612),
.Y(n_5533)
);

AOI22xp5_ASAP7_75t_L g5534 ( 
.A1(n_5532),
.A2(n_5525),
.B1(n_5530),
.B2(n_5529),
.Y(n_5534)
);

XOR2x2_ASAP7_75t_L g5535 ( 
.A(n_5531),
.B(n_610),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_5535),
.Y(n_5536)
);

AOI22xp5_ASAP7_75t_L g5537 ( 
.A1(n_5536),
.A2(n_5534),
.B1(n_5533),
.B2(n_615),
.Y(n_5537)
);

OAI322xp33_ASAP7_75t_L g5538 ( 
.A1(n_5537),
.A2(n_613),
.A3(n_614),
.B1(n_615),
.B2(n_616),
.C1(n_617),
.C2(n_618),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_5538),
.Y(n_5539)
);

XOR2x2_ASAP7_75t_L g5540 ( 
.A(n_5539),
.B(n_613),
.Y(n_5540)
);

OAI221xp5_ASAP7_75t_L g5541 ( 
.A1(n_5540),
.A2(n_617),
.B1(n_618),
.B2(n_619),
.C(n_620),
.Y(n_5541)
);

OAI21xp5_ASAP7_75t_L g5542 ( 
.A1(n_5541),
.A2(n_621),
.B(n_622),
.Y(n_5542)
);

XNOR2xp5_ASAP7_75t_L g5543 ( 
.A(n_5542),
.B(n_645),
.Y(n_5543)
);

OAI21xp5_ASAP7_75t_L g5544 ( 
.A1(n_5543),
.A2(n_623),
.B(n_624),
.Y(n_5544)
);

BUFx2_ASAP7_75t_L g5545 ( 
.A(n_5544),
.Y(n_5545)
);

AOI21xp5_ASAP7_75t_L g5546 ( 
.A1(n_5545),
.A2(n_623),
.B(n_624),
.Y(n_5546)
);

OAI221xp5_ASAP7_75t_L g5547 ( 
.A1(n_5546),
.A2(n_626),
.B1(n_627),
.B2(n_628),
.C(n_629),
.Y(n_5547)
);

AOI221xp5_ASAP7_75t_L g5548 ( 
.A1(n_5546),
.A2(n_627),
.B1(n_628),
.B2(n_629),
.C(n_630),
.Y(n_5548)
);

AOI22xp33_ASAP7_75t_L g5549 ( 
.A1(n_5547),
.A2(n_631),
.B1(n_632),
.B2(n_633),
.Y(n_5549)
);

AOI211xp5_ASAP7_75t_L g5550 ( 
.A1(n_5549),
.A2(n_5548),
.B(n_632),
.C(n_633),
.Y(n_5550)
);


endmodule