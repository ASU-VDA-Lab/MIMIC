module real_jpeg_23231_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_50),
.B1(n_52),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_57),
.B1(n_73),
.B2(n_87),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_2),
.A2(n_22),
.B1(n_28),
.B2(n_73),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_39),
.B1(n_50),
.B2(n_52),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_6),
.A2(n_22),
.B1(n_28),
.B2(n_39),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_7),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_69)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_9),
.B1(n_42),
.B2(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_42),
.B1(n_50),
.B2(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_22),
.B1(n_28),
.B2(n_42),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_9),
.B(n_49),
.C(n_52),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_48),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_37),
.C(n_76),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_22),
.C(n_34),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_11),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_9),
.B(n_67),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_9),
.B(n_79),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_120),
.B1(n_259),
.B2(n_260),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_119),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_101),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_16),
.B(n_101),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_62),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_30),
.B(n_45),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_18),
.A2(n_45),
.B1(n_46),
.B2(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_18),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_18),
.A2(n_31),
.B1(n_104),
.B2(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_27),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_20),
.B(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_21),
.A2(n_27),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_21),
.B(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_21),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_22),
.B(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_30),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_31),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B(n_40),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_32),
.B(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_32),
.A2(n_40),
.B(n_137),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

OA22x2_ASAP7_75t_SL g78 ( 
.A1(n_36),
.A2(n_37),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_37),
.B(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_41),
.A2(n_43),
.B1(n_67),
.B2(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_41),
.B(n_94),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_43),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_58),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_48),
.A2(n_54),
.B1(n_59),
.B2(n_116),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_52),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_52),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_59),
.Y(n_88)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_61),
.B(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_81),
.B2(n_82),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_65),
.B(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_70),
.A2(n_115),
.B1(n_125),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_177),
.C(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_70),
.A2(n_167),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_70),
.B(n_115),
.C(n_157),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_78),
.B(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_97),
.B(n_99),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_80),
.Y(n_140)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_117),
.C(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_83),
.A2(n_84),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_83),
.A2(n_84),
.B1(n_138),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_129),
.C(n_138),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_100),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_106),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_105),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_115),
.C(n_117),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_108),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_112),
.A2(n_113),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_112),
.A2(n_113),
.B1(n_190),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_184),
.C(n_190),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_113),
.B(n_162),
.C(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_117),
.A2(n_118),
.B1(n_153),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_117),
.A2(n_118),
.B1(n_136),
.B2(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_118),
.B(n_136),
.C(n_228),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_120),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_143),
.B(n_258),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_141),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_122),
.B(n_141),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_126),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_128),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_129),
.A2(n_130),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_136),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_164),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_136),
.A2(n_150),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_253),
.B(n_257),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_180),
.B(n_239),
.C(n_252),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_169),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_146),
.B(n_169),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_156),
.B2(n_168),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_149),
.B(n_155),
.C(n_168),
.Y(n_240)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_166),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_161),
.A2(n_162),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_213),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.C(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_171),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_176),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_179),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_177),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_238),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_199),
.B(n_237),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_183),
.B(n_196),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_185),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_230),
.B(n_236),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_224),
.B(n_229),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_216),
.B(n_223),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_208),
.B(n_215),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_205),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_212),
.B(n_214),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_241),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_251),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_249),
.C(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);


endmodule