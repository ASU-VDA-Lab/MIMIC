module fake_jpeg_1364_n_224 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_224);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_20),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_2),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_88),
.B(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_59),
.B1(n_58),
.B2(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_70),
.B1(n_68),
.B2(n_73),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_65),
.CON(n_94),
.SN(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx6f_ASAP7_75t_SL g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_100),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_95),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_92),
.B1(n_98),
.B2(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_111),
.B1(n_113),
.B2(n_117),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_109),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_106),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_66),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_63),
.C(n_74),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_78),
.C(n_61),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_59),
.B1(n_99),
.B2(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_63),
.B1(n_74),
.B2(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_64),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_79),
.B1(n_56),
.B2(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_61),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_4),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_128),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_67),
.C(n_72),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_129),
.C(n_130),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_71),
.C(n_62),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_57),
.C(n_60),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_136),
.Y(n_148)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_1),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_95),
.C(n_55),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_3),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_3),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_95),
.C(n_55),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_150),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_116),
.B(n_107),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_116),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_10),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_75),
.C(n_60),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_100),
.B1(n_75),
.B2(n_60),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_158),
.B1(n_161),
.B2(n_33),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_25),
.B1(n_51),
.B2(n_50),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_156),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_157),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_141),
.B1(n_132),
.B2(n_120),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_23),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_6),
.C(n_7),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_160),
.B(n_9),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_7),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_169),
.B(n_182),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_8),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_177),
.B1(n_151),
.B2(n_159),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_12),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_34),
.C(n_49),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_181),
.C(n_165),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_30),
.C(n_48),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_11),
.Y(n_182)
);

OAI22x1_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_27),
.B1(n_47),
.B2(n_44),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_26),
.B1(n_43),
.B2(n_40),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_188),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_162),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_149),
.B1(n_145),
.B2(n_147),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_196),
.B1(n_170),
.B2(n_175),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_13),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_53),
.B1(n_39),
.B2(n_38),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_168),
.B1(n_37),
.B2(n_35),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_199),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_168),
.A3(n_184),
.B1(n_171),
.B2(n_175),
.C1(n_183),
.C2(n_185),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_204),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_203),
.C(n_196),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_168),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_14),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_187),
.B1(n_190),
.B2(n_195),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_200),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_212),
.B1(n_14),
.B2(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_205),
.C(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_214),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_15),
.C(n_18),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_207),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_217),
.B(n_216),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_221),
.B(n_19),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_19),
.B(n_20),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_21),
.Y(n_224)
);


endmodule