module real_jpeg_4439_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g182 ( 
.A(n_0),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_0),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_0),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_0),
.Y(n_296)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_0),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_0),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_1),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_1),
.A2(n_127),
.B1(n_218),
.B2(n_287),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_1),
.A2(n_218),
.B1(n_298),
.B2(n_394),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g454 ( 
.A1(n_1),
.A2(n_218),
.B1(n_455),
.B2(n_457),
.Y(n_454)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_2),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_2),
.Y(n_204)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_3),
.A2(n_89),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_3),
.A2(n_89),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_4),
.A2(n_33),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_4),
.A2(n_203),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_4),
.A2(n_203),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_4),
.A2(n_203),
.B1(n_428),
.B2(n_431),
.Y(n_427)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_20),
.B(n_513),
.Y(n_19)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_6),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_7),
.Y(n_388)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_140),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_10),
.A2(n_140),
.B1(n_273),
.B2(n_284),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_10),
.A2(n_140),
.B1(n_195),
.B2(n_318),
.Y(n_317)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_12),
.Y(n_517)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_13),
.A2(n_176),
.B1(n_233),
.B2(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_13),
.B(n_388),
.C(n_389),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_13),
.B(n_70),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_13),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_13),
.B(n_114),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_13),
.B(n_226),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_14),
.A2(n_55),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_14),
.A2(n_55),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_14),
.A2(n_55),
.B1(n_232),
.B2(n_239),
.Y(n_292)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_16),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_16),
.A2(n_49),
.B1(n_183),
.B2(n_188),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_16),
.A2(n_49),
.B1(n_238),
.B2(n_243),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_16),
.A2(n_49),
.B1(n_223),
.B2(n_335),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_17),
.A2(n_84),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_17),
.A2(n_84),
.B1(n_183),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_17),
.A2(n_84),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_18),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_18),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_18),
.A2(n_207),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_18),
.A2(n_207),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_18),
.A2(n_207),
.B1(n_319),
.B2(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_156),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_154),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_131),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_23),
.B(n_131),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_119),
.B2(n_120),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_56),
.C(n_90),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_26),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_27),
.A2(n_44),
.B1(n_50),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_27),
.A2(n_37),
.B1(n_202),
.B2(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_27),
.A2(n_268),
.B(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_28),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_28),
.A2(n_263),
.B(n_267),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_32),
.Y(n_170)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_33),
.Y(n_208)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_34),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_34),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_37),
.B(n_176),
.Y(n_323)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_41),
.Y(n_166)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_41),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_43),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_43),
.Y(n_220)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_43),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_43),
.Y(n_337)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_50),
.A2(n_202),
.B(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_51),
.B(n_206),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_51),
.B(n_139),
.Y(n_370)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_56),
.A2(n_90),
.B1(n_91),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_79),
.B1(n_85),
.B2(n_86),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_57),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_57),
.A2(n_79),
.B1(n_85),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_57),
.A2(n_85),
.B1(n_215),
.B2(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_57),
.A2(n_85),
.B1(n_283),
.B2(n_334),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_70),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_62),
.Y(n_468)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_64),
.Y(n_226)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_69),
.Y(n_272)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_70),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

AOI22x1_ASAP7_75t_L g280 ( 
.A1(n_70),
.A2(n_122),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_70),
.A2(n_122),
.B1(n_148),
.B2(n_359),
.Y(n_358)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_73),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_74),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_74),
.Y(n_259)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_74),
.Y(n_408)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_74),
.Y(n_471)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_95),
.B1(n_98),
.B2(n_101),
.Y(n_94)
);

INVx11_ASAP7_75t_L g406 ( 
.A(n_75),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_76),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_76),
.Y(n_246)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_77),
.Y(n_472)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_80),
.Y(n_273)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_85),
.B(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_85),
.A2(n_270),
.B(n_315),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_137),
.C(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_90),
.A2(n_91),
.B1(n_145),
.B2(n_146),
.Y(n_502)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_113),
.B(n_115),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_92),
.A2(n_113),
.B1(n_230),
.B2(n_236),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_92),
.A2(n_381),
.B(n_383),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_92),
.A2(n_113),
.B1(n_405),
.B2(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_92),
.A2(n_383),
.B(n_454),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_93),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_93),
.A2(n_114),
.B1(n_237),
.B2(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_93),
.A2(n_114),
.B1(n_292),
.B2(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_93),
.A2(n_114),
.B1(n_342),
.B2(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_104),
.A2(n_256),
.B(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_112),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_108),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_109),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_111),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_111),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_113),
.A2(n_230),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_114),
.B(n_257),
.Y(n_383)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_115),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_117),
.Y(n_345)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_117),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_214),
.B(n_221),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_122),
.B(n_281),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_122),
.A2(n_221),
.B(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_129),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_143),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_508)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_136),
.A2(n_137),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_143),
.A2(n_144),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_497),
.B(n_510),
.Y(n_156)
);

OAI311xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_327),
.A3(n_374),
.B1(n_491),
.C1(n_496),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_305),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_160),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_274),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_161),
.B(n_274),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_227),
.C(n_254),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_162),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_199),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_163),
.B(n_200),
.C(n_213),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_164),
.A2(n_177),
.B1(n_178),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_164),
.Y(n_312)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.A3(n_168),
.B1(n_171),
.B2(n_175),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_SL g263 ( 
.A1(n_175),
.A2(n_176),
.B(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_176),
.A2(n_179),
.B(n_397),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_SL g460 ( 
.A1(n_176),
.A2(n_335),
.B(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_186),
.B1(n_189),
.B2(n_192),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_179),
.A2(n_249),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_179),
.A2(n_297),
.B(n_347),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_179),
.A2(n_393),
.B(n_397),
.Y(n_392)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_180),
.A2(n_193),
.B1(n_248),
.B2(n_252),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_180),
.A2(n_187),
.B1(n_317),
.B2(n_322),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_180),
.B(n_400),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_180),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_182),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_182),
.Y(n_423)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_182),
.Y(n_435)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_185),
.Y(n_302)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_185),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_185),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_198),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_212),
.B2(n_213),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_205),
.B(n_370),
.Y(n_369)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_227),
.A2(n_228),
.B1(n_254),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_247),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_229),
.B(n_247),
.Y(n_278)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_242),
.Y(n_386)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_246),
.Y(n_382)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_250),
.Y(n_401)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_251),
.Y(n_390)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.C(n_269),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_255),
.B(n_269),
.Y(n_308)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g466 ( 
.A1(n_259),
.A2(n_273),
.A3(n_462),
.B1(n_467),
.B2(n_469),
.Y(n_466)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_260),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_261),
.A2(n_262),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_275),
.B(n_290),
.C(n_303),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_290),
.B1(n_303),
.B2(n_304),
.Y(n_276)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_278),
.B(n_280),
.C(n_289),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_293),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_324),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_306),
.B(n_324),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.C(n_313),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_307),
.B(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_310),
.A2(n_311),
.B1(n_313),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_313),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.C(n_323),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_314),
.B(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_316),
.B(n_323),
.Y(n_482)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_317),
.Y(n_465)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_371),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_328),
.A2(n_371),
.B(n_492),
.C(n_495),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_352),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_329),
.B(n_352),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_339),
.C(n_351),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g373 ( 
.A(n_330),
.B(n_339),
.CI(n_351),
.CON(n_373),
.SN(n_373)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_333),
.C(n_338),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_346),
.B2(n_350),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_346),
.Y(n_366)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_346),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_346),
.A2(n_350),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_346),
.A2(n_366),
.B(n_369),
.Y(n_500)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_353),
.B(n_356),
.C(n_364),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_364),
.B2(n_365),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_360),
.B(n_363),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_361),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_363),
.B(n_500),
.CI(n_501),
.CON(n_499),
.SN(n_499)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_363),
.B(n_500),
.C(n_501),
.Y(n_509)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_372),
.B(n_373),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g519 ( 
.A(n_373),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_485),
.B(n_490),
.Y(n_374)
);

AO21x1_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_474),
.B(n_484),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_448),
.B(n_473),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_411),
.B(n_447),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_391),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_379),
.B(n_391),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_380),
.A2(n_384),
.B1(n_385),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_402),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_403),
.C(n_410),
.Y(n_449)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_409),
.B2(n_410),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_406),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_439),
.B(n_446),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_425),
.B(n_438),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_424),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_421),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

INVx8_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_437),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_437),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_433),
.B(n_436),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_427),
.Y(n_441)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx5_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_435),
.A2(n_436),
.B(n_465),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_444),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_444),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_450),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_463),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_458),
.B2(n_459),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_458),
.C(n_463),
.Y(n_475)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_466),
.Y(n_480)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_472),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_475),
.B(n_476),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_478),
.B1(n_481),
.B2(n_483),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_480),
.C(n_483),
.Y(n_486)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_481),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_486),
.B(n_487),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_505),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_504),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_504),
.Y(n_511)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_499),
.Y(n_520)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_502),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_511),
.B(n_512),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_509),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_509),
.Y(n_512)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_517),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx13_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);


endmodule