module fake_netlist_1_2979_n_679 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_679);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_679;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_47), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_28), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_48), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_3), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_7), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_44), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_22), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_57), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_6), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_24), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_41), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_34), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_72), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_18), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_1), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_21), .Y(n_92) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_13), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_39), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_35), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_51), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_67), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_69), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_55), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_61), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_16), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_71), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_14), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_26), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_31), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_59), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_2), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_25), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_58), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_5), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_7), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_104), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_112), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_85), .B(n_0), .Y(n_130) );
NAND2xp33_ASAP7_75t_R g131 ( .A(n_86), .B(n_0), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_112), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_82), .B(n_1), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_85), .B(n_3), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_122), .B(n_4), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_122), .B(n_4), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_81), .B(n_5), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_112), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_78), .B(n_8), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_78), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_105), .B(n_8), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_96), .A2(n_40), .B(n_74), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_88), .B(n_9), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_123), .B(n_10), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_99), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_107), .B(n_10), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_110), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_92), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_119), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_108), .B(n_11), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_79), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_98), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_165), .B(n_97), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_165), .B(n_87), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_142), .B(n_116), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_130), .B(n_102), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_126), .B(n_111), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
INVx5_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_126), .B(n_115), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_142), .B(n_100), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_129), .B(n_109), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_128), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_129), .B(n_94), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_128), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_140), .B(n_94), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_140), .A2(n_117), .B1(n_106), .B2(n_103), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_146), .B(n_80), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_130), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_134), .Y(n_197) );
INVx1_ASAP7_75t_SL g198 ( .A(n_133), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_134), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_149), .B(n_86), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_127), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_149), .A2(n_124), .B1(n_91), .B2(n_114), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_153), .B(n_89), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_153), .B(n_89), .Y(n_209) );
NOR2xp33_ASAP7_75t_SL g210 ( .A(n_159), .B(n_120), .Y(n_210) );
INVx4_ASAP7_75t_SL g211 ( .A(n_138), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
AND2x6_ASAP7_75t_L g213 ( .A(n_138), .B(n_113), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_127), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_166), .B(n_120), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_159), .B(n_118), .Y(n_216) );
AND2x6_ASAP7_75t_L g217 ( .A(n_138), .B(n_101), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_138), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_160), .B(n_118), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_146), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
INVxp67_ASAP7_75t_SL g222 ( .A(n_160), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_133), .B(n_124), .C(n_114), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_162), .B(n_101), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_166), .B(n_91), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_125), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_125), .Y(n_227) );
NAND3xp33_ASAP7_75t_L g228 ( .A(n_133), .B(n_11), .C(n_12), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_161), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_125), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_222), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_226), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_227), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_230), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_174), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_222), .Y(n_237) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_210), .B(n_154), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_214), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_197), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g241 ( .A1(n_198), .A2(n_155), .B1(n_154), .B2(n_161), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_192), .B(n_154), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_173), .A2(n_155), .B1(n_131), .B2(n_162), .Y(n_243) );
BUFx4f_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
BUFx4f_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_192), .B(n_155), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
AOI22x1_ASAP7_75t_L g249 ( .A1(n_218), .A2(n_156), .B1(n_158), .B2(n_147), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_197), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_217), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_218), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_168), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_221), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_200), .B(n_125), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_201), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_168), .Y(n_258) );
OR2x6_ASAP7_75t_L g259 ( .A(n_173), .B(n_144), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_200), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_209), .B(n_125), .Y(n_262) );
AND2x6_ASAP7_75t_L g263 ( .A(n_178), .B(n_136), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_229), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_223), .A2(n_131), .B1(n_164), .B2(n_144), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_175), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_174), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_225), .B(n_141), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_217), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_217), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_219), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_217), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_224), .B(n_141), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_213), .A2(n_148), .B1(n_164), .B2(n_157), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_171), .B(n_167), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_224), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_177), .Y(n_278) );
INVx5_ASAP7_75t_L g279 ( .A(n_213), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_177), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_211), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_175), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_210), .B(n_136), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_211), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_202), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_195), .B(n_157), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_202), .B(n_148), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_179), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_177), .Y(n_290) );
BUFx12f_ASAP7_75t_L g291 ( .A(n_195), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_175), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_213), .A2(n_167), .B1(n_136), .B2(n_139), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_181), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_228), .B(n_151), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_215), .B(n_139), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_177), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_236), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_231), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_288), .B(n_190), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_259), .B(n_211), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_291), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_291), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_281), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_253), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_233), .A2(n_193), .B1(n_169), .B2(n_184), .C(n_186), .Y(n_307) );
INVx4_ASAP7_75t_SL g308 ( .A(n_263), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_241), .B(n_193), .C(n_216), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_274), .B(n_176), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_274), .B(n_206), .Y(n_311) );
CKINVDCx8_ASAP7_75t_R g312 ( .A(n_239), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_259), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_281), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_259), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_257), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_287), .B(n_189), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_287), .B(n_196), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_256), .A2(n_212), .B(n_208), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_287), .B(n_205), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_288), .B(n_207), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_268), .B(n_199), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_239), .B(n_176), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_281), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_236), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_268), .B(n_184), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_246), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_267), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_244), .B(n_180), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_248), .Y(n_332) );
CKINVDCx11_ASAP7_75t_R g333 ( .A(n_284), .Y(n_333) );
AND3x1_ASAP7_75t_SL g334 ( .A(n_286), .B(n_13), .C(n_14), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_257), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_240), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_243), .B(n_186), .Y(n_337) );
INVx5_ASAP7_75t_L g338 ( .A(n_263), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_238), .A2(n_180), .B1(n_167), .B2(n_136), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_260), .B(n_180), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_263), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_261), .B(n_180), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_238), .A2(n_167), .B1(n_136), .B2(n_143), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_271), .B(n_167), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_286), .A2(n_139), .B1(n_143), .B2(n_150), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_267), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_264), .B(n_139), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_255), .Y(n_348) );
CKINVDCx16_ASAP7_75t_R g349 ( .A(n_335), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_332), .Y(n_350) );
INVx4_ASAP7_75t_SL g351 ( .A(n_301), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_310), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_320), .A2(n_277), .B(n_272), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_348), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_299), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_305), .A2(n_247), .B1(n_242), .B2(n_263), .Y(n_356) );
OAI211xp5_ASAP7_75t_L g357 ( .A1(n_307), .A2(n_265), .B(n_275), .C(n_264), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_313), .A2(n_263), .B1(n_289), .B2(n_276), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_343), .A2(n_151), .B(n_249), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_328), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_338), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_324), .B(n_284), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_337), .A2(n_263), .B1(n_251), .B2(n_240), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_309), .A2(n_251), .B1(n_245), .B2(n_244), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_327), .A2(n_283), .B(n_262), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_336), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_L g368 ( .A1(n_322), .A2(n_296), .B(n_283), .C(n_143), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_316), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_300), .A2(n_245), .B1(n_244), .B2(n_252), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_303), .B(n_279), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_302), .B(n_279), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_304), .Y(n_374) );
NOR2xp67_ASAP7_75t_L g375 ( .A(n_304), .B(n_279), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_344), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_306), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_319), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_345), .A2(n_245), .B1(n_293), .B2(n_273), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_273), .B1(n_269), .B2(n_270), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_373), .A2(n_300), .B1(n_322), .B2(n_329), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_373), .A2(n_329), .B1(n_315), .B2(n_340), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_351), .B(n_308), .Y(n_384) );
BUFx4f_ASAP7_75t_SL g385 ( .A(n_369), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_363), .A2(n_339), .B1(n_323), .B2(n_347), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_357), .A2(n_311), .B(n_340), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_376), .A2(n_150), .B1(n_139), .B2(n_143), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_376), .A2(n_321), .B1(n_317), .B2(n_318), .C(n_143), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_349), .A2(n_312), .B1(n_338), .B2(n_279), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_353), .A2(n_338), .B1(n_341), .B2(n_326), .Y(n_393) );
OR2x6_ASAP7_75t_L g394 ( .A(n_366), .B(n_341), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_366), .A2(n_334), .B1(n_338), .B2(n_279), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_350), .B(n_342), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_374), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_350), .A2(n_150), .B1(n_295), .B2(n_163), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_354), .A2(n_295), .B1(n_163), .B2(n_147), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_355), .B(n_333), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_356), .A2(n_346), .B1(n_326), .B2(n_295), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
OR2x6_ASAP7_75t_L g404 ( .A(n_361), .B(n_314), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_354), .B(n_314), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_355), .B(n_333), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_360), .A2(n_295), .B1(n_163), .B2(n_147), .Y(n_407) );
NOR2xp67_ASAP7_75t_R g408 ( .A(n_351), .B(n_304), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_396), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_385), .B(n_375), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_399), .A2(n_359), .B(n_407), .Y(n_412) );
OAI31xp33_ASAP7_75t_L g413 ( .A1(n_386), .A2(n_362), .A3(n_379), .B(n_371), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_405), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_384), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_395), .B(n_156), .C(n_364), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_389), .B(n_351), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_385), .A2(n_334), .B1(n_380), .B2(n_367), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_389), .B(n_378), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_384), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_382), .B(n_367), .Y(n_421) );
OAI33xp33_ASAP7_75t_L g422 ( .A1(n_400), .A2(n_158), .A3(n_377), .B1(n_137), .B2(n_145), .B3(n_135), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_388), .A2(n_398), .B(n_399), .Y(n_423) );
NAND4xp25_ASAP7_75t_L g424 ( .A(n_406), .B(n_163), .C(n_158), .D(n_372), .Y(n_424) );
OAI22xp5_ASAP7_75t_SL g425 ( .A1(n_387), .A2(n_358), .B1(n_370), .B2(n_377), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_392), .A2(n_163), .B(n_368), .C(n_365), .Y(n_426) );
OA21x2_ASAP7_75t_L g427 ( .A1(n_407), .A2(n_359), .B(n_151), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_382), .A2(n_378), .B1(n_346), .B2(n_270), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_383), .A2(n_280), .B1(n_278), .B2(n_290), .C(n_249), .Y(n_429) );
OAI321xp33_ASAP7_75t_L g430 ( .A1(n_398), .A2(n_156), .A3(n_331), .B1(n_135), .B2(n_137), .C(n_145), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_383), .B(n_232), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_397), .B(n_156), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_384), .B(n_308), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_403), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_391), .A2(n_252), .B1(n_269), .B2(n_325), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_401), .B(n_156), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_404), .B(n_156), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_390), .A2(n_297), .B1(n_331), .B2(n_325), .C(n_235), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_401), .B(n_156), .Y(n_440) );
AOI211xp5_ASAP7_75t_SL g441 ( .A1(n_402), .A2(n_308), .B(n_297), .C(n_135), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
AND2x4_ASAP7_75t_SL g443 ( .A(n_404), .B(n_330), .Y(n_443) );
OAI31xp33_ASAP7_75t_SL g444 ( .A1(n_393), .A2(n_235), .A3(n_234), .B(n_232), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_418), .B(n_390), .C(n_132), .D(n_145), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_409), .B(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_410), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_421), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_421), .Y(n_451) );
OAI31xp33_ASAP7_75t_L g452 ( .A1(n_424), .A2(n_297), .A3(n_234), .B(n_137), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_414), .B(n_419), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_434), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_412), .B(n_404), .Y(n_459) );
AOI21xp5_ASAP7_75t_SL g460 ( .A1(n_419), .A2(n_394), .B(n_330), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_413), .A2(n_132), .B(n_304), .C(n_204), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_437), .B(n_394), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_423), .B(n_132), .C(n_16), .D(n_17), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_427), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_431), .A2(n_292), .B(n_294), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_437), .B(n_15), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_15), .Y(n_468) );
AND2x4_ASAP7_75t_SL g469 ( .A(n_417), .B(n_330), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_419), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_432), .B(n_132), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_425), .A2(n_330), .B1(n_298), .B2(n_285), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_442), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_438), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_432), .B(n_438), .C(n_426), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_436), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_442), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_415), .B(n_204), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_415), .B(n_204), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_436), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_415), .B(n_20), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_415), .B(n_23), .Y(n_482) );
OAI21x1_ASAP7_75t_L g483 ( .A1(n_427), .A2(n_258), .B(n_294), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_415), .B(n_27), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_422), .A2(n_298), .B1(n_188), .B2(n_183), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_417), .A2(n_298), .B1(n_285), .B2(n_188), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_440), .B(n_29), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_444), .B(n_188), .C(n_183), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_417), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g492 ( .A1(n_411), .A2(n_181), .B1(n_183), .B2(n_203), .C1(n_298), .C2(n_194), .Y(n_492) );
OA211x2_ASAP7_75t_L g493 ( .A1(n_416), .A2(n_30), .B(n_33), .C(n_37), .Y(n_493) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_430), .A2(n_292), .B(n_282), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g495 ( .A1(n_420), .A2(n_191), .A3(n_172), .B1(n_182), .B2(n_187), .B3(n_170), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_459), .B(n_420), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_451), .B(n_427), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_449), .B(n_443), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_451), .B(n_441), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_450), .B(n_443), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_463), .B(n_435), .C(n_429), .D(n_439), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_456), .Y(n_502) );
NAND3xp33_ASAP7_75t_L g503 ( .A(n_495), .B(n_428), .C(n_181), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_445), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_449), .B(n_433), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_490), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_459), .B(n_433), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_469), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_445), .B(n_433), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_457), .B(n_38), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_448), .B(n_203), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_457), .B(n_42), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_465), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_465), .B(n_203), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_453), .B(n_45), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_453), .B(n_46), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_454), .B(n_49), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_473), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_454), .B(n_50), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_455), .B(n_52), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_458), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_458), .B(n_53), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_476), .B(n_54), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_455), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_477), .B(n_56), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_476), .B(n_62), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_473), .A2(n_64), .B(n_65), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_480), .B(n_66), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_447), .B(n_485), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_446), .B(n_254), .C(n_266), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_470), .B(n_68), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_485), .B(n_70), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_464), .B(n_75), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_491), .B(n_254), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_468), .B(n_250), .C(n_258), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_468), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_491), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_467), .B(n_266), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_470), .B(n_282), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_462), .B(n_250), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_474), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_475), .B(n_250), .C(n_452), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_462), .B(n_250), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_483), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_469), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_460), .B(n_250), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_489), .A2(n_488), .B1(n_472), .B2(n_493), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_481), .B(n_482), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_471), .A2(n_461), .B(n_488), .C(n_482), .Y(n_552) );
NAND2x1_ASAP7_75t_SL g553 ( .A(n_518), .B(n_484), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_502), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_513), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_497), .B(n_466), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_529), .B(n_466), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_537), .B(n_460), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_501), .B(n_518), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_496), .B(n_478), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_518), .B(n_478), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_524), .B(n_492), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_504), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_541), .B(n_486), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_496), .B(n_479), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_541), .B(n_479), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_503), .B(n_487), .C(n_494), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_496), .B(n_494), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_508), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_496), .B(n_494), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_507), .B(n_494), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
NOR2xp33_ASAP7_75t_R g573 ( .A(n_548), .B(n_550), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_544), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_503), .B(n_552), .C(n_545), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_509), .B(n_506), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_509), .B(n_505), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_549), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_498), .B(n_499), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_500), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_498), .B(n_507), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_520), .Y(n_584) );
XOR2xp5_ASAP7_75t_L g585 ( .A(n_551), .B(n_520), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_538), .B(n_521), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_521), .B(n_551), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_532), .B(n_526), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_514), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_545), .A2(n_536), .B(n_549), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_532), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_532), .B(n_536), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_551), .B(n_526), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_534), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_499), .B(n_551), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_523), .B(n_528), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_554), .B(n_546), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_576), .B(n_516), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_559), .B(n_516), .Y(n_602) );
OAI31xp33_ASAP7_75t_L g603 ( .A1(n_575), .A2(n_559), .A3(n_593), .B(n_588), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_581), .B(n_522), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_563), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_572), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_586), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_583), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_562), .B(n_525), .C(n_532), .D(n_523), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_578), .B(n_519), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
AOI322xp5_ASAP7_75t_L g612 ( .A1(n_584), .A2(n_569), .A3(n_580), .B1(n_597), .B2(n_593), .C1(n_579), .C2(n_587), .Y(n_612) );
CKINVDCx16_ASAP7_75t_R g613 ( .A(n_573), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_586), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_582), .B(n_528), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_589), .B(n_522), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_558), .B(n_533), .Y(n_617) );
NAND2xp33_ASAP7_75t_L g618 ( .A(n_573), .B(n_533), .Y(n_618) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_567), .B(n_510), .C(n_512), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_588), .A2(n_512), .B1(n_540), .B2(n_546), .Y(n_620) );
AOI211x1_ASAP7_75t_L g621 ( .A1(n_590), .A2(n_527), .B(n_534), .C(n_517), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_577), .Y(n_622) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_591), .B(n_515), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_595), .B(n_587), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_553), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_566), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_557), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_594), .B(n_542), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_591), .B(n_519), .Y(n_630) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_591), .B(n_540), .Y(n_631) );
AO21x1_ASAP7_75t_L g632 ( .A1(n_561), .A2(n_511), .B(n_539), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_585), .B(n_531), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g634 ( .A(n_560), .B(n_543), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_561), .A2(n_547), .B(n_598), .C(n_571), .Y(n_635) );
XNOR2x1_ASAP7_75t_L g636 ( .A(n_560), .B(n_565), .Y(n_636) );
OAI322xp33_ASAP7_75t_L g637 ( .A1(n_592), .A2(n_564), .A3(n_596), .B1(n_556), .B2(n_565), .C1(n_570), .C2(n_568), .Y(n_637) );
XOR2x2_ASAP7_75t_L g638 ( .A(n_571), .B(n_568), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_556), .B(n_571), .Y(n_639) );
XNOR2x1_ASAP7_75t_L g640 ( .A(n_570), .B(n_239), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_588), .A2(n_575), .B1(n_585), .B2(n_591), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_559), .A2(n_575), .B1(n_573), .B2(n_562), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_554), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_559), .A2(n_575), .B1(n_418), .B2(n_463), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_585), .B(n_214), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_643), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_601), .Y(n_647) );
XOR2xp5_ASAP7_75t_L g648 ( .A(n_613), .B(n_645), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_618), .A2(n_603), .B(n_641), .Y(n_649) );
AOI32xp33_ASAP7_75t_L g650 ( .A1(n_642), .A2(n_640), .A3(n_636), .B1(n_630), .B2(n_635), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_612), .B(n_626), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_619), .A2(n_633), .B(n_609), .C(n_632), .Y(n_652) );
AO22x2_ASAP7_75t_L g653 ( .A1(n_619), .A2(n_621), .B1(n_622), .B2(n_614), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_637), .A2(n_620), .B(n_602), .C(n_639), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_644), .A2(n_617), .B(n_599), .Y(n_655) );
CKINVDCx16_ASAP7_75t_R g656 ( .A(n_644), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_617), .A2(n_625), .B1(n_630), .B2(n_620), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_606), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_656), .B(n_627), .Y(n_659) );
OAI211xp5_ASAP7_75t_L g660 ( .A1(n_650), .A2(n_604), .B(n_623), .C(n_615), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_658), .Y(n_661) );
AOI211xp5_ASAP7_75t_SL g662 ( .A1(n_649), .A2(n_615), .B(n_600), .C(n_616), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_651), .A2(n_638), .B1(n_610), .B2(n_628), .Y(n_663) );
INVxp33_ASAP7_75t_SL g664 ( .A(n_648), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_647), .Y(n_665) );
OR3x2_ASAP7_75t_L g666 ( .A(n_653), .B(n_624), .C(n_629), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_665), .B(n_652), .Y(n_667) );
NAND3xp33_ASAP7_75t_SL g668 ( .A(n_660), .B(n_657), .C(n_654), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_664), .B(n_655), .C(n_653), .D(n_646), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_659), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_670), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_667), .B(n_661), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_668), .Y(n_673) );
OAI221xp5_ASAP7_75t_R g674 ( .A1(n_673), .A2(n_663), .B1(n_669), .B2(n_666), .C(n_662), .Y(n_674) );
AND3x4_ASAP7_75t_L g675 ( .A(n_672), .B(n_663), .C(n_607), .Y(n_675) );
XNOR2x1_ASAP7_75t_L g676 ( .A(n_675), .B(n_672), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_676), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_671), .B1(n_674), .B2(n_631), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_605), .B1(n_608), .B2(n_634), .C(n_611), .Y(n_679) );
endmodule