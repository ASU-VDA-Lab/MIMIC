module fake_jpeg_22771_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_121;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_50),
.A2(n_57),
.B1(n_28),
.B2(n_2),
.Y(n_114)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_68),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_53),
.B(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_58),
.B(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_81),
.B1(n_18),
.B2(n_30),
.Y(n_100)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_71),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_38),
.B1(n_26),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_37),
.B1(n_33),
.B2(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_74),
.Y(n_110)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_33),
.CON(n_81),
.SN(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_27),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_43),
.B(n_19),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_17),
.B(n_16),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_59),
.B1(n_68),
.B2(n_65),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_104),
.Y(n_133)
);

OA22x2_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_36),
.B1(n_30),
.B2(n_20),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_56),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_59),
.B1(n_75),
.B2(n_77),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_114),
.B1(n_15),
.B2(n_7),
.Y(n_151)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_81),
.B1(n_52),
.B2(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_56),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_36),
.C(n_30),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_36),
.C(n_20),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_28),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_122),
.B(n_123),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_70),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_108),
.Y(n_173)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_130),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_79),
.B1(n_57),
.B2(n_50),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_1),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_131),
.B(n_136),
.Y(n_183)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_135),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_88),
.B(n_86),
.C(n_55),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_146),
.B1(n_151),
.B2(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_139),
.Y(n_167)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_55),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_91),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_55),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_149),
.B1(n_101),
.B2(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_148),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_6),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_153),
.Y(n_169)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_6),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_152),
.Y(n_180)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_112),
.C(n_90),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_171),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_161),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_8),
.Y(n_208)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_174),
.B1(n_177),
.B2(n_149),
.Y(n_193)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_101),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_111),
.B1(n_120),
.B2(n_118),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_108),
.B1(n_102),
.B2(n_106),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_6),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_144),
.B1(n_131),
.B2(n_143),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_193),
.B1(n_195),
.B2(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_128),
.B1(n_144),
.B2(n_102),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_204),
.B1(n_208),
.B2(n_184),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_127),
.B1(n_118),
.B2(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_202),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_207),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_170),
.B1(n_183),
.B2(n_164),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_220),
.B1(n_154),
.B2(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_217),
.B1(n_222),
.B2(n_224),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_221),
.C(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_171),
.B1(n_169),
.B2(n_156),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_169),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

OAI22x1_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_188),
.B1(n_160),
.B2(n_189),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_172),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_158),
.B(n_90),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_204),
.A3(n_181),
.B1(n_168),
.B2(n_163),
.C1(n_161),
.C2(n_189),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_203),
.B1(n_194),
.B2(n_190),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_238),
.B1(n_243),
.B2(n_148),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_95),
.C(n_121),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_235),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_206),
.B1(n_186),
.B2(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_239),
.B1(n_103),
.B2(n_9),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_215),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_158),
.B1(n_155),
.B2(n_182),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_225),
.B(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_162),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_241),
.B(n_240),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_247),
.B(n_257),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_225),
.B(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_138),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_221),
.B1(n_219),
.B2(n_95),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_253),
.C(n_242),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_121),
.C(n_104),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_93),
.B1(n_103),
.B2(n_11),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_239),
.B(n_237),
.C(n_228),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_232),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_8),
.B(n_9),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_264),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_234),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_266),
.B1(n_247),
.B2(n_245),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_260),
.A2(n_229),
.B(n_246),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_268),
.A2(n_261),
.B(n_257),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_265),
.B1(n_230),
.B2(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_274),
.C(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_255),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_270),
.B(n_241),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_278),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_229),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_277),
.B(n_230),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_271),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_267),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_264),
.B(n_12),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_238),
.B(n_277),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_285),
.B(n_282),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_11),
.B(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_13),
.Y(n_290)
);


endmodule