module fake_jpeg_2830_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_59),
.Y(n_95)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_74),
.B(n_73),
.C(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_97),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_66),
.B1(n_69),
.B2(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_83),
.B1(n_66),
.B2(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_77),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_112),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_113),
.B1(n_76),
.B2(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_70),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_83),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_85),
.B1(n_60),
.B2(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_67),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_22),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_67),
.B1(n_68),
.B2(n_4),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_69),
.B1(n_98),
.B2(n_77),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_127),
.B1(n_129),
.B2(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_131),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_81),
.B1(n_84),
.B2(n_78),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_47),
.B1(n_46),
.B2(n_45),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_81),
.B(n_84),
.C(n_72),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_136),
.B(n_120),
.C(n_135),
.D(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_57),
.B1(n_55),
.B2(n_53),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_1),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_52),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_148),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_151),
.C(n_163),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_101),
.B(n_113),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_153),
.B(n_33),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_147),
.B1(n_156),
.B2(n_8),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_130),
.B1(n_122),
.B2(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_67),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_157),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_2),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_3),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_44),
.C(n_43),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_5),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_41),
.C(n_40),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_171),
.C(n_183),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

OAI321xp33_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_21),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_35),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_181),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_7),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_145),
.B1(n_156),
.B2(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_151),
.B1(n_9),
.B2(n_11),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_31),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_24),
.C(n_23),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_8),
.C(n_11),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_191),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_12),
.C(n_14),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_12),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_169),
.B1(n_173),
.B2(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_21),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_175),
.Y(n_198)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_176),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_166),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_167),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_168),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_185),
.B(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_206),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_196),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_195),
.B(n_172),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_207),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_211),
.B(n_203),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_214),
.B(n_196),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_185),
.C(n_179),
.Y(n_216)
);


endmodule