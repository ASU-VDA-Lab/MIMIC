module fake_jpeg_19349_n_289 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_21),
.B1(n_17),
.B2(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_40),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_45),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

AO22x1_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_33),
.B1(n_30),
.B2(n_19),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_22),
.B1(n_18),
.B2(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_18),
.B1(n_33),
.B2(n_25),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_49),
.Y(n_77)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_21),
.Y(n_78)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_25),
.B1(n_32),
.B2(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_25),
.B1(n_20),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_103)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_30),
.C(n_20),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_40),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_83),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_24),
.B(n_23),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_54),
.C(n_6),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_26),
.B1(n_34),
.B2(n_17),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_93),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_28),
.CI(n_19),
.CON(n_87),
.SN(n_87)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_102),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_34),
.B1(n_27),
.B2(n_26),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_99),
.B1(n_103),
.B2(n_0),
.Y(n_128)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_23),
.B1(n_34),
.B2(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_27),
.B1(n_9),
.B2(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_109),
.B1(n_49),
.B2(n_59),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_68),
.C(n_70),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_0),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_62),
.B(n_11),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_49),
.B(n_66),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_112),
.A2(n_127),
.B(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_76),
.B1(n_89),
.B2(n_84),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_49),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_132),
.C(n_135),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_134),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_54),
.B1(n_69),
.B2(n_72),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_107),
.B1(n_87),
.B2(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_15),
.B(n_5),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_124),
.CON(n_154),
.SN(n_154)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_68),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_85),
.B1(n_77),
.B2(n_72),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_71),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_68),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_71),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_85),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_92),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_98),
.B1(n_105),
.B2(n_97),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_190)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_156),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_144),
.C(n_55),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_87),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_86),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_151),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_169),
.B1(n_118),
.B2(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_161),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_89),
.B1(n_51),
.B2(n_101),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_118),
.B(n_81),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_92),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_77),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_165),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_139),
.B1(n_137),
.B2(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_12),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_128),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_84),
.B1(n_101),
.B2(n_81),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_172),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_123),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_193),
.B1(n_187),
.B2(n_186),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_193),
.B(n_154),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_178),
.B1(n_184),
.B2(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_139),
.B1(n_121),
.B2(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_186),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_127),
.B1(n_71),
.B2(n_70),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_70),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_167),
.C(n_141),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_155),
.B1(n_150),
.B2(n_145),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_12),
.B(n_13),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_144),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_202),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_203),
.B1(n_216),
.B2(n_172),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_180),
.B(n_174),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_199),
.A2(n_200),
.B(n_217),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_164),
.B(n_167),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_209),
.B1(n_169),
.B2(n_158),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_143),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_147),
.B1(n_163),
.B2(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_215),
.C(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_196),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_205),
.B(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_179),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_167),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_173),
.B1(n_176),
.B2(n_184),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_141),
.B(n_145),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_212),
.B1(n_158),
.B2(n_181),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_224),
.C(n_236),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_165),
.C(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_194),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_183),
.B1(n_182),
.B2(n_191),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_199),
.B1(n_213),
.B2(n_216),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_171),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_237),
.B(n_218),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_202),
.C(n_215),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_200),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_217),
.C(n_213),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_245),
.C(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_198),
.C(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_241),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_158),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_181),
.B1(n_171),
.B2(n_158),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_259),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_262),
.C(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_242),
.B(n_248),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_235),
.B(n_231),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_246),
.B1(n_251),
.B2(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_266),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_226),
.B1(n_221),
.B2(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_221),
.B1(n_240),
.B2(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_275),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_264),
.B(n_224),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_170),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_267),
.C(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_239),
.C(n_270),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_263),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_273),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_281),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_271),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_283),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_285),
.B(n_266),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_261),
.Y(n_289)
);


endmodule