module fake_jpeg_5037_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

AOI21xp33_ASAP7_75t_L g8 ( 
.A1(n_3),
.A2(n_0),
.B(n_1),
.Y(n_8)
);

BUFx24_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

AOI21xp33_ASAP7_75t_L g12 ( 
.A1(n_1),
.A2(n_0),
.B(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx6p67_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_21),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_12),
.B(n_13),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_15),
.B(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_5),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_29),
.C(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_21),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_27),
.C(n_28),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_11),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_25),
.B(n_11),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_43),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_17),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_39),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_47)
);

AOI21x1_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_13),
.B(n_34),
.Y(n_48)
);


endmodule