module fake_jpeg_31910_n_63 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NAND2x1p5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_9),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_21),
.B(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_43),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_22),
.C(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_10),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_24),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_48),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_21),
.B(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_53),
.B1(n_11),
.B2(n_13),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_41),
.C(n_44),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.C(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_51),
.C(n_45),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_13),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_3),
.B(n_4),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B(n_3),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_11),
.A3(n_5),
.B1(n_14),
.B2(n_0),
.C1(n_17),
.C2(n_23),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_17),
.Y(n_63)
);


endmodule