module real_aes_10680_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1632;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_0), .Y(n_947) );
AOI21xp33_ASAP7_75t_L g902 ( .A1(n_1), .A2(n_598), .B(n_680), .Y(n_902) );
INVx1_ASAP7_75t_L g927 ( .A(n_1), .Y(n_927) );
INVx1_ASAP7_75t_L g602 ( .A(n_2), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_2), .A2(n_82), .B1(n_640), .B2(n_642), .C(n_643), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_3), .A2(n_276), .B1(n_598), .B2(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g658 ( .A(n_3), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_4), .A2(n_334), .B1(n_1124), .B2(n_1126), .C(n_1132), .Y(n_1123) );
AOI21xp33_ASAP7_75t_L g1156 ( .A1(n_4), .A2(n_600), .B(n_801), .Y(n_1156) );
AOI22xp33_ASAP7_75t_SL g1238 ( .A1(n_5), .A2(n_85), .B1(n_1033), .B2(n_1233), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1254 ( .A(n_5), .Y(n_1254) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_6), .A2(n_7), .B1(n_1298), .B2(n_1311), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_8), .Y(n_296) );
AND2x2_ASAP7_75t_L g323 ( .A(n_8), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_8), .B(n_211), .Y(n_327) );
INVx1_ASAP7_75t_L g382 ( .A(n_8), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_9), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g937 ( .A1(n_10), .A2(n_938), .B(n_940), .C(n_970), .Y(n_937) );
INVxp67_ASAP7_75t_L g368 ( .A(n_11), .Y(n_368) );
OAI222xp33_ASAP7_75t_L g417 ( .A1(n_11), .A2(n_51), .B1(n_267), .B2(n_418), .C1(n_422), .C2(n_428), .Y(n_417) );
INVx1_ASAP7_75t_L g1102 ( .A(n_12), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_13), .A2(n_23), .B1(n_1233), .B2(n_1512), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_13), .A2(n_212), .B1(n_1249), .B2(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1107 ( .A(n_14), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_15), .Y(n_955) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_16), .A2(n_254), .B1(n_1305), .B2(n_1308), .Y(n_1319) );
AOI221xp5_ASAP7_75t_SL g1618 ( .A1(n_17), .A2(n_43), .B1(n_669), .B2(n_1619), .C(n_1620), .Y(n_1618) );
AOI22xp33_ASAP7_75t_L g1636 ( .A1(n_17), .A2(n_43), .B1(n_791), .B2(n_804), .Y(n_1636) );
OAI221xp5_ASAP7_75t_L g1135 ( .A1(n_18), .A2(n_27), .B1(n_329), .B2(n_641), .C(n_644), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_18), .Y(n_1163) );
CKINVDCx14_ASAP7_75t_R g1323 ( .A(n_19), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_20), .A2(n_93), .B1(n_500), .B2(n_502), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_20), .A2(n_35), .B1(n_530), .B2(n_548), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_21), .A2(n_44), .B1(n_441), .B2(n_442), .C(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g660 ( .A(n_21), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_22), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g1531 ( .A1(n_23), .A2(n_104), .B1(n_979), .B2(n_980), .C(n_1532), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1608 ( .A1(n_24), .A2(n_214), .B1(n_1609), .B2(n_1611), .Y(n_1608) );
AOI221xp5_ASAP7_75t_L g1624 ( .A1(n_24), .A2(n_214), .B1(n_1031), .B2(n_1625), .C(n_1627), .Y(n_1624) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_25), .A2(n_236), .B1(n_678), .B2(n_679), .C(n_680), .Y(n_677) );
INVx1_ASAP7_75t_L g706 ( .A(n_25), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_26), .A2(n_826), .B1(n_882), .B2(n_886), .C(n_892), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_26), .A2(n_192), .B1(n_558), .B2(n_919), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_27), .Y(n_1162) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_28), .A2(n_163), .B1(n_556), .B2(n_558), .C(n_560), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_28), .A2(n_235), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g398 ( .A(n_29), .Y(n_398) );
OR2x2_ASAP7_75t_L g432 ( .A(n_29), .B(n_396), .Y(n_432) );
INVx1_ASAP7_75t_L g736 ( .A(n_30), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_30), .A2(n_242), .B1(n_789), .B2(n_791), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g1184 ( .A1(n_31), .A2(n_201), .B1(n_1185), .B2(n_1186), .C(n_1188), .Y(n_1184) );
INVx1_ASAP7_75t_L g1195 ( .A(n_31), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_32), .A2(n_67), .B1(n_494), .B2(n_496), .Y(n_493) );
INVx1_ASAP7_75t_L g546 ( .A(n_32), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_33), .A2(n_253), .B1(n_840), .B2(n_841), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_33), .A2(n_253), .B1(n_642), .B2(n_643), .C(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g371 ( .A(n_34), .Y(n_371) );
OAI222xp33_ASAP7_75t_L g573 ( .A1(n_35), .A2(n_163), .B1(n_170), .B2(n_574), .C1(n_576), .C2(n_580), .Y(n_573) );
INVx1_ASAP7_75t_L g322 ( .A(n_36), .Y(n_322) );
OR2x2_ASAP7_75t_L g326 ( .A(n_36), .B(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g337 ( .A(n_36), .Y(n_337) );
BUFx2_ASAP7_75t_L g510 ( .A(n_36), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_37), .A2(n_222), .B1(n_328), .B2(n_853), .C(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g990 ( .A(n_37), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g1515 ( .A1(n_38), .A2(n_165), .B1(n_1235), .B2(n_1236), .Y(n_1515) );
INVxp33_ASAP7_75t_SL g1539 ( .A(n_38), .Y(n_1539) );
INVx1_ASAP7_75t_L g1171 ( .A(n_39), .Y(n_1171) );
INVxp33_ASAP7_75t_SL g1509 ( .A(n_40), .Y(n_1509) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_40), .A2(n_221), .B1(n_1056), .B2(n_1077), .C(n_1526), .Y(n_1525) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_41), .A2(n_186), .B1(n_541), .B2(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1148 ( .A(n_41), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_42), .Y(n_750) );
INVx1_ASAP7_75t_L g650 ( .A(n_44), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_45), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_46), .A2(n_72), .B1(n_684), .B2(n_685), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_46), .A2(n_72), .B1(n_640), .B2(n_642), .C(n_644), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_47), .A2(n_157), .B1(n_622), .B2(n_792), .Y(n_901) );
INVx1_ASAP7_75t_L g929 ( .A(n_47), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g1232 ( .A1(n_48), .A2(n_198), .B1(n_1033), .B2(n_1233), .Y(n_1232) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_48), .A2(n_260), .B1(n_1077), .B2(n_1256), .C(n_1258), .Y(n_1255) );
INVx1_ASAP7_75t_L g344 ( .A(n_49), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_50), .A2(n_100), .B1(n_317), .B2(n_652), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_50), .A2(n_100), .B1(n_618), .B2(n_894), .Y(n_1141) );
INVxp67_ASAP7_75t_L g366 ( .A(n_51), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_52), .A2(n_217), .B1(n_500), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g859 ( .A(n_52), .Y(n_859) );
INVx1_ASAP7_75t_L g1177 ( .A(n_53), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1082 ( .A(n_54), .Y(n_1082) );
INVx1_ASAP7_75t_L g521 ( .A(n_55), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_55), .A2(n_94), .B1(n_565), .B2(n_569), .C(n_570), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_56), .A2(n_937), .B1(n_1003), .B2(n_1004), .Y(n_936) );
INVx1_ASAP7_75t_L g1004 ( .A(n_56), .Y(n_1004) );
INVx1_ASAP7_75t_L g1127 ( .A(n_57), .Y(n_1127) );
AOI21xp33_ASAP7_75t_L g1146 ( .A1(n_57), .A2(n_441), .B(n_891), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1237 ( .A1(n_58), .A2(n_105), .B1(n_1235), .B2(n_1236), .Y(n_1237) );
INVxp33_ASAP7_75t_SL g1264 ( .A(n_58), .Y(n_1264) );
INVx1_ASAP7_75t_L g1572 ( .A(n_59), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1640 ( .A1(n_59), .A2(n_208), .B1(n_794), .B2(n_805), .Y(n_1640) );
OAI22xp33_ASAP7_75t_L g903 ( .A1(n_60), .A2(n_192), .B1(n_615), .B2(n_618), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_60), .A2(n_273), .B1(n_912), .B2(n_917), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g1622 ( .A(n_61), .Y(n_1622) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_62), .A2(n_124), .B1(n_1021), .B2(n_1023), .Y(n_1020) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_62), .A2(n_147), .B1(n_891), .B2(n_1051), .C(n_1053), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_63), .A2(n_73), .B1(n_441), .B2(n_443), .C(n_679), .Y(n_828) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_63), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_64), .A2(n_210), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_64), .A2(n_279), .B1(n_745), .B2(n_1087), .Y(n_1086) );
AO22x2_ASAP7_75t_L g724 ( .A1(n_65), .A2(n_725), .B1(n_726), .B2(n_812), .Y(n_724) );
INVx1_ASAP7_75t_L g812 ( .A(n_65), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_66), .A2(n_95), .B1(n_1298), .B2(n_1311), .Y(n_1320) );
INVx1_ASAP7_75t_L g544 ( .A(n_67), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_68), .Y(n_760) );
INVx1_ASAP7_75t_L g946 ( .A(n_69), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_69), .A2(n_143), .B1(n_799), .B2(n_998), .C(n_1000), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_70), .Y(n_1084) );
AOI22xp5_ASAP7_75t_SL g1316 ( .A1(n_71), .A2(n_87), .B1(n_1292), .B2(n_1298), .Y(n_1316) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_73), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_74), .A2(n_268), .B1(n_611), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g712 ( .A(n_74), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_75), .A2(n_204), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_75), .A2(n_204), .B1(n_804), .B2(n_805), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_76), .Y(n_748) );
INVx1_ASAP7_75t_L g964 ( .A(n_77), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_77), .A2(n_250), .B1(n_615), .B2(n_618), .Y(n_1002) );
INVxp33_ASAP7_75t_SL g1013 ( .A(n_78), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_78), .A2(n_213), .B1(n_790), .B2(n_792), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_79), .Y(n_1011) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_79), .A2(n_219), .B1(n_685), .B2(n_1041), .C(n_1043), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1173 ( .A1(n_80), .A2(n_148), .B1(n_552), .B2(n_1104), .C(n_1174), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_80), .A2(n_101), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
CKINVDCx16_ASAP7_75t_R g1296 ( .A(n_81), .Y(n_1296) );
INVx1_ASAP7_75t_L g603 ( .A(n_82), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g1129 ( .A(n_83), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1564 ( .A(n_84), .Y(n_1564) );
INVxp33_ASAP7_75t_L g1263 ( .A(n_85), .Y(n_1263) );
INVx1_ASAP7_75t_L g1176 ( .A(n_86), .Y(n_1176) );
AOI221xp5_ASAP7_75t_L g1197 ( .A1(n_86), .A2(n_148), .B1(n_979), .B2(n_1198), .C(n_1199), .Y(n_1197) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_88), .A2(n_161), .B1(n_458), .B2(n_460), .C(n_462), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_88), .A2(n_178), .B1(n_469), .B2(n_474), .C(n_478), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_89), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g1554 ( .A1(n_90), .A2(n_208), .B1(n_1555), .B2(n_1558), .Y(n_1554) );
INVx1_ASAP7_75t_L g1639 ( .A(n_90), .Y(n_1639) );
INVx1_ASAP7_75t_L g396 ( .A(n_91), .Y(n_396) );
INVx1_ASAP7_75t_L g446 ( .A(n_91), .Y(n_446) );
INVx1_ASAP7_75t_L g823 ( .A(n_92), .Y(n_823) );
INVx1_ASAP7_75t_L g563 ( .A(n_93), .Y(n_563) );
INVx1_ASAP7_75t_L g517 ( .A(n_94), .Y(n_517) );
INVx1_ASAP7_75t_L g1189 ( .A(n_96), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_96), .A2(n_201), .B1(n_422), .B2(n_838), .C(n_1194), .Y(n_1193) );
AO221x2_ASAP7_75t_L g1321 ( .A1(n_97), .A2(n_265), .B1(n_1298), .B2(n_1311), .C(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g887 ( .A(n_98), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_98), .A2(n_172), .B1(n_558), .B2(n_910), .Y(n_909) );
NAND2xp33_ASAP7_75t_SL g596 ( .A(n_99), .B(n_502), .Y(n_596) );
INVx1_ASAP7_75t_L g633 ( .A(n_99), .Y(n_633) );
INVxp67_ASAP7_75t_SL g1175 ( .A(n_101), .Y(n_1175) );
INVxp67_ASAP7_75t_SL g1217 ( .A(n_102), .Y(n_1217) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_102), .A2(n_232), .B1(n_992), .B2(n_1245), .Y(n_1244) );
OAI221xp5_ASAP7_75t_L g744 ( .A1(n_103), .A2(n_745), .B1(n_746), .B2(n_752), .C(n_759), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_103), .A2(n_137), .B1(n_799), .B2(n_802), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g1513 ( .A1(n_104), .A2(n_212), .B1(n_1235), .B2(n_1514), .Y(n_1513) );
INVxp67_ASAP7_75t_SL g1243 ( .A(n_105), .Y(n_1243) );
OAI22xp33_ASAP7_75t_L g1139 ( .A1(n_106), .A2(n_164), .B1(n_325), .B2(n_931), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_106), .A2(n_224), .B1(n_420), .B2(n_611), .Y(n_1155) );
INVx1_ASAP7_75t_L g1182 ( .A(n_107), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1204 ( .A1(n_107), .A2(n_159), .B1(n_600), .B2(n_795), .C(n_1205), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_108), .A2(n_224), .B1(n_932), .B2(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1153 ( .A(n_108), .Y(n_1153) );
XNOR2xp5_ASAP7_75t_L g310 ( .A(n_109), .B(n_311), .Y(n_310) );
INVxp33_ASAP7_75t_SL g1017 ( .A(n_110), .Y(n_1017) );
AOI21xp33_ASAP7_75t_L g1046 ( .A1(n_110), .A2(n_1001), .B(n_1047), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_111), .A2(n_878), .B1(n_933), .B2(n_934), .Y(n_877) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_111), .Y(n_933) );
INVxp67_ASAP7_75t_L g339 ( .A(n_112), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_112), .A2(n_181), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_113), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_114), .A2(n_177), .B1(n_460), .B2(n_498), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g540 ( .A1(n_114), .A2(n_335), .B(n_541), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g1167 ( .A1(n_115), .A2(n_1168), .B(n_1191), .Y(n_1167) );
INVx1_ASAP7_75t_L g1211 ( .A(n_115), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_116), .A2(n_255), .B1(n_1305), .B2(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1190 ( .A(n_117), .Y(n_1190) );
CKINVDCx5p33_ASAP7_75t_R g1520 ( .A(n_118), .Y(n_1520) );
INVx1_ASAP7_75t_L g969 ( .A(n_119), .Y(n_969) );
OAI211xp5_ASAP7_75t_SL g971 ( .A1(n_119), .A2(n_972), .B(n_974), .C(n_982), .Y(n_971) );
INVx1_ASAP7_75t_L g1508 ( .A(n_120), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_121), .A2(n_245), .B1(n_836), .B2(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g851 ( .A(n_121), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_122), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_123), .A2(n_176), .B1(n_1031), .B2(n_1033), .Y(n_1030) );
INVxp33_ASAP7_75t_SL g1058 ( .A(n_123), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_124), .A2(n_127), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
AOI22xp33_ASAP7_75t_SL g1516 ( .A1(n_125), .A2(n_141), .B1(n_1233), .B2(n_1517), .Y(n_1516) );
INVxp33_ASAP7_75t_L g1538 ( .A(n_125), .Y(n_1538) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_126), .A2(n_223), .B1(n_598), .B2(n_679), .C(n_680), .Y(n_834) );
INVx1_ASAP7_75t_L g850 ( .A(n_126), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_127), .A2(n_147), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g741 ( .A(n_128), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_128), .A2(n_146), .B1(n_794), .B2(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g288 ( .A(n_129), .Y(n_288) );
INVx1_ASAP7_75t_L g1061 ( .A(n_130), .Y(n_1061) );
INVx1_ASAP7_75t_L g625 ( .A(n_131), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_132), .Y(n_697) );
INVx1_ASAP7_75t_L g722 ( .A(n_133), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_134), .A2(n_193), .B1(n_1026), .B2(n_1027), .Y(n_1029) );
INVxp67_ASAP7_75t_SL g1039 ( .A(n_134), .Y(n_1039) );
INVxp67_ASAP7_75t_SL g1500 ( .A(n_135), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1524 ( .A1(n_135), .A2(n_280), .B1(n_992), .B2(n_1245), .Y(n_1524) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_136), .A2(n_203), .B1(n_452), .B2(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g703 ( .A(n_136), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_137), .A2(n_547), .B1(n_732), .B2(n_734), .C(n_739), .Y(n_731) );
OAI221xp5_ASAP7_75t_SL g1180 ( .A1(n_138), .A2(n_251), .B1(n_543), .B2(n_866), .C(n_1181), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_138), .A2(n_251), .B1(n_790), .B2(n_1207), .Y(n_1206) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_139), .A2(n_237), .B1(n_1305), .B2(n_1308), .Y(n_1315) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_140), .A2(n_227), .B1(n_506), .B2(n_507), .Y(n_595) );
INVx1_ASAP7_75t_L g638 ( .A(n_140), .Y(n_638) );
INVxp67_ASAP7_75t_SL g1536 ( .A(n_141), .Y(n_1536) );
XOR2xp5_ASAP7_75t_L g1120 ( .A(n_142), .B(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g944 ( .A(n_143), .Y(n_944) );
INVx1_ASAP7_75t_L g1015 ( .A(n_144), .Y(n_1015) );
OAI222xp33_ASAP7_75t_L g313 ( .A1(n_145), .A2(n_182), .B1(n_271), .B2(n_314), .C1(n_325), .C2(n_328), .Y(n_313) );
INVx1_ASAP7_75t_L g404 ( .A(n_145), .Y(n_404) );
INVx1_ASAP7_75t_L g740 ( .A(n_146), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_149), .A2(n_150), .B1(n_1292), .B2(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1506 ( .A(n_151), .Y(n_1506) );
CKINVDCx14_ASAP7_75t_R g1324 ( .A(n_152), .Y(n_1324) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_153), .A2(n_240), .B1(n_1305), .B2(n_1308), .Y(n_1304) );
XNOR2xp5_ASAP7_75t_L g485 ( .A(n_154), .B(n_486), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_155), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_156), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_157), .A2(n_263), .B1(n_931), .B2(n_932), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_158), .A2(n_264), .B1(n_789), .B2(n_1056), .Y(n_1070) );
INVx1_ASAP7_75t_L g1091 ( .A(n_158), .Y(n_1091) );
INVx1_ASAP7_75t_L g1183 ( .A(n_159), .Y(n_1183) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_160), .Y(n_696) );
OAI332xp33_ASAP7_75t_L g333 ( .A1(n_161), .A2(n_334), .A3(n_338), .B1(n_349), .B2(n_358), .B3(n_367), .C1(n_376), .C2(n_383), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_162), .Y(n_688) );
INVx1_ASAP7_75t_L g1158 ( .A(n_164), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1523 ( .A(n_165), .Y(n_1523) );
CKINVDCx5p33_ASAP7_75t_R g1568 ( .A(n_166), .Y(n_1568) );
CKINVDCx5p33_ASAP7_75t_R g1240 ( .A(n_167), .Y(n_1240) );
INVx1_ASAP7_75t_L g827 ( .A(n_168), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_169), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_170), .A2(n_235), .B1(n_552), .B2(n_553), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_171), .Y(n_766) );
INVx1_ASAP7_75t_L g884 ( .A(n_172), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g1621 ( .A(n_173), .Y(n_1621) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_174), .A2(n_184), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g533 ( .A(n_174), .Y(n_533) );
INVxp67_ASAP7_75t_SL g959 ( .A(n_175), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_175), .A2(n_205), .B1(n_979), .B2(n_980), .C(n_981), .Y(n_978) );
INVxp67_ASAP7_75t_SL g1049 ( .A(n_176), .Y(n_1049) );
INVx1_ASAP7_75t_L g539 ( .A(n_177), .Y(n_539) );
INVx1_ASAP7_75t_L g456 ( .A(n_178), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_179), .A2(n_243), .B1(n_443), .B2(n_690), .C(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g717 ( .A(n_179), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g890 ( .A1(n_180), .A2(n_790), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_180), .A2(n_262), .B1(n_912), .B2(n_914), .Y(n_911) );
INVx1_ASAP7_75t_L g350 ( .A(n_181), .Y(n_350) );
INVx1_ASAP7_75t_L g450 ( .A(n_182), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_183), .A2(n_279), .B1(n_1072), .B2(n_1073), .Y(n_1075) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_183), .A2(n_210), .B1(n_732), .B2(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g535 ( .A(n_184), .Y(n_535) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_185), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_185), .B(n_288), .Y(n_1279) );
AND3x2_ASAP7_75t_L g1295 ( .A(n_185), .B(n_288), .C(n_1282), .Y(n_1295) );
INVx1_ASAP7_75t_L g1145 ( .A(n_186), .Y(n_1145) );
CKINVDCx16_ASAP7_75t_R g1299 ( .A(n_187), .Y(n_1299) );
AOI22xp5_ASAP7_75t_SL g1331 ( .A1(n_188), .A2(n_200), .B1(n_1292), .B2(n_1298), .Y(n_1331) );
INVx2_ASAP7_75t_L g301 ( .A(n_189), .Y(n_301) );
INVx1_ASAP7_75t_L g842 ( .A(n_190), .Y(n_842) );
AOI22xp5_ASAP7_75t_SL g1330 ( .A1(n_191), .A2(n_258), .B1(n_1305), .B2(n_1308), .Y(n_1330) );
INVxp33_ASAP7_75t_SL g1059 ( .A(n_193), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_194), .Y(n_1226) );
INVx1_ASAP7_75t_L g1170 ( .A(n_195), .Y(n_1170) );
INVxp33_ASAP7_75t_SL g1227 ( .A(n_196), .Y(n_1227) );
AOI221xp5_ASAP7_75t_L g1246 ( .A1(n_196), .A2(n_244), .B1(n_1247), .B2(n_1249), .C(n_1250), .Y(n_1246) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_197), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_198), .A2(n_220), .B1(n_1207), .B2(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1282 ( .A(n_199), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_202), .A2(n_270), .B1(n_541), .B2(n_1131), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_202), .A2(n_270), .B1(n_615), .B2(n_826), .Y(n_1142) );
INVx1_ASAP7_75t_L g707 ( .A(n_203), .Y(n_707) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_205), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_206), .A2(n_256), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
INVx1_ASAP7_75t_L g1097 ( .A(n_206), .Y(n_1097) );
AO221x2_ASAP7_75t_L g1387 ( .A1(n_207), .A2(n_281), .B1(n_1345), .B2(n_1388), .C(n_1389), .Y(n_1387) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_209), .Y(n_676) );
INVx1_ASAP7_75t_L g303 ( .A(n_211), .Y(n_303) );
INVx2_ASAP7_75t_L g324 ( .A(n_211), .Y(n_324) );
INVxp33_ASAP7_75t_SL g1018 ( .A(n_213), .Y(n_1018) );
OR2x2_ASAP7_75t_L g879 ( .A(n_215), .B(n_627), .Y(n_879) );
CKINVDCx14_ASAP7_75t_R g1391 ( .A(n_216), .Y(n_1391) );
INVx1_ASAP7_75t_L g867 ( .A(n_217), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_218), .A2(n_818), .B1(n_875), .B2(n_876), .Y(n_817) );
INVx1_ASAP7_75t_L g876 ( .A(n_218), .Y(n_876) );
INVxp67_ASAP7_75t_SL g1010 ( .A(n_219), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g1234 ( .A1(n_220), .A2(n_260), .B1(n_1235), .B2(n_1236), .Y(n_1234) );
INVxp33_ASAP7_75t_SL g1504 ( .A(n_221), .Y(n_1504) );
INVx1_ASAP7_75t_L g993 ( .A(n_222), .Y(n_993) );
INVx1_ASAP7_75t_L g848 ( .A(n_223), .Y(n_848) );
OAI211xp5_ASAP7_75t_L g1584 ( .A1(n_225), .A2(n_1585), .B(n_1587), .C(n_1592), .Y(n_1584) );
INVx1_ASAP7_75t_L g1631 ( .A(n_225), .Y(n_1631) );
CKINVDCx16_ASAP7_75t_R g1289 ( .A(n_226), .Y(n_1289) );
INVx1_ASAP7_75t_L g631 ( .A(n_227), .Y(n_631) );
INVx1_ASAP7_75t_L g1111 ( .A(n_228), .Y(n_1111) );
INVx1_ASAP7_75t_L g957 ( .A(n_229), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_230), .Y(n_616) );
XOR2xp5_ASAP7_75t_L g1065 ( .A(n_231), .B(n_1066), .Y(n_1065) );
INVxp67_ASAP7_75t_SL g1220 ( .A(n_232), .Y(n_1220) );
INVx1_ASAP7_75t_L g1224 ( .A(n_233), .Y(n_1224) );
INVx1_ASAP7_75t_L g1105 ( .A(n_234), .Y(n_1105) );
INVx1_ASAP7_75t_L g704 ( .A(n_236), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g1569 ( .A(n_238), .Y(n_1569) );
AOI22xp5_ASAP7_75t_L g1494 ( .A1(n_239), .A2(n_1495), .B1(n_1540), .B2(n_1541), .Y(n_1494) );
CKINVDCx5p33_ASAP7_75t_R g1540 ( .A(n_239), .Y(n_1540) );
XOR2x2_ASAP7_75t_L g1212 ( .A(n_240), .B(n_1213), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1601 ( .A1(n_241), .A2(n_257), .B1(n_1602), .B2(n_1604), .Y(n_1601) );
INVx1_ASAP7_75t_L g1628 ( .A(n_241), .Y(n_1628) );
INVx1_ASAP7_75t_L g738 ( .A(n_242), .Y(n_738) );
INVx1_ASAP7_75t_L g713 ( .A(n_243), .Y(n_713) );
INVxp33_ASAP7_75t_SL g1222 ( .A(n_244), .Y(n_1222) );
INVx1_ASAP7_75t_L g846 ( .A(n_245), .Y(n_846) );
INVx1_ASAP7_75t_L g961 ( .A(n_246), .Y(n_961) );
OAI211xp5_ASAP7_75t_L g987 ( .A1(n_246), .A2(n_988), .B(n_989), .C(n_994), .Y(n_987) );
INVx1_ASAP7_75t_L g411 ( .A(n_247), .Y(n_411) );
INVx1_ASAP7_75t_L g1283 ( .A(n_248), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_248), .B(n_1281), .Y(n_1288) );
INVx1_ASAP7_75t_L g833 ( .A(n_249), .Y(n_833) );
INVx1_ASAP7_75t_L g966 ( .A(n_250), .Y(n_966) );
INVx1_ASAP7_75t_L g355 ( .A(n_252), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g1547 ( .A1(n_255), .A2(n_1548), .B1(n_1550), .B2(n_1642), .Y(n_1547) );
AO22x2_ASAP7_75t_L g1550 ( .A1(n_255), .A2(n_1551), .B1(n_1552), .B2(n_1641), .Y(n_1550) );
INVxp67_ASAP7_75t_L g1641 ( .A(n_255), .Y(n_1641) );
INVx1_ASAP7_75t_L g1095 ( .A(n_256), .Y(n_1095) );
INVx1_ASAP7_75t_L g1574 ( .A(n_257), .Y(n_1574) );
INVx2_ASAP7_75t_L g300 ( .A(n_259), .Y(n_300) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_261), .A2(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g637 ( .A(n_261), .Y(n_637) );
INVx1_ASAP7_75t_L g885 ( .A(n_262), .Y(n_885) );
INVx1_ASAP7_75t_L g899 ( .A(n_263), .Y(n_899) );
INVx1_ASAP7_75t_L g1090 ( .A(n_264), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_266), .Y(n_943) );
INVxp67_ASAP7_75t_L g359 ( .A(n_267), .Y(n_359) );
INVx1_ASAP7_75t_L g718 ( .A(n_268), .Y(n_718) );
INVx1_ASAP7_75t_L g698 ( .A(n_269), .Y(n_698) );
INVx1_ASAP7_75t_L g415 ( .A(n_271), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g1284 ( .A(n_272), .Y(n_1284) );
OAI211xp5_ASAP7_75t_SL g893 ( .A1(n_273), .A2(n_894), .B(n_895), .C(n_898), .Y(n_893) );
BUFx3_ASAP7_75t_L g401 ( .A(n_274), .Y(n_401) );
INVx1_ASAP7_75t_L g426 ( .A(n_274), .Y(n_426) );
BUFx3_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
INVx1_ASAP7_75t_L g421 ( .A(n_275), .Y(n_421) );
INVx1_ASAP7_75t_L g653 ( .A(n_276), .Y(n_653) );
INVx1_ASAP7_75t_L g822 ( .A(n_277), .Y(n_822) );
INVx1_ASAP7_75t_L g1036 ( .A(n_278), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1501 ( .A(n_280), .Y(n_1501) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_304), .B(n_1268), .Y(n_282) );
HB1xp67_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x4_ASAP7_75t_L g1549 ( .A(n_286), .B(n_292), .Y(n_1549) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g1546 ( .A(n_287), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_287), .B(n_289), .Y(n_1644) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_289), .B(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x6_ASAP7_75t_L g1581 ( .A(n_294), .B(n_510), .Y(n_1581) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g743 ( .A(n_295), .B(n_303), .Y(n_743) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g335 ( .A(n_296), .B(n_336), .Y(n_335) );
INVx8_ASAP7_75t_L g1573 ( .A(n_297), .Y(n_1573) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
OR2x2_ASAP7_75t_L g325 ( .A(n_298), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_SL g357 ( .A(n_298), .Y(n_357) );
INVx1_ASAP7_75t_L g370 ( .A(n_298), .Y(n_370) );
BUFx2_ASAP7_75t_L g657 ( .A(n_298), .Y(n_657) );
INVx2_ASAP7_75t_SL g858 ( .A(n_298), .Y(n_858) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_298), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g1174 ( .A1(n_298), .A2(n_374), .B1(n_1175), .B2(n_1176), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_298), .A2(n_374), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
OR2x6_ASAP7_75t_L g1576 ( .A(n_298), .B(n_1557), .Y(n_1576) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g318 ( .A(n_300), .Y(n_318) );
AND2x4_ASAP7_75t_L g347 ( .A(n_300), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
INVx1_ASAP7_75t_L g387 ( .A(n_300), .Y(n_387) );
AND2x2_ASAP7_75t_L g473 ( .A(n_300), .B(n_301), .Y(n_473) );
INVx1_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_301), .B(n_318), .Y(n_343) );
INVx2_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
INVx1_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
INVx1_ASAP7_75t_L g481 ( .A(n_301), .Y(n_481) );
AND2x4_ASAP7_75t_L g1570 ( .A(n_302), .B(n_481), .Y(n_1570) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_814), .B2(n_1267), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
XNOR2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_670), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_587), .B2(n_588), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_484), .B1(n_485), .B2(n_586), .Y(n_309) );
INVx1_ASAP7_75t_L g586 ( .A(n_310), .Y(n_586) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_388), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_333), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_315), .A2(n_470), .B1(n_637), .B2(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_315), .A2(n_470), .B1(n_850), .B2(n_851), .Y(n_849) );
INVx1_ASAP7_75t_L g1138 ( .A(n_315), .Y(n_1138) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x2_ASAP7_75t_L g708 ( .A(n_316), .B(n_321), .Y(n_708) );
AND2x2_ASAP7_75t_L g928 ( .A(n_316), .B(n_321), .Y(n_928) );
INVx2_ASAP7_75t_SL g1626 ( .A(n_316), .Y(n_1626) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g534 ( .A(n_317), .B(n_323), .Y(n_534) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_317), .Y(n_552) );
INVx1_ASAP7_75t_L g913 ( .A(n_317), .Y(n_913) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_317), .Y(n_1026) );
BUFx6f_ASAP7_75t_L g1185 ( .A(n_317), .Y(n_1185) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g331 ( .A(n_318), .Y(n_331) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g384 ( .A(n_321), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g470 ( .A(n_321), .B(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g476 ( .A(n_321), .B(n_477), .Y(n_476) );
AND2x6_ASAP7_75t_L g634 ( .A(n_321), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g847 ( .A(n_321), .B(n_364), .Y(n_847) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_321), .B(n_541), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g1179 ( .A1(n_321), .A2(n_921), .B1(n_1180), .B2(n_1184), .Y(n_1179) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g379 ( .A(n_322), .Y(n_379) );
OR2x2_ASAP7_75t_L g579 ( .A(n_322), .B(n_432), .Y(n_579) );
INVx2_ASAP7_75t_L g530 ( .A(n_323), .Y(n_530) );
AND2x4_ASAP7_75t_L g733 ( .A(n_323), .B(n_557), .Y(n_733) );
INVx1_ASAP7_75t_L g336 ( .A(n_324), .Y(n_336) );
INVx1_ASAP7_75t_L g381 ( .A(n_324), .Y(n_381) );
AND2x4_ASAP7_75t_L g627 ( .A(n_325), .B(n_574), .Y(n_627) );
INVx2_ASAP7_75t_L g1178 ( .A(n_325), .Y(n_1178) );
INVx3_ASAP7_75t_L g332 ( .A(n_326), .Y(n_332) );
INVx1_ASAP7_75t_L g549 ( .A(n_327), .Y(n_549) );
BUFx4f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx4f_ASAP7_75t_L g642 ( .A(n_329), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_330), .A2(n_566), .B1(n_1082), .B2(n_1084), .Y(n_1113) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x6_ASAP7_75t_L g569 ( .A(n_331), .B(n_548), .Y(n_569) );
AND2x4_ASAP7_75t_L g479 ( .A(n_332), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g482 ( .A(n_332), .B(n_483), .Y(n_482) );
NAND2x1_ASAP7_75t_SL g641 ( .A(n_332), .B(n_566), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_332), .B(n_635), .Y(n_644) );
AND2x4_ASAP7_75t_L g923 ( .A(n_332), .B(n_924), .Y(n_923) );
OAI33xp33_ASAP7_75t_L g645 ( .A1(n_334), .A2(n_646), .A3(n_654), .B1(n_661), .B2(n_663), .B3(n_667), .Y(n_645) );
OAI33xp33_ASAP7_75t_L g710 ( .A1(n_334), .A2(n_378), .A3(n_711), .B1(n_714), .B2(n_719), .B3(n_721), .Y(n_710) );
OAI33xp33_ASAP7_75t_L g855 ( .A1(n_334), .A2(n_376), .A3(n_856), .B1(n_863), .B2(n_868), .B3(n_872), .Y(n_855) );
OAI33xp33_ASAP7_75t_L g950 ( .A1(n_334), .A2(n_661), .A3(n_951), .B1(n_956), .B2(n_960), .B3(n_965), .Y(n_950) );
OR2x6_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g1557 ( .A(n_336), .Y(n_1557) );
BUFx2_ASAP7_75t_L g467 ( .A(n_337), .Y(n_467) );
INVx2_ASAP7_75t_L g491 ( .A(n_337), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_344), .B2(n_345), .Y(n_338) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g864 ( .A(n_341), .Y(n_864) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_341), .Y(n_1101) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g543 ( .A(n_342), .Y(n_543) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
INVx1_ASAP7_75t_L g649 ( .A(n_343), .Y(n_649) );
OAI221xp5_ASAP7_75t_SL g438 ( .A1(n_344), .A2(n_355), .B1(n_422), .B2(n_439), .C(n_440), .Y(n_438) );
INVx2_ASAP7_75t_SL g1514 ( .A(n_345), .Y(n_1514) );
INVx4_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g737 ( .A(n_346), .Y(n_737) );
INVx2_ASAP7_75t_SL g757 ( .A(n_346), .Y(n_757) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_346), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_346), .Y(n_1092) );
BUFx3_ASAP7_75t_L g1630 ( .A(n_346), .Y(n_1630) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
INVx1_ASAP7_75t_L g532 ( .A(n_347), .Y(n_532) );
INVx1_ASAP7_75t_L g1561 ( .A(n_347), .Y(n_1561) );
AND2x4_ASAP7_75t_L g386 ( .A(n_348), .B(n_387), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_355), .B2(n_356), .Y(n_349) );
OR2x6_ASAP7_75t_L g547 ( .A(n_351), .B(n_548), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_351), .A2(n_664), .B1(n_688), .B2(n_696), .Y(n_721) );
INVx1_ASAP7_75t_L g861 ( .A(n_351), .Y(n_861) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g538 ( .A(n_352), .Y(n_538) );
BUFx2_ASAP7_75t_L g666 ( .A(n_352), .Y(n_666) );
INVx2_ASAP7_75t_L g1094 ( .A(n_352), .Y(n_1094) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_353), .B(n_354), .Y(n_375) );
INVx1_ASAP7_75t_L g925 ( .A(n_354), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_356), .A2(n_665), .B1(n_740), .B2(n_741), .C(n_742), .Y(n_739) );
OAI22xp5_ASAP7_75t_SL g1620 ( .A1(n_356), .A2(n_1621), .B1(n_1622), .B2(n_1623), .Y(n_1620) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_363), .B2(n_366), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_360), .A2(n_952), .B1(n_953), .B2(n_955), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_360), .A2(n_961), .B1(n_962), .B2(n_964), .Y(n_960) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g1555 ( .A(n_362), .B(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g954 ( .A(n_363), .Y(n_954) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g915 ( .A(n_364), .Y(n_915) );
INVx2_ASAP7_75t_L g1187 ( .A(n_364), .Y(n_1187) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g477 ( .A(n_365), .Y(n_477) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_365), .Y(n_554) );
OAI22xp5_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_369), .B1(n_371), .B2(n_372), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g1106 ( .A1(n_369), .A2(n_374), .B1(n_751), .B2(n_1107), .C(n_1108), .Y(n_1106) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g749 ( .A(n_370), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_371), .A2(n_417), .B1(n_431), .B2(n_433), .C(n_436), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_372), .A2(n_664), .B1(n_712), .B2(n_713), .Y(n_711) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g1623 ( .A(n_373), .Y(n_1623) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g659 ( .A(n_374), .Y(n_659) );
BUFx3_ASAP7_75t_L g874 ( .A(n_374), .Y(n_874) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI33xp33_ASAP7_75t_L g1019 ( .A1(n_377), .A2(n_908), .A3(n_1020), .B1(n_1025), .B2(n_1029), .B3(n_1030), .Y(n_1019) );
AOI33xp33_ASAP7_75t_L g1228 ( .A1(n_377), .A2(n_1229), .A3(n_1232), .B1(n_1234), .B2(n_1237), .B3(n_1238), .Y(n_1228) );
AOI33xp33_ASAP7_75t_L g1510 ( .A1(n_377), .A2(n_1229), .A3(n_1511), .B1(n_1513), .B2(n_1515), .B3(n_1516), .Y(n_1510) );
INVx6_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx5_ASAP7_75t_L g662 ( .A(n_378), .Y(n_662) );
OR2x6_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_379), .B(n_394), .Y(n_516) );
INVx2_ASAP7_75t_L g561 ( .A(n_380), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g1567 ( .A(n_381), .Y(n_1567) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_384), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_845) );
INVx1_ASAP7_75t_L g932 ( .A(n_384), .Y(n_932) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_385), .Y(n_1034) );
BUFx6f_ASAP7_75t_L g1517 ( .A(n_385), .Y(n_1517) );
AOI222xp33_ASAP7_75t_L g1563 ( .A1(n_385), .A2(n_1564), .B1(n_1565), .B2(n_1568), .C1(n_1569), .C2(n_1570), .Y(n_1563) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g483 ( .A(n_386), .Y(n_483) );
BUFx3_ASAP7_75t_L g559 ( .A(n_386), .Y(n_559) );
BUFx3_ASAP7_75t_L g635 ( .A(n_386), .Y(n_635) );
BUFx6f_ASAP7_75t_L g1131 ( .A(n_386), .Y(n_1131) );
AND2x4_ASAP7_75t_L g1578 ( .A(n_386), .B(n_1579), .Y(n_1578) );
AOI21xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_464), .B(n_468), .Y(n_388) );
NAND4xp25_ASAP7_75t_SL g389 ( .A(n_390), .B(n_416), .C(n_438), .D(n_447), .Y(n_389) );
AOI222xp33_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_404), .B1(n_405), .B2(n_411), .C1(n_412), .C2(n_415), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_391), .A2(n_1177), .B1(n_1204), .B2(n_1206), .Y(n_1203) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g575 ( .A(n_393), .B(n_510), .Y(n_575) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .Y(n_393) );
AND2x4_ASAP7_75t_L g407 ( .A(n_394), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g412 ( .A(n_394), .B(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
AND2x4_ASAP7_75t_L g601 ( .A(n_394), .B(n_408), .Y(n_601) );
INVx1_ASAP7_75t_L g985 ( .A(n_394), .Y(n_985) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_394), .B(n_413), .Y(n_1042) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g463 ( .A(n_397), .B(n_446), .Y(n_463) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g1591 ( .A(n_398), .Y(n_1591) );
HB1xp67_ASAP7_75t_L g1596 ( .A(n_398), .Y(n_1596) );
INVx1_ASAP7_75t_L g1607 ( .A(n_398), .Y(n_1607) );
INVx6_ASAP7_75t_L g461 ( .A(n_399), .Y(n_461) );
INVx2_ASAP7_75t_L g599 ( .A(n_399), .Y(n_599) );
BUFx2_ASAP7_75t_L g694 ( .A(n_399), .Y(n_694) );
AND2x4_ASAP7_75t_L g1603 ( .A(n_399), .B(n_1595), .Y(n_1603) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g414 ( .A(n_400), .Y(n_414) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g420 ( .A(n_401), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g435 ( .A(n_401), .B(n_403), .Y(n_435) );
INVx1_ASAP7_75t_L g410 ( .A(n_402), .Y(n_410) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g430 ( .A(n_403), .B(n_426), .Y(n_430) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx4_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g685 ( .A(n_407), .Y(n_685) );
INVx1_ASAP7_75t_SL g840 ( .A(n_407), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_407), .A2(n_412), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI222xp33_ASAP7_75t_L g1192 ( .A1(n_407), .A2(n_412), .B1(n_431), .B2(n_1170), .C1(n_1171), .C2(n_1193), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g1161 ( .A1(n_408), .A2(n_413), .B1(n_1162), .B2(n_1163), .Y(n_1161) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g514 ( .A(n_409), .Y(n_514) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g1598 ( .A(n_410), .Y(n_1598) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_411), .A2(n_479), .B(n_482), .Y(n_478) );
AOI322xp5_ASAP7_75t_L g594 ( .A1(n_412), .A2(n_595), .A3(n_596), .B1(n_597), .B2(n_601), .C1(n_602), .C2(n_603), .Y(n_594) );
INVx2_ASAP7_75t_L g684 ( .A(n_412), .Y(n_684) );
INVx2_ASAP7_75t_SL g841 ( .A(n_412), .Y(n_841) );
INVx2_ASAP7_75t_L g520 ( .A(n_413), .Y(n_520) );
BUFx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x6_ASAP7_75t_L g1599 ( .A(n_414), .B(n_1591), .Y(n_1599) );
OR2x2_ASAP7_75t_L g580 ( .A(n_418), .B(n_579), .Y(n_580) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx4f_ASAP7_75t_L g692 ( .A(n_419), .Y(n_692) );
AND2x2_ASAP7_75t_L g832 ( .A(n_419), .B(n_431), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_419), .A2(n_434), .B1(n_1190), .B2(n_1195), .Y(n_1194) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_420), .Y(n_441) );
INVx2_ASAP7_75t_SL g495 ( .A(n_420), .Y(n_495) );
BUFx3_ASAP7_75t_L g506 ( .A(n_420), .Y(n_506) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_420), .Y(n_622) );
BUFx2_ASAP7_75t_L g682 ( .A(n_420), .Y(n_682) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_420), .Y(n_790) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_420), .Y(n_836) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_420), .Y(n_996) );
AND2x6_ASAP7_75t_L g1612 ( .A(n_420), .B(n_1590), .Y(n_1612) );
INVx1_ASAP7_75t_L g427 ( .A(n_421), .Y(n_427) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g578 ( .A(n_424), .Y(n_578) );
OR2x2_ASAP7_75t_L g615 ( .A(n_424), .B(n_432), .Y(n_615) );
INVx1_ASAP7_75t_L g1150 ( .A(n_424), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1609 ( .A(n_424), .B(n_1610), .Y(n_1609) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
AND2x2_ASAP7_75t_L g585 ( .A(n_425), .B(n_427), .Y(n_585) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g1078 ( .A(n_428), .Y(n_1078) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g439 ( .A(n_429), .Y(n_439) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_429), .Y(n_496) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_429), .Y(n_830) );
INVx1_ASAP7_75t_L g838 ( .A(n_429), .Y(n_838) );
BUFx6f_ASAP7_75t_L g1207 ( .A(n_429), .Y(n_1207) );
AND2x6_ASAP7_75t_L g1605 ( .A(n_429), .B(n_1606), .Y(n_1605) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
INVx1_ASAP7_75t_L g508 ( .A(n_430), .Y(n_508) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_430), .Y(n_792) );
AND2x4_ASAP7_75t_L g433 ( .A(n_431), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g621 ( .A(n_431), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g618 ( .A(n_432), .B(n_455), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_433), .A2(n_436), .B1(n_605), .B2(n_606), .C(n_610), .Y(n_604) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_433), .Y(n_687) );
INVx2_ASAP7_75t_SL g826 ( .A(n_433), .Y(n_826) );
BUFx6f_ASAP7_75t_L g973 ( .A(n_433), .Y(n_973) );
AND2x4_ASAP7_75t_L g436 ( .A(n_434), .B(n_437), .Y(n_436) );
BUFx4f_ASAP7_75t_L g442 ( .A(n_434), .Y(n_442) );
INVx1_ASAP7_75t_L g459 ( .A(n_434), .Y(n_459) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
INVx1_ASAP7_75t_L g691 ( .A(n_434), .Y(n_691) );
INVx2_ASAP7_75t_SL g797 ( .A(n_434), .Y(n_797) );
BUFx3_ASAP7_75t_L g802 ( .A(n_434), .Y(n_802) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_435), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_436), .A2(n_687), .B1(n_688), .B2(n_689), .C(n_693), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_436), .A2(n_825), .B1(n_827), .B2(n_828), .C(n_829), .Y(n_824) );
INVx1_ASAP7_75t_L g892 ( .A(n_436), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g1196 ( .A1(n_436), .A2(n_1197), .B(n_1200), .Y(n_1196) );
BUFx3_ASAP7_75t_L g1164 ( .A(n_437), .Y(n_1164) );
BUFx3_ASAP7_75t_L g449 ( .A(n_441), .Y(n_449) );
INVx2_ASAP7_75t_L g1052 ( .A(n_441), .Y(n_1052) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g1199 ( .A(n_444), .Y(n_1199) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
INVx2_ASAP7_75t_L g609 ( .A(n_445), .Y(n_609) );
INVx2_ASAP7_75t_SL g891 ( .A(n_445), .Y(n_891) );
INVx1_ASAP7_75t_L g1532 ( .A(n_445), .Y(n_1532) );
INVx1_ASAP7_75t_L g1616 ( .A(n_446), .Y(n_1616) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B1(n_451), .B2(n_456), .C(n_457), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g611 ( .A(n_455), .Y(n_611) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g980 ( .A(n_459), .Y(n_980) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_461), .Y(n_501) );
INVx2_ASAP7_75t_L g795 ( .A(n_461), .Y(n_795) );
INVx2_ASAP7_75t_L g801 ( .A(n_461), .Y(n_801) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_461), .Y(n_1047) );
INVx1_ASAP7_75t_L g1535 ( .A(n_461), .Y(n_1535) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g509 ( .A(n_463), .B(n_510), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_463), .Y(n_600) );
INVx2_ASAP7_75t_SL g680 ( .A(n_463), .Y(n_680) );
AND2x4_ASAP7_75t_L g808 ( .A(n_463), .B(n_510), .Y(n_808) );
INVx2_ASAP7_75t_L g1001 ( .A(n_463), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_463), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_464), .A2(n_674), .B1(n_698), .B2(n_699), .Y(n_673) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI31xp33_ASAP7_75t_L g1241 ( .A1(n_465), .A2(n_1242), .A3(n_1253), .B(n_1262), .Y(n_1241) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_466), .A2(n_527), .B(n_550), .Y(n_526) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g1116 ( .A(n_467), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1615 ( .A(n_467), .B(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_470), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_470), .A2(n_927), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_470), .A2(n_708), .B1(n_946), .B2(n_947), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_470), .A2(n_708), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_470), .A2(n_708), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1507 ( .A1(n_470), .A2(n_928), .B1(n_1508), .B2(n_1509), .Y(n_1507) );
BUFx2_ASAP7_75t_L g910 ( .A(n_471), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_471), .A2(n_483), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
BUFx3_ASAP7_75t_L g1233 ( .A(n_471), .Y(n_1233) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g541 ( .A(n_472), .Y(n_541) );
INVx2_ASAP7_75t_L g572 ( .A(n_472), .Y(n_572) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_473), .Y(n_557) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_475), .A2(n_634), .B1(n_943), .B2(n_944), .Y(n_942) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g632 ( .A(n_476), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_476), .A2(n_634), .B1(n_703), .B2(n_704), .Y(n_702) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_476), .Y(n_1014) );
BUFx2_ASAP7_75t_L g1223 ( .A(n_476), .Y(n_1223) );
BUFx2_ASAP7_75t_L g1505 ( .A(n_476), .Y(n_1505) );
BUFx3_ASAP7_75t_L g669 ( .A(n_477), .Y(n_669) );
INVx2_ASAP7_75t_L g866 ( .A(n_477), .Y(n_866) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_477), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_479), .A2(n_482), .B1(n_896), .B2(n_897), .C(n_923), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_479), .A2(n_482), .B1(n_923), .B2(n_1010), .C(n_1011), .Y(n_1009) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_479), .A2(n_482), .B1(n_923), .B2(n_1170), .C(n_1171), .Y(n_1169) );
INVx1_ASAP7_75t_L g1219 ( .A(n_479), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1497 ( .A1(n_479), .A2(n_1498), .B1(n_1500), .B2(n_1501), .C(n_1502), .Y(n_1497) );
AND2x2_ASAP7_75t_L g761 ( .A(n_480), .B(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g567 ( .A(n_481), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_482), .A2(n_1216), .B1(n_1217), .B2(n_1218), .C(n_1220), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1502 ( .A(n_482), .Y(n_1502) );
INVx1_ASAP7_75t_L g1024 ( .A(n_483), .Y(n_1024) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR4xp75_ASAP7_75t_L g486 ( .A(n_487), .B(n_526), .C(n_573), .D(n_581), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_511), .Y(n_487) );
AOI33xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_493), .A3(n_497), .B1(n_499), .B2(n_505), .B3(n_509), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
BUFx2_ASAP7_75t_L g624 ( .A(n_491), .Y(n_624) );
INVx2_ASAP7_75t_L g769 ( .A(n_491), .Y(n_769) );
OR2x6_ASAP7_75t_L g787 ( .A(n_491), .B(n_609), .Y(n_787) );
AND2x4_ASAP7_75t_L g908 ( .A(n_491), .B(n_743), .Y(n_908) );
AND2x2_ASAP7_75t_L g921 ( .A(n_491), .B(n_561), .Y(n_921) );
AND2x4_ASAP7_75t_L g1231 ( .A(n_491), .B(n_743), .Y(n_1231) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g781 ( .A(n_495), .Y(n_781) );
INVx1_ASAP7_75t_L g979 ( .A(n_495), .Y(n_979) );
INVx2_ASAP7_75t_SL g977 ( .A(n_496), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_498), .B(n_525), .Y(n_811) );
INVx1_ASAP7_75t_L g999 ( .A(n_498), .Y(n_999) );
INVx1_ASAP7_75t_L g1257 ( .A(n_498), .Y(n_1257) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g678 ( .A(n_501), .Y(n_678) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g679 ( .A(n_503), .Y(n_679) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g524 ( .A(n_504), .Y(n_524) );
BUFx6f_ASAP7_75t_L g986 ( .A(n_504), .Y(n_986) );
BUFx6f_ASAP7_75t_L g1205 ( .A(n_504), .Y(n_1205) );
AND2x4_ASAP7_75t_L g1588 ( .A(n_504), .B(n_1589), .Y(n_1588) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_507), .Y(n_1056) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_579), .Y(n_582) );
OR2x6_ASAP7_75t_L g775 ( .A(n_508), .B(n_579), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_517), .B1(n_518), .B2(n_521), .C(n_522), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g784 ( .A(n_513), .Y(n_784) );
INVx1_ASAP7_75t_L g1083 ( .A(n_513), .Y(n_1083) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OR2x6_ASAP7_75t_L g519 ( .A(n_516), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g525 ( .A(n_516), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_518), .A2(n_760), .B1(n_763), .B2(n_784), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g1081 ( .A1(n_518), .A2(n_522), .B1(n_1082), .B2(n_1083), .C(n_1084), .Y(n_1081) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g992 ( .A(n_520), .B(n_985), .Y(n_992) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_523), .Y(n_1053) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI221x1_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_533), .B1(n_534), .B2(n_535), .C(n_536), .Y(n_527) );
INVx3_ASAP7_75t_L g730 ( .A(n_528), .Y(n_730) );
INVx3_ASAP7_75t_L g1087 ( .A(n_528), .Y(n_1087) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
AND2x4_ASAP7_75t_L g562 ( .A(n_529), .B(n_559), .Y(n_562) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g545 ( .A(n_531), .Y(n_545) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g652 ( .A(n_532), .Y(n_652) );
INVx3_ASAP7_75t_L g729 ( .A(n_534), .Y(n_729) );
INVx3_ASAP7_75t_L g1115 ( .A(n_534), .Y(n_1115) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_542), .B(n_547), .Y(n_536) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_539), .B(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g968 ( .A(n_538), .Y(n_968) );
AOI21xp33_ASAP7_75t_L g1112 ( .A1(n_538), .A2(n_548), .B(n_1113), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_541), .B(n_762), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_542) );
INVx2_ASAP7_75t_L g716 ( .A(n_543), .Y(n_716) );
INVx1_ASAP7_75t_L g917 ( .A(n_545), .Y(n_917) );
INVx1_ASAP7_75t_L g568 ( .A(n_548), .Y(n_568) );
INVx1_ASAP7_75t_L g762 ( .A(n_548), .Y(n_762) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI221xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_555), .B1(n_562), .B2(n_563), .C(n_564), .Y(n_550) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g963 ( .A(n_554), .Y(n_963) );
INVx2_ASAP7_75t_L g1104 ( .A(n_554), .Y(n_1104) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g920 ( .A(n_557), .Y(n_920) );
BUFx6f_ASAP7_75t_L g1022 ( .A(n_557), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1512 ( .A(n_558), .Y(n_1512) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g751 ( .A(n_560), .Y(n_751) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx8_ASAP7_75t_L g745 ( .A(n_562), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
CKINVDCx11_ASAP7_75t_R g764 ( .A(n_569), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x6_ASAP7_75t_L g767 ( .A(n_575), .B(n_768), .Y(n_767) );
AOI222xp33_ASAP7_75t_L g1117 ( .A1(n_575), .A2(n_774), .B1(n_778), .B2(n_1105), .C1(n_1108), .C2(n_1111), .Y(n_1117) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g883 ( .A(n_578), .Y(n_883) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_578), .Y(n_976) );
INVx2_ASAP7_75t_L g1251 ( .A(n_578), .Y(n_1251) );
OR2x6_ASAP7_75t_L g583 ( .A(n_579), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g779 ( .A(n_579), .Y(n_779) );
CKINVDCx6p67_ASAP7_75t_R g776 ( .A(n_583), .Y(n_776) );
OAI21xp33_ASAP7_75t_L g1144 ( .A1(n_584), .A2(n_1145), .B(n_1146), .Y(n_1144) );
OAI221xp5_ASAP7_75t_L g1250 ( .A1(n_584), .A2(n_1224), .B1(n_1226), .B2(n_1251), .C(n_1252), .Y(n_1250) );
INVx1_ASAP7_75t_L g1586 ( .A(n_584), .Y(n_1586) );
BUFx3_ASAP7_75t_L g1635 ( .A(n_584), .Y(n_1635) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx4f_ASAP7_75t_L g889 ( .A(n_585), .Y(n_889) );
INVx1_ASAP7_75t_L g1154 ( .A(n_585), .Y(n_1154) );
INVx1_ASAP7_75t_L g1160 ( .A(n_585), .Y(n_1160) );
BUFx2_ASAP7_75t_L g1528 ( .A(n_585), .Y(n_1528) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
XNOR2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g1389 ( .A1(n_590), .A2(n_1390), .B1(n_1391), .B2(n_1392), .Y(n_1389) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_628), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_623), .B1(n_625), .B2(n_626), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_604), .C(n_612), .D(n_619), .Y(n_593) );
AND2x2_ASAP7_75t_L g778 ( .A(n_598), .B(n_779), .Y(n_778) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_598), .Y(n_1072) );
A2O1A1Ixp33_ASAP7_75t_L g1157 ( .A1(n_598), .A2(n_1158), .B(n_1159), .C(n_1164), .Y(n_1157) );
INVx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g1261 ( .A(n_599), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_601), .A2(n_990), .B1(n_991), .B2(n_993), .Y(n_989) );
INVx2_ASAP7_75t_L g1245 ( .A(n_601), .Y(n_1245) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_605), .A2(n_613), .B1(n_664), .B2(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g1151 ( .A(n_611), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_616), .B2(n_617), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_614), .A2(n_617), .B1(n_696), .B2(n_697), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_614), .A2(n_617), .B1(n_822), .B2(n_823), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_614), .A2(n_617), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_614), .A2(n_617), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_614), .A2(n_617), .B1(n_1538), .B2(n_1539), .Y(n_1537) );
INVx6_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_616), .A2(n_620), .B1(n_647), .B2(n_668), .Y(n_667) );
INVx4_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_621), .A2(n_676), .B1(n_677), .B2(n_681), .C(n_683), .Y(n_675) );
INVx1_ASAP7_75t_L g988 ( .A(n_621), .Y(n_988) );
AOI21xp33_ASAP7_75t_SL g1038 ( .A1(n_621), .A2(n_1039), .B(n_1040), .Y(n_1038) );
AOI211xp5_ASAP7_75t_L g1242 ( .A1(n_621), .A2(n_1243), .B(n_1244), .C(n_1246), .Y(n_1242) );
AOI211xp5_ASAP7_75t_L g1522 ( .A1(n_621), .A2(n_1523), .B(n_1524), .C(n_1525), .Y(n_1522) );
BUFx3_ASAP7_75t_L g804 ( .A(n_622), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_623), .A2(n_626), .B1(n_820), .B2(n_842), .Y(n_819) );
INVx2_ASAP7_75t_L g1060 ( .A(n_623), .Y(n_1060) );
CKINVDCx8_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
OAI31xp33_ASAP7_75t_L g727 ( .A1(n_624), .A2(n_728), .A3(n_731), .B(n_744), .Y(n_727) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g699 ( .A(n_627), .Y(n_699) );
INVx5_ASAP7_75t_L g939 ( .A(n_627), .Y(n_939) );
INVx1_ASAP7_75t_L g1519 ( .A(n_627), .Y(n_1519) );
NOR3xp33_ASAP7_75t_SL g628 ( .A(n_629), .B(n_639), .C(n_645), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_636), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_634), .A2(n_1013), .B1(n_1014), .B2(n_1015), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_634), .A2(n_1222), .B1(n_1223), .B2(n_1224), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_634), .A2(n_1504), .B1(n_1505), .B2(n_1506), .Y(n_1503) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g854 ( .A(n_641), .Y(n_854) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g949 ( .A(n_644), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B1(n_651), .B2(n_653), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g755 ( .A(n_649), .Y(n_755) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_649), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_651), .A2(n_715), .B1(n_717), .B2(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g871 ( .A(n_652), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_SL g664 ( .A(n_656), .Y(n_664) );
INVx1_ASAP7_75t_L g1096 ( .A(n_656), .Y(n_1096) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
BUFx3_ASAP7_75t_L g958 ( .A(n_659), .Y(n_958) );
INVx1_ASAP7_75t_L g1632 ( .A(n_661), .Y(n_1632) );
CKINVDCx8_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g747 ( .A(n_666), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_668), .A2(n_676), .B1(n_697), .B2(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_723), .B1(n_724), .B2(n_813), .Y(n_670) );
INVx2_ASAP7_75t_L g813 ( .A(n_671), .Y(n_813) );
XOR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_722), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_700), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_686), .C(n_695), .Y(n_674) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_709), .C(n_710), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_716), .Y(n_720) );
INVx2_ASAP7_75t_L g735 ( .A(n_716), .Y(n_735) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND3xp33_ASAP7_75t_SL g726 ( .A(n_727), .B(n_765), .C(n_771), .Y(n_726) );
CKINVDCx6p67_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_734) );
BUFx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g1099 ( .A(n_743), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_749), .B2(n_750), .C(n_751), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_748), .A2(n_758), .B1(n_774), .B2(n_776), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_750), .A2(n_756), .B1(n_778), .B2(n_780), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g1126 ( .A1(n_755), .A2(n_1127), .B1(n_1128), .B2(n_1129), .C(n_1130), .Y(n_1126) );
INVx1_ASAP7_75t_L g1236 ( .A(n_757), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_763), .B2(n_764), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
NOR2xp67_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx2_ASAP7_75t_L g905 ( .A(n_769), .Y(n_905) );
INVx1_ASAP7_75t_L g1110 ( .A(n_770), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_782), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_777), .Y(n_772) );
CKINVDCx6p67_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_776), .A2(n_780), .B1(n_1102), .B2(n_1107), .Y(n_1118) );
AND2x2_ASAP7_75t_L g780 ( .A(n_779), .B(n_781), .Y(n_780) );
NAND3xp33_ASAP7_75t_SL g782 ( .A(n_783), .B(n_785), .C(n_809), .Y(n_782) );
AOI33xp33_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .A3(n_793), .B1(n_798), .B2(n_803), .B3(n_807), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g1069 ( .A(n_787), .Y(n_1069) );
OAI22xp5_ASAP7_75t_SL g1633 ( .A1(n_787), .A2(n_1080), .B1(n_1634), .B2(n_1637), .Y(n_1633) );
BUFx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_790), .Y(n_1077) );
INVx1_ASAP7_75t_L g1248 ( .A(n_790), .Y(n_1248) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g806 ( .A(n_792), .Y(n_806) );
BUFx3_ASAP7_75t_L g1249 ( .A(n_792), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_795), .Y(n_1055) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g1198 ( .A(n_797), .Y(n_1198) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx6f_ASAP7_75t_L g1201 ( .A(n_801), .Y(n_1201) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_806), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
BUFx4f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx4_ASAP7_75t_L g1080 ( .A(n_808), .Y(n_1080) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_SL g1267 ( .A(n_814), .Y(n_1267) );
XNOR2x1_ASAP7_75t_L g814 ( .A(n_815), .B(n_1063), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_935), .Y(n_815) );
XOR2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_877), .Y(n_816) );
INVx1_ASAP7_75t_L g875 ( .A(n_818), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_843), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_831), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_822), .A2(n_827), .B1(n_873), .B2(n_874), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_823), .A2(n_833), .B1(n_869), .B2(n_871), .Y(n_868) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AOI221xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_834), .B2(n_835), .C(n_839), .Y(n_831) );
INVx1_ASAP7_75t_L g894 ( .A(n_832), .Y(n_894) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g1202 ( .A(n_838), .Y(n_1202) );
NOR3xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_852), .C(n_855), .Y(n_843) );
NAND2xp5_ASAP7_75t_SL g844 ( .A(n_845), .B(n_849), .Y(n_844) );
INVx2_ASAP7_75t_L g931 ( .A(n_847), .Y(n_931) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_859), .B1(n_860), .B2(n_862), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_864), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1089) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OAI22xp33_ASAP7_75t_L g956 ( .A1(n_873), .A2(n_957), .B1(n_958), .B2(n_959), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_873), .A2(n_966), .B1(n_967), .B2(n_969), .Y(n_965) );
INVx1_ASAP7_75t_L g934 ( .A(n_878), .Y(n_934) );
NAND4xp75_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .C(n_906), .D(n_926), .Y(n_878) );
OAI31xp33_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_893), .A3(n_903), .B(n_904), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g1634 ( .A1(n_883), .A2(n_1621), .B1(n_1622), .B2(n_1635), .C(n_1636), .Y(n_1634) );
OAI21xp33_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B(n_890), .Y(n_886) );
INVx2_ASAP7_75t_SL g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g900 ( .A(n_889), .Y(n_900) );
INVx2_ASAP7_75t_L g1044 ( .A(n_889), .Y(n_1044) );
BUFx2_ASAP7_75t_L g981 ( .A(n_891), .Y(n_981) );
INVx1_ASAP7_75t_L g1259 ( .A(n_891), .Y(n_1259) );
OAI211xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .B(n_901), .C(n_902), .Y(n_898) );
OAI31xp33_ASAP7_75t_L g970 ( .A1(n_904), .A2(n_971), .A3(n_987), .B(n_1002), .Y(n_970) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
AOI31xp33_ASAP7_75t_SL g1191 ( .A1(n_905), .A2(n_1192), .A3(n_1196), .B(n_1203), .Y(n_1191) );
AND2x2_ASAP7_75t_SL g906 ( .A(n_907), .B(n_922), .Y(n_906) );
AOI33xp33_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .A3(n_911), .B1(n_916), .B2(n_918), .B3(n_921), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g1172 ( .A1(n_908), .A2(n_1173), .B1(n_1177), .B2(n_1178), .Y(n_1172) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g1132 ( .A(n_921), .B(n_1133), .C(n_1134), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_923), .Y(n_1216) );
INVx1_ASAP7_75t_L g1499 ( .A(n_923), .Y(n_1499) );
AND2x4_ASAP7_75t_L g1565 ( .A(n_924), .B(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_1005), .B1(n_1006), .B2(n_1062), .Y(n_935) );
INVx1_ASAP7_75t_L g1062 ( .A(n_936), .Y(n_1062) );
INVx1_ASAP7_75t_L g1003 ( .A(n_937), .Y(n_1003) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_939), .A2(n_1036), .B(n_1037), .Y(n_1035) );
AOI21xp5_ASAP7_75t_L g1239 ( .A1(n_939), .A2(n_1240), .B(n_1241), .Y(n_1239) );
NOR3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_948), .C(n_950), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_945), .Y(n_941) );
OAI221xp5_ASAP7_75t_L g994 ( .A1(n_943), .A2(n_947), .B1(n_977), .B2(n_995), .C(n_997), .Y(n_994) );
INVx2_ASAP7_75t_SL g953 ( .A(n_954), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g974 ( .A1(n_955), .A2(n_957), .B1(n_975), .B2(n_977), .C(n_978), .Y(n_974) );
OAI22xp33_ASAP7_75t_SL g1627 ( .A1(n_958), .A2(n_1628), .B1(n_1629), .B2(n_1631), .Y(n_1627) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_973), .A2(n_983), .B1(n_1049), .B2(n_1050), .C(n_1054), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_973), .A2(n_983), .B1(n_1254), .B2(n_1255), .C(n_1260), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1530 ( .A1(n_973), .A2(n_983), .B1(n_1531), .B2(n_1533), .C(n_1536), .Y(n_1530) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
AND2x4_ASAP7_75t_L g983 ( .A(n_984), .B(n_986), .Y(n_983) );
INVx1_ASAP7_75t_SL g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1074 ( .A(n_986), .Y(n_1074) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1001), .Y(n_1529) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_1006), .Y(n_1005) );
XNOR2x1_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1061), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1035), .Y(n_1007) );
AND4x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .C(n_1016), .D(n_1019), .Y(n_1008) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_1015), .A2(n_1044), .B(n_1045), .C(n_1046), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1022), .Y(n_1032) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1619 ( .A(n_1026), .Y(n_1619) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
AOI31xp33_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1048), .A3(n_1057), .B(n_1060), .Y(n_1037) );
INVx3_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
AOI31xp33_ASAP7_75t_L g1521 ( .A1(n_1060), .A2(n_1522), .A3(n_1530), .B(n_1537), .Y(n_1521) );
AO22x2_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1212), .B1(n_1265), .B2(n_1266), .Y(n_1063) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1064), .Y(n_1265) );
XNOR2xp5_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1119), .Y(n_1064) );
NAND4xp75_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1085), .C(n_1117), .D(n_1118), .Y(n_1066) );
AND2x2_ASAP7_75t_SL g1067 ( .A(n_1068), .B(n_1081), .Y(n_1067) );
AOI33xp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .A3(n_1071), .B1(n_1075), .B2(n_1076), .B3(n_1079), .Y(n_1068) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1077), .Y(n_1638) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
OAI31xp33_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1088), .A3(n_1114), .B(n_1116), .Y(n_1085) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1093), .B1(n_1100), .B2(n_1106), .C(n_1109), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B1(n_1096), .B2(n_1097), .C(n_1098), .Y(n_1093) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B1(n_1103), .B2(n_1105), .Y(n_1100) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
AOI21xp5_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1111), .B(n_1112), .Y(n_1109) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1116), .Y(n_1165) );
XNOR2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1166), .Y(n_1119) );
NAND3xp33_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1136), .C(n_1140), .Y(n_1121) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1135), .Y(n_1122) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_1129), .A2(n_1148), .B1(n_1149), .B2(n_1151), .Y(n_1147) );
NOR2xp33_ASAP7_75t_SL g1136 ( .A(n_1137), .B(n_1139), .Y(n_1136) );
OAI31xp33_ASAP7_75t_SL g1140 ( .A1(n_1141), .A2(n_1142), .A3(n_1143), .B(n_1165), .Y(n_1140) );
OAI211xp5_ASAP7_75t_SL g1143 ( .A1(n_1144), .A2(n_1147), .B(n_1152), .C(n_1157), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1526 ( .A1(n_1149), .A2(n_1506), .B1(n_1508), .B2(n_1527), .C(n_1529), .Y(n_1526) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
OAI211xp5_ASAP7_75t_L g1152 ( .A1(n_1153), .A2(n_1154), .B(n_1155), .C(n_1156), .Y(n_1152) );
NAND2xp33_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
NAND2xp5_ASAP7_75t_SL g1166 ( .A(n_1167), .B(n_1208), .Y(n_1166) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1168), .Y(n_1210) );
NAND3xp33_ASAP7_75t_SL g1168 ( .A(n_1169), .B(n_1172), .C(n_1179), .Y(n_1168) );
BUFx3_ASAP7_75t_L g1235 ( .A(n_1185), .Y(n_1235) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1191), .Y(n_1209) );
NAND3xp33_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .C(n_1211), .Y(n_1208) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1212), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1239), .Y(n_1213) );
AND4x1_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1221), .C(n_1225), .D(n_1228), .Y(n_1214) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1617 ( .A1(n_1229), .A2(n_1618), .B1(n_1624), .B2(n_1632), .C(n_1633), .Y(n_1617) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_1269), .A2(n_1491), .B1(n_1494), .B2(n_1542), .C(n_1547), .Y(n_1268) );
NOR2xp67_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1429), .Y(n_1269) );
OAI21xp33_ASAP7_75t_L g1270 ( .A1(n_1271), .A2(n_1385), .B(n_1393), .Y(n_1270) );
NOR5xp2_ASAP7_75t_SL g1271 ( .A(n_1272), .B(n_1325), .C(n_1353), .D(n_1365), .E(n_1373), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1300), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_1273), .A2(n_1378), .B1(n_1407), .B2(n_1409), .Y(n_1406) );
OAI211xp5_ASAP7_75t_L g1436 ( .A1(n_1273), .A2(n_1368), .B(n_1437), .C(n_1439), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1273), .B(n_1440), .Y(n_1456) );
HB1xp67_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx2_ASAP7_75t_SL g1348 ( .A(n_1274), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1274), .B(n_1314), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1274), .B(n_1329), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1274), .B(n_1427), .Y(n_1426) );
AND2x4_ASAP7_75t_L g1435 ( .A(n_1274), .B(n_1328), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1444 ( .A(n_1274), .B(n_1427), .Y(n_1444) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1274), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_1274), .B(n_1418), .Y(n_1481) );
CKINVDCx5p33_ASAP7_75t_R g1274 ( .A(n_1275), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1275), .B(n_1328), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1275), .B(n_1329), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1290), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1284), .B1(n_1285), .B2(n_1289), .Y(n_1276) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_1277), .Y(n_1390) );
BUFx6f_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
OAI22xp5_ASAP7_75t_L g1322 ( .A1(n_1278), .A2(n_1287), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1280), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1279), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1279), .Y(n_1307) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1280), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1283), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1283), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g1392 ( .A(n_1285), .Y(n_1392) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1288), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1296), .B1(n_1297), .B2(n_1299), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
BUFx3_ASAP7_75t_L g1388 ( .A(n_1292), .Y(n_1388) );
AND2x4_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1295), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1293), .B(n_1295), .Y(n_1311) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
AND2x4_ASAP7_75t_L g1298 ( .A(n_1294), .B(n_1295), .Y(n_1298) );
INVx2_ASAP7_75t_L g1345 ( .A(n_1297), .Y(n_1345) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1312), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1302), .B(n_1339), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1302), .B(n_1351), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1302), .B(n_1336), .Y(n_1464) );
INVxp67_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
BUFx3_ASAP7_75t_L g1335 ( .A(n_1303), .Y(n_1335) );
BUFx2_ASAP7_75t_L g1350 ( .A(n_1303), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1303), .B(n_1339), .Y(n_1378) );
AOI222xp33_ASAP7_75t_L g1411 ( .A1(n_1303), .A2(n_1349), .B1(n_1364), .B2(n_1380), .C1(n_1412), .C2(n_1413), .Y(n_1411) );
NOR3xp33_ASAP7_75t_L g1466 ( .A(n_1303), .B(n_1367), .C(n_1447), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1310), .Y(n_1303) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1307), .Y(n_1305) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_1307), .B(n_1309), .Y(n_1308) );
BUFx2_ASAP7_75t_L g1343 ( .A(n_1308), .Y(n_1343) );
HB1xp67_ASAP7_75t_L g1643 ( .A(n_1309), .Y(n_1643) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1317), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1313), .B(n_1370), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1313), .B(n_1348), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1313), .B(n_1435), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1313), .B(n_1485), .Y(n_1484) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
BUFx2_ASAP7_75t_L g1332 ( .A(n_1314), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1314), .B(n_1335), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1314), .B(n_1350), .Y(n_1399) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1314), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1314), .B(n_1363), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1316), .Y(n_1314) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1317), .Y(n_1339) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1317), .B(n_1376), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1321), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1318), .B(n_1337), .Y(n_1336) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1318), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1318), .B(n_1335), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1318), .B(n_1321), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1318), .B(n_1335), .Y(n_1382) );
OAI321xp33_ASAP7_75t_L g1442 ( .A1(n_1318), .A2(n_1443), .A3(n_1445), .B1(n_1447), .B2(n_1449), .C(n_1450), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1320), .Y(n_1318) );
INVx2_ASAP7_75t_SL g1337 ( .A(n_1321), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1321), .B(n_1352), .Y(n_1351) );
OAI222xp33_ASAP7_75t_L g1394 ( .A1(n_1321), .A2(n_1328), .B1(n_1395), .B2(n_1397), .C1(n_1400), .C2(n_1401), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1321), .B(n_1335), .Y(n_1485) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1333), .B1(n_1340), .B2(n_1346), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1332), .Y(n_1326) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1327), .Y(n_1441) );
OAI311xp33_ASAP7_75t_L g1462 ( .A1(n_1327), .A2(n_1385), .A3(n_1463), .B1(n_1465), .C1(n_1468), .Y(n_1462) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
NOR2xp33_ASAP7_75t_L g1383 ( .A(n_1328), .B(n_1384), .Y(n_1383) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1328), .B(n_1446), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1328), .B(n_1341), .Y(n_1448) );
INVx3_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1340 ( .A(n_1329), .B(n_1341), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1329), .B(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1329), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
NAND2xp5_ASAP7_75t_SL g1356 ( .A(n_1332), .B(n_1357), .Y(n_1356) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1332), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1332), .B(n_1396), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1332), .B(n_1414), .Y(n_1413) );
AOI221xp5_ASAP7_75t_L g1430 ( .A1(n_1332), .A2(n_1431), .B1(n_1436), .B2(n_1441), .C(n_1442), .Y(n_1430) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1338), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1334), .B(n_1427), .Y(n_1440) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1334), .Y(n_1449) );
OAI21xp5_ASAP7_75t_SL g1468 ( .A1(n_1334), .A2(n_1469), .B(n_1470), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1336), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1335), .B(n_1337), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1335), .B(n_1369), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1335), .B(n_1410), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1454 ( .A(n_1335), .B(n_1352), .Y(n_1454) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1336), .Y(n_1375) );
NAND3xp33_ASAP7_75t_SL g1450 ( .A(n_1336), .B(n_1404), .C(n_1451), .Y(n_1450) );
AOI321xp33_ASAP7_75t_L g1457 ( .A1(n_1337), .A2(n_1348), .A3(n_1370), .B1(n_1458), .B2(n_1459), .C(n_1460), .Y(n_1457) );
NOR2x1_ASAP7_75t_L g1469 ( .A(n_1337), .B(n_1350), .Y(n_1469) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1338), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1339), .B(n_1362), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1339), .B(n_1399), .Y(n_1438) );
NOR2xp33_ASAP7_75t_L g1459 ( .A(n_1340), .B(n_1348), .Y(n_1459) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1340), .Y(n_1482) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1341), .Y(n_1360) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1341), .Y(n_1363) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1341), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1344), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1349), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1407 ( .A(n_1347), .B(n_1408), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1347), .B(n_1438), .Y(n_1437) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1348), .B(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1348), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1473 ( .A(n_1348), .B(n_1474), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1349), .B(n_1367), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_1350), .B(n_1352), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1351), .B(n_1399), .Y(n_1398) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1351), .Y(n_1432) );
A2O1A1Ixp33_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1356), .B(n_1358), .C(n_1361), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1357), .B(n_1367), .Y(n_1401) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
AOI211xp5_ASAP7_75t_L g1472 ( .A1(n_1359), .A2(n_1473), .B(n_1475), .C(n_1487), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1359), .B(n_1480), .Y(n_1486) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1360), .Y(n_1404) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1360), .Y(n_1418) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1362), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1364), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1363), .B(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1363), .Y(n_1424) );
AOI32xp33_ASAP7_75t_L g1465 ( .A1(n_1364), .A2(n_1382), .A3(n_1458), .B1(n_1466), .B2(n_1467), .Y(n_1465) );
AOI21xp33_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1368), .B(n_1371), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1367), .B(n_1396), .Y(n_1400) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1367), .B(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1370), .B(n_1399), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1370), .B(n_1477), .Y(n_1476) );
A2O1A1Ixp33_ASAP7_75t_L g1373 ( .A1(n_1374), .A2(n_1377), .B(n_1379), .C(n_1381), .Y(n_1373) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1376), .Y(n_1374) );
NOR3xp33_ASAP7_75t_L g1460 ( .A(n_1375), .B(n_1424), .C(n_1461), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1375), .B(n_1432), .Y(n_1467) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1376), .Y(n_1477) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1379), .B(n_1421), .Y(n_1420) );
CKINVDCx5p33_ASAP7_75t_R g1379 ( .A(n_1380), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1383), .Y(n_1381) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx3_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1387), .B(n_1403), .Y(n_1402) );
INVx3_ASAP7_75t_L g1417 ( .A(n_1387), .Y(n_1417) );
AOI21xp5_ASAP7_75t_L g1452 ( .A1(n_1387), .A2(n_1453), .B(n_1462), .Y(n_1452) );
O2A1O1Ixp33_ASAP7_75t_L g1478 ( .A1(n_1387), .A2(n_1479), .B(n_1481), .C(n_1482), .Y(n_1478) );
BUFx2_ASAP7_75t_SL g1493 ( .A(n_1392), .Y(n_1493) );
AOI221xp5_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1402), .B1(n_1405), .B2(n_1415), .C(n_1419), .Y(n_1393) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1396), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
OAI222xp33_ASAP7_75t_L g1475 ( .A1(n_1401), .A2(n_1433), .B1(n_1476), .B2(n_1478), .C1(n_1483), .C2(n_1486), .Y(n_1475) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1404), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1411), .Y(n_1405) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
OAI211xp5_ASAP7_75t_L g1429 ( .A1(n_1417), .A2(n_1430), .B(n_1452), .C(n_1472), .Y(n_1429) );
O2A1O1Ixp33_ASAP7_75t_L g1487 ( .A1(n_1417), .A2(n_1474), .B(n_1488), .C(n_1489), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1418), .B(n_1435), .Y(n_1434) );
OAI21xp33_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1422), .B(n_1423), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1425), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1428), .Y(n_1425) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1426), .Y(n_1461) );
NOR2xp33_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1433), .Y(n_1431) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
OAI211xp5_ASAP7_75t_L g1453 ( .A1(n_1454), .A2(n_1455), .B(n_1456), .C(n_1457), .Y(n_1453) );
INVx2_ASAP7_75t_L g1490 ( .A(n_1464), .Y(n_1490) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
CKINVDCx5p33_ASAP7_75t_R g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_SL g1492 ( .A(n_1493), .Y(n_1492) );
INVx2_ASAP7_75t_L g1541 ( .A(n_1495), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1518), .Y(n_1495) );
AND4x1_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1503), .C(n_1507), .D(n_1510), .Y(n_1496) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
AOI21xp33_ASAP7_75t_SL g1518 ( .A1(n_1519), .A2(n_1520), .B(n_1521), .Y(n_1518) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
HB1xp67_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
CKINVDCx14_ASAP7_75t_R g1542 ( .A(n_1543), .Y(n_1542) );
INVx2_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
CKINVDCx5p33_ASAP7_75t_R g1544 ( .A(n_1545), .Y(n_1544) );
OAI21xp5_ASAP7_75t_L g1642 ( .A1(n_1546), .A2(n_1643), .B(n_1644), .Y(n_1642) );
BUFx2_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx2_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1617), .Y(n_1552) );
O2A1O1Ixp33_ASAP7_75t_L g1553 ( .A1(n_1554), .A2(n_1562), .B(n_1580), .C(n_1582), .Y(n_1553) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
AND2x4_ASAP7_75t_L g1559 ( .A(n_1557), .B(n_1560), .Y(n_1559) );
INVx5_ASAP7_75t_SL g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
NAND3xp33_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1571), .C(n_1577), .Y(n_1562) );
AOI22xp33_ASAP7_75t_L g1592 ( .A1(n_1564), .A2(n_1569), .B1(n_1593), .B2(n_1599), .Y(n_1592) );
INVxp67_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1567), .Y(n_1579) );
OAI221xp5_ASAP7_75t_L g1637 ( .A1(n_1568), .A2(n_1635), .B1(n_1638), .B2(n_1639), .C(n_1640), .Y(n_1637) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_1572), .A2(n_1573), .B1(n_1574), .B2(n_1575), .Y(n_1571) );
INVx5_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
CKINVDCx11_ASAP7_75t_R g1577 ( .A(n_1578), .Y(n_1577) );
CKINVDCx16_ASAP7_75t_R g1580 ( .A(n_1581), .Y(n_1580) );
AOI21xp5_ASAP7_75t_L g1582 ( .A1(n_1583), .A2(n_1600), .B(n_1613), .Y(n_1582) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
INVx2_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
CKINVDCx8_ASAP7_75t_R g1587 ( .A(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1590), .Y(n_1610) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
BUFx4f_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
AND2x4_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1597), .Y(n_1594) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
NOR2xp33_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1608), .Y(n_1600) );
INVx4_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx4_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_SL g1606 ( .A(n_1607), .Y(n_1606) );
CKINVDCx6p67_ASAP7_75t_R g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
BUFx6f_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx3_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
endmodule