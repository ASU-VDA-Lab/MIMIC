module fake_netlist_6_3825_n_1247 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1247);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1247;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_50),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_8),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_177),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_87),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_28),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_62),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_64),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_44),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_86),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_34),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_135),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_51),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_70),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_24),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_22),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_37),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_13),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_164),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_132),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_81),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_78),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_48),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_73),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_28),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_66),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_47),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_75),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_109),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_33),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_236),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_179),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_212),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_218),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_184),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_220),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_184),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_183),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_192),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_183),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_200),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_214),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_239),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_242),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_246),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_249),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_250),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_251),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

BUFx8_ASAP7_75t_SL g298 ( 
.A(n_248),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_254),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_265),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_259),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_255),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_261),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_240),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_241),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_239),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_237),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_310),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_292),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_309),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_273),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_273),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_309),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_295),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_273),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_267),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_311),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_299),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_313),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_274),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_314),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_302),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_287),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_305),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_289),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_275),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_275),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_291),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_303),
.Y(n_370)
);

CKINVDCx6p67_ASAP7_75t_R g371 ( 
.A(n_356),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_313),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_303),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_303),
.Y(n_378)
);

BUFx12f_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_340),
.B(n_303),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_303),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_329),
.B(n_199),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_286),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_364),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_334),
.B(n_300),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_320),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_344),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_303),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

BUFx12f_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_300),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_288),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_324),
.B(n_301),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_271),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_325),
.B(n_301),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_326),
.B(n_306),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_367),
.B(n_284),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_330),
.B(n_306),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

BUFx8_ASAP7_75t_SL g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_403),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_307),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_413),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_332),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_393),
.A2(n_331),
.B1(n_327),
.B2(n_357),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_348),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

CKINVDCx11_ASAP7_75t_R g428 ( 
.A(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_384),
.A2(n_359),
.B(n_348),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_412),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_403),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_408),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_393),
.Y(n_440)
);

AOI22x1_ASAP7_75t_SL g441 ( 
.A1(n_371),
.A2(n_365),
.B1(n_360),
.B2(n_331),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_359),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_307),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_335),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_335),
.Y(n_445)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_375),
.B(n_215),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_406),
.A2(n_327),
.B1(n_368),
.B2(n_358),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_363),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_363),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_345),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_345),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_392),
.B(n_366),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_409),
.A2(n_358),
.B1(n_368),
.B2(n_323),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_366),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_293),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_392),
.A2(n_194),
.B1(n_191),
.B2(n_196),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_411),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

BUFx12f_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_375),
.B(n_293),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

AND2x2_ASAP7_75t_SL g471 ( 
.A(n_375),
.B(n_215),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_397),
.B(n_294),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_391),
.B(n_304),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_382),
.B(n_181),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_382),
.B(n_182),
.Y(n_476)
);

OA21x2_ASAP7_75t_L g477 ( 
.A1(n_378),
.A2(n_312),
.B(n_276),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_397),
.B(n_294),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_382),
.B(n_189),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_382),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

AND3x2_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_204),
.C(n_193),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_386),
.A2(n_230),
.B1(n_206),
.B2(n_208),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_373),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_399),
.B(n_210),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_394),
.A2(n_198),
.B1(n_188),
.B2(n_232),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_373),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_394),
.B(n_203),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_373),
.B(n_213),
.Y(n_494)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_385),
.A2(n_312),
.B(n_276),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_377),
.B(n_397),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_397),
.B(n_296),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_396),
.B(n_217),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_370),
.A2(n_318),
.B(n_226),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_376),
.A2(n_198),
.B1(n_222),
.B2(n_229),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_388),
.B(n_296),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_459),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_398),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_430),
.A2(n_235),
.B(n_233),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_417),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_410),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_428),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_428),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_420),
.B(n_410),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_439),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_419),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_497),
.A2(n_318),
.B(n_316),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_455),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_420),
.B(n_377),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_440),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_420),
.B(n_377),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_417),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_441),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_445),
.B(n_362),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_452),
.B(n_279),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_423),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_458),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_427),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_415),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_462),
.B(n_377),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_459),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_442),
.B(n_388),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_464),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_433),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_464),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_R g552 ( 
.A(n_495),
.B(n_433),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_451),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_462),
.B(n_388),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_450),
.B(n_388),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_466),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_473),
.B(n_185),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_451),
.B(n_388),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_418),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_466),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_447),
.Y(n_562)
);

CKINVDCx6p67_ASAP7_75t_R g563 ( 
.A(n_453),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_460),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_416),
.B(n_388),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_459),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_473),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_488),
.B(n_390),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_567),
.B(n_474),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_505),
.B(n_446),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_523),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_538),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_511),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_511),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_512),
.B(n_474),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_559),
.B(n_446),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_454),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_516),
.Y(n_580)
);

INVxp33_ASAP7_75t_SL g581 ( 
.A(n_510),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_536),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_489),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_536),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_529),
.B(n_471),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_537),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_541),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_542),
.A2(n_456),
.B1(n_493),
.B2(n_499),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_516),
.B(n_461),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_515),
.B(n_471),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_541),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_503),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_557),
.B(n_499),
.C(n_484),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_515),
.B(n_472),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_515),
.B(n_472),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_528),
.B(n_460),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_546),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_563),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_549),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_539),
.B(n_544),
.Y(n_605)
);

AO22x2_ASAP7_75t_L g606 ( 
.A1(n_518),
.A2(n_497),
.B1(n_490),
.B2(n_434),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_506),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

HB1xp67_ASAP7_75t_SL g609 ( 
.A(n_510),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_580),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_599),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_594),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_576),
.B(n_563),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_600),
.B(n_605),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_578),
.B(n_554),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_594),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_573),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_484),
.C(n_485),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_592),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_590),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_599),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_571),
.B(n_523),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_594),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_579),
.B(n_548),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_574),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_579),
.B(n_525),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_571),
.B(n_562),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_583),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_586),
.A2(n_531),
.B1(n_532),
.B2(n_530),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_594),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_601),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_601),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_533),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_596),
.A2(n_569),
.B1(n_564),
.B2(n_478),
.Y(n_635)
);

BUFx8_ASAP7_75t_SL g636 ( 
.A(n_609),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_575),
.B(n_535),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_573),
.B(n_562),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_577),
.B(n_553),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_575),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_591),
.A2(n_498),
.B1(n_469),
.B2(n_472),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_592),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_570),
.B(n_526),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_582),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_581),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_603),
.B(n_487),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_584),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_572),
.Y(n_651)
);

BUFx4f_ASAP7_75t_L g652 ( 
.A(n_572),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_597),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_608),
.B(n_435),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_584),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_526),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_608),
.B(n_435),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_605),
.B(n_517),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_585),
.B(n_469),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_577),
.B(n_495),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_592),
.B(n_522),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_594),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_592),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_577),
.B(n_540),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_585),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_594),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_587),
.B(n_469),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_588),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_589),
.B(n_565),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_608),
.B(n_522),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_588),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_588),
.B(n_522),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_593),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_593),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_593),
.B(n_434),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_592),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_595),
.B(n_438),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_595),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_592),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_595),
.B(n_438),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_589),
.A2(n_476),
.B1(n_481),
.B2(n_475),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_577),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_602),
.B(n_506),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_607),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_607),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_607),
.A2(n_520),
.B1(n_517),
.B2(n_556),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_607),
.B(n_520),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_602),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_602),
.B(n_415),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_611),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_632),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_633),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_640),
.Y(n_697)
);

INVxp33_ASAP7_75t_L g698 ( 
.A(n_615),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_643),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_647),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_657),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_667),
.Y(n_702)
);

XNOR2xp5_ASAP7_75t_L g703 ( 
.A(n_648),
.B(n_513),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g704 ( 
.A(n_636),
.B(n_513),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_626),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_671),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_674),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_676),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_690),
.B(n_604),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_621),
.B(n_604),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_641),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_677),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_681),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_621),
.B(n_604),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_691),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_646),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_650),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_616),
.B(n_606),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_618),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_688),
.B(n_507),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_616),
.B(n_606),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_670),
.Y(n_723)
);

XOR2x2_ASAP7_75t_L g724 ( 
.A(n_645),
.B(n_514),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_634),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_624),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_619),
.A2(n_501),
.B(n_555),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_637),
.Y(n_729)
);

INVxp33_ASAP7_75t_SL g730 ( 
.A(n_660),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_661),
.B(n_524),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_691),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_637),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_SL g734 ( 
.A(n_651),
.B(n_514),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_627),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_691),
.Y(n_736)
);

XOR2xp5_ASAP7_75t_L g737 ( 
.A(n_654),
.B(n_527),
.Y(n_737)
);

XNOR2x2_ASAP7_75t_L g738 ( 
.A(n_628),
.B(n_606),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_669),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_627),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_651),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_686),
.Y(n_742)
);

XNOR2xp5_ASAP7_75t_L g743 ( 
.A(n_689),
.B(n_550),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_686),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_652),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_649),
.B(n_545),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_623),
.B(n_524),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_655),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_613),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_655),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_638),
.B(n_482),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_658),
.B(n_524),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_672),
.B(n_606),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_653),
.B(n_211),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_673),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_625),
.B(n_211),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_659),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_610),
.B(n_211),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_663),
.B(n_540),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_685),
.B(n_225),
.Y(n_760)
);

XNOR2xp5_ASAP7_75t_L g761 ( 
.A(n_614),
.B(n_550),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_630),
.B(n_483),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_675),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_659),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_620),
.B(n_468),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_678),
.Y(n_766)
);

XNOR2x2_ASAP7_75t_L g767 ( 
.A(n_619),
.B(n_606),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_678),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_692),
.A2(n_508),
.B(n_500),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_680),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_630),
.B(n_540),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_688),
.B(n_436),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_635),
.B(n_415),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_663),
.B(n_503),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_629),
.B(n_437),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_629),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_760),
.B(n_684),
.C(n_227),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_693),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_735),
.B(n_680),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_763),
.B(n_687),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_694),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_695),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_726),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_717),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_740),
.B(n_683),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_755),
.B(n_763),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_730),
.A2(n_652),
.B1(n_642),
.B2(n_639),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_767),
.A2(n_184),
.B1(n_756),
.B2(n_743),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_698),
.B(n_683),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_612),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_746),
.B(n_612),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_769),
.A2(n_519),
.B(n_508),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_697),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_748),
.B(n_750),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_714),
.B(n_687),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_757),
.B(n_617),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_771),
.B(n_617),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_764),
.B(n_639),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_714),
.B(n_624),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_722),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_723),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_719),
.B(n_639),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_705),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_726),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_699),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_745),
.B(n_552),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_726),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_728),
.B(n_624),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_754),
.B(n_758),
.C(n_776),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_719),
.B(n_639),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_741),
.B(n_556),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_709),
.B(n_631),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_762),
.B(n_631),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_700),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_701),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_702),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_746),
.A2(n_227),
.B1(n_180),
.B2(n_225),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_776),
.B(n_631),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_711),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_706),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_707),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_762),
.B(n_668),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_747),
.B(n_668),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_771),
.B(n_668),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_725),
.B(n_666),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_727),
.B(n_666),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_710),
.B(n_751),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_708),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_751),
.B(n_620),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_775),
.B(n_644),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_716),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_712),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_752),
.B(n_739),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_731),
.B(n_664),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_749),
.B(n_662),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_775),
.B(n_190),
.C(n_185),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_726),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_718),
.B(n_500),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_773),
.B(n_644),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_773),
.B(n_665),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_749),
.B(n_561),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_732),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_713),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_742),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_753),
.B(n_202),
.C(n_190),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_736),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_729),
.B(n_666),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_778),
.Y(n_849)
);

AND2x6_ASAP7_75t_L g850 ( 
.A(n_788),
.B(n_733),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_787),
.B(n_744),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_828),
.B(n_790),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_778),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_782),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_783),
.Y(n_855)
);

OAI221xp5_ASAP7_75t_L g856 ( 
.A1(n_789),
.A2(n_734),
.B1(n_761),
.B2(n_737),
.C(n_753),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_834),
.B(n_753),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_843),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_828),
.B(n_718),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_794),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_794),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_843),
.Y(n_862)
);

AO22x2_ASAP7_75t_L g863 ( 
.A1(n_814),
.A2(n_721),
.B1(n_738),
.B2(n_766),
.Y(n_863)
);

CKINVDCx16_ASAP7_75t_R g864 ( 
.A(n_824),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_814),
.A2(n_721),
.B1(n_770),
.B2(n_768),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_789),
.A2(n_741),
.B1(n_724),
.B2(n_704),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_847),
.B(n_715),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_847),
.B(n_715),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_791),
.B(n_774),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_806),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_813),
.Y(n_871)
);

OAI221xp5_ASAP7_75t_L g872 ( 
.A1(n_818),
.A2(n_703),
.B1(n_561),
.B2(n_551),
.C(n_221),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_836),
.B(n_759),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_810),
.A2(n_759),
.B1(n_774),
.B2(n_476),
.Y(n_874)
);

AO22x2_ASAP7_75t_L g875 ( 
.A1(n_823),
.A2(n_772),
.B1(n_679),
.B2(n_682),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_806),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_795),
.B(n_772),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_805),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_781),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_845),
.B(n_720),
.Y(n_880)
);

AO22x2_ASAP7_75t_L g881 ( 
.A1(n_823),
.A2(n_679),
.B1(n_682),
.B2(n_665),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_815),
.Y(n_882)
);

AO22x2_ASAP7_75t_L g883 ( 
.A1(n_796),
.A2(n_846),
.B1(n_831),
.B2(n_830),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_785),
.B(n_720),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_777),
.A2(n_476),
.B1(n_481),
.B2(n_475),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_801),
.B(n_720),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_815),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_817),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_805),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_817),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_843),
.B(n_503),
.Y(n_891)
);

OAI221xp5_ASAP7_75t_L g892 ( 
.A1(n_818),
.A2(n_551),
.B1(n_221),
.B2(n_223),
.C(n_202),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_800),
.A2(n_720),
.B1(n_279),
.B2(n_2),
.Y(n_893)
);

OAI221xp5_ASAP7_75t_L g894 ( 
.A1(n_837),
.A2(n_842),
.B1(n_809),
.B2(n_830),
.C(n_831),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_802),
.B(n_720),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_816),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_843),
.B(n_803),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_796),
.A2(n_568),
.B1(n_664),
.B2(n_507),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_797),
.B(n_666),
.Y(n_899)
);

AO22x2_ASAP7_75t_L g900 ( 
.A1(n_840),
.A2(n_841),
.B1(n_800),
.B2(n_822),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_821),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_811),
.B(n_662),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_836),
.B(n_662),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_792),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_829),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_833),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_844),
.Y(n_907)
);

CKINVDCx16_ASAP7_75t_R g908 ( 
.A(n_835),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_792),
.B(n_780),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_780),
.B(n_519),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_804),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_820),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_832),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_809),
.A2(n_476),
.B1(n_475),
.B2(n_481),
.Y(n_914)
);

AO22x2_ASAP7_75t_L g915 ( 
.A1(n_840),
.A2(n_568),
.B1(n_507),
.B2(n_2),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_779),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_799),
.B(n_521),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_786),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_825),
.Y(n_919)
);

AO22x2_ASAP7_75t_L g920 ( 
.A1(n_841),
.A2(n_568),
.B1(n_1),
.B2(n_3),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_784),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_808),
.B(n_521),
.Y(n_922)
);

AO22x2_ASAP7_75t_L g923 ( 
.A1(n_839),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_L g924 ( 
.A(n_825),
.B(n_547),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_826),
.B(n_0),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_924),
.A2(n_812),
.B(n_827),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_883),
.A2(n_848),
.B(n_807),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_852),
.B(n_798),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_L g929 ( 
.A(n_850),
.B(n_798),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_897),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_919),
.B(n_798),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_866),
.A2(n_819),
.B(n_798),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_883),
.A2(n_765),
.B(n_819),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_863),
.A2(n_765),
.B(n_793),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_864),
.B(n_798),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_849),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_853),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_856),
.A2(n_825),
.B(n_228),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_908),
.B(n_825),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_894),
.B(n_4),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_863),
.A2(n_492),
.B(n_468),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_875),
.A2(n_492),
.B(n_558),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_L g943 ( 
.A(n_892),
.B(n_228),
.C(n_223),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_875),
.A2(n_881),
.B(n_900),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_850),
.A2(n_825),
.B(n_476),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_916),
.B(n_838),
.Y(n_946)
);

AOI21xp33_ASAP7_75t_L g947 ( 
.A1(n_900),
.A2(n_838),
.B(n_205),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_881),
.A2(n_508),
.B(n_500),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_909),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_860),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_918),
.B(n_5),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_898),
.A2(n_449),
.B(n_448),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_861),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_870),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_871),
.B(n_6),
.Y(n_955)
);

BUFx8_ASAP7_75t_L g956 ( 
.A(n_850),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_859),
.B(n_6),
.Y(n_957)
);

O2A1O1Ixp5_ASAP7_75t_L g958 ( 
.A1(n_925),
.A2(n_278),
.B(n_316),
.C(n_317),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_898),
.A2(n_496),
.B(n_477),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_876),
.Y(n_960)
);

BUFx8_ASAP7_75t_L g961 ( 
.A(n_917),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_874),
.A2(n_495),
.B1(n_543),
.B2(n_521),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_882),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_872),
.A2(n_225),
.B(n_231),
.C(n_9),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_915),
.A2(n_494),
.B1(n_475),
.B2(n_481),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_904),
.B(n_7),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_873),
.B(n_8),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_885),
.A2(n_203),
.B(n_205),
.C(n_231),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_915),
.A2(n_494),
.B1(n_475),
.B2(n_481),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_851),
.B(n_9),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_911),
.B(n_10),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_912),
.B(n_10),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_887),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_888),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_L g975 ( 
.A1(n_880),
.A2(n_317),
.B(n_432),
.C(n_13),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_890),
.Y(n_976)
);

OAI321xp33_ASAP7_75t_L g977 ( 
.A1(n_914),
.A2(n_203),
.A3(n_205),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_884),
.A2(n_494),
.B(n_231),
.Y(n_978)
);

NAND2x1p5_ASAP7_75t_L g979 ( 
.A(n_878),
.B(n_521),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_923),
.A2(n_496),
.B(n_477),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_936),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_931),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_937),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_949),
.B(n_889),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_965),
.A2(n_923),
.B1(n_920),
.B2(n_893),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_944),
.B(n_862),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_950),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_939),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_928),
.B(n_865),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_927),
.B(n_865),
.Y(n_990)
);

INVxp33_ASAP7_75t_L g991 ( 
.A(n_967),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_935),
.B(n_867),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_979),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_960),
.Y(n_994)
);

INVx5_ASAP7_75t_L g995 ( 
.A(n_931),
.Y(n_995)
);

AND3x1_ASAP7_75t_SL g996 ( 
.A(n_956),
.B(n_855),
.C(n_854),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_961),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_946),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_956),
.B(n_858),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_943),
.A2(n_940),
.B1(n_932),
.B2(n_938),
.Y(n_1000)
);

BUFx8_ASAP7_75t_L g1001 ( 
.A(n_966),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_SL g1002 ( 
.A(n_947),
.B(n_899),
.C(n_895),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_974),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_970),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_979),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_953),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_954),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_930),
.B(n_868),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_971),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_964),
.A2(n_920),
.B(n_886),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_930),
.B(n_921),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_963),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_973),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_976),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_972),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_961),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_933),
.A2(n_877),
.B(n_913),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_951),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_957),
.B(n_896),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_955),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_929),
.Y(n_1021)
);

CKINVDCx8_ASAP7_75t_R g1022 ( 
.A(n_945),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_926),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_975),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_977),
.B(n_902),
.C(n_901),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_969),
.B(n_903),
.Y(n_1026)
);

OR2x4_ASAP7_75t_L g1027 ( 
.A(n_945),
.B(n_905),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_977),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_978),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_934),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_968),
.B(n_907),
.C(n_906),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_959),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_978),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_962),
.B(n_11),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_942),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_980),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_952),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_R g1038 ( 
.A(n_958),
.B(n_11),
.Y(n_1038)
);

AND2x6_ASAP7_75t_SL g1039 ( 
.A(n_941),
.B(n_869),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_948),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_931),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_947),
.A2(n_879),
.B(n_910),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_979),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_939),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_981),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_982),
.B(n_857),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_985),
.A2(n_990),
.B(n_1024),
.C(n_1010),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1029),
.B(n_922),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_1000),
.A2(n_205),
.B(n_203),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_997),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_1035),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_1051)
);

NOR2xp67_ASAP7_75t_L g1052 ( 
.A(n_995),
.B(n_12),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_1030),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_1001),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1029),
.A2(n_496),
.B(n_891),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1018),
.B(n_891),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_SL g1057 ( 
.A(n_1023),
.B(n_891),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1033),
.A2(n_17),
.B(n_19),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_SL g1059 ( 
.A(n_1017),
.B(n_20),
.C(n_21),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_982),
.B(n_20),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_999),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1033),
.A2(n_1028),
.B(n_989),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1050),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_1047),
.A2(n_1036),
.B(n_986),
.C(n_1015),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1050),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1046),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1052),
.B(n_995),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1045),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1049),
.A2(n_1028),
.B1(n_1021),
.B2(n_1037),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_1059),
.A2(n_1028),
.B(n_991),
.C(n_1025),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_1054),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1056),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_1061),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1059),
.A2(n_1021),
.B(n_1031),
.C(n_984),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_1062),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1060),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1057),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1051),
.A2(n_1020),
.B(n_1032),
.C(n_1040),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1048),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1058),
.B(n_1022),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_1048),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1053),
.B(n_1009),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_1055),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1053),
.A2(n_1027),
.B1(n_995),
.B2(n_1041),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1061),
.B(n_1016),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1047),
.A2(n_1041),
.B1(n_1044),
.B2(n_988),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1050),
.B(n_998),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1084),
.A2(n_1012),
.B(n_1040),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_SL g1089 ( 
.A1(n_1074),
.A2(n_1070),
.B(n_1064),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1080),
.A2(n_1019),
.B(n_1026),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1074),
.A2(n_1002),
.B(n_1039),
.C(n_1009),
.Y(n_1091)
);

AND2x6_ASAP7_75t_L g1092 ( 
.A(n_1071),
.B(n_1009),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1086),
.A2(n_1043),
.B1(n_1008),
.B2(n_993),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1071),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1088),
.A2(n_1065),
.B(n_1063),
.Y(n_1095)
);

AO21x2_ASAP7_75t_L g1096 ( 
.A1(n_1089),
.A2(n_1080),
.B(n_1082),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1095),
.A2(n_1073),
.B(n_1093),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_1095),
.B(n_1071),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1098),
.A2(n_1085),
.A3(n_1091),
.B(n_1096),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_1071),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_1073),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1100),
.B(n_1096),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_1102),
.B(n_1081),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1102),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1101),
.Y(n_1105)
);

NAND2xp33_ASAP7_75t_R g1106 ( 
.A(n_1103),
.B(n_1094),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_1104),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_1104),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_R g1109 ( 
.A(n_1108),
.B(n_1067),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_1106),
.B(n_1105),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1109),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1110),
.B(n_1085),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_L g1113 ( 
.A(n_1112),
.B(n_1107),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1111),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_1113),
.B(n_1096),
.C(n_1070),
.Y(n_1115)
);

NAND4xp25_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_1090),
.C(n_1069),
.D(n_1078),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1115),
.B(n_1092),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_1116),
.B(n_1098),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1117),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1118),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1120),
.B(n_1092),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_1072),
.C(n_1081),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1120),
.B(n_1092),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1121),
.B(n_1087),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1122),
.B(n_1075),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1124),
.B(n_1087),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1126),
.B(n_1001),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1127),
.B(n_1125),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1128),
.B(n_1076),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1129),
.B(n_1066),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1130),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1132),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1133),
.B(n_1079),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1134),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_1136),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1135),
.A2(n_1068),
.B1(n_1083),
.B2(n_1077),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1137),
.B(n_21),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_L g1141 ( 
.A(n_1137),
.B(n_1067),
.Y(n_1141)
);

OAI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1141),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_1142)
);

NAND2x1_ASAP7_75t_L g1143 ( 
.A(n_1140),
.B(n_502),
.Y(n_1143)
);

NAND4xp25_ASAP7_75t_L g1144 ( 
.A(n_1139),
.B(n_23),
.C(n_25),
.D(n_26),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1142),
.B(n_26),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1144),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1145),
.A2(n_1143),
.B1(n_1004),
.B2(n_30),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1146),
.Y(n_1148)
);

INVxp33_ASAP7_75t_L g1149 ( 
.A(n_1148),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1147),
.B(n_27),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_R g1151 ( 
.A(n_1150),
.B(n_27),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1149),
.B(n_29),
.Y(n_1152)
);

NAND4xp75_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_29),
.C(n_30),
.D(n_31),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1152),
.B(n_1004),
.Y(n_1154)
);

AOI211xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1153),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_SL g1156 ( 
.A1(n_1154),
.A2(n_32),
.B(n_34),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1155),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1156),
.B(n_35),
.C(n_36),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1156),
.B(n_35),
.Y(n_1159)
);

NAND4xp25_ASAP7_75t_SL g1160 ( 
.A(n_1158),
.B(n_36),
.C(n_37),
.D(n_38),
.Y(n_1160)
);

AOI211xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1157),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1159),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1162),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1160),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1164),
.A2(n_1161),
.B(n_39),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1163),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1166),
.B(n_40),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1165),
.A2(n_494),
.B1(n_502),
.B2(n_43),
.Y(n_1168)
);

NOR2x1_ASAP7_75t_L g1169 ( 
.A(n_1167),
.B(n_502),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1168),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1170),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.C(n_46),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1169),
.B(n_49),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1172),
.B(n_54),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1171),
.B(n_390),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1174),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1173),
.Y(n_1176)
);

XNOR2x1_ASAP7_75t_L g1177 ( 
.A(n_1174),
.B(n_55),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1176),
.A2(n_1034),
.B(n_1038),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1175),
.A2(n_56),
.B(n_57),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1177),
.A2(n_59),
.B(n_60),
.Y(n_1180)
);

NAND4xp25_ASAP7_75t_L g1181 ( 
.A(n_1180),
.B(n_61),
.C(n_63),
.D(n_65),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1179),
.B(n_67),
.Y(n_1182)
);

AOI31xp33_ASAP7_75t_L g1183 ( 
.A1(n_1182),
.A2(n_1178),
.A3(n_69),
.B(n_71),
.Y(n_1183)
);

OA211x2_ASAP7_75t_L g1184 ( 
.A1(n_1181),
.A2(n_68),
.B(n_72),
.C(n_74),
.Y(n_1184)
);

OR3x2_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_76),
.C(n_77),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1183),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1186),
.B(n_79),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1185),
.A2(n_494),
.B1(n_83),
.B2(n_84),
.Y(n_1188)
);

OAI211xp5_ASAP7_75t_L g1189 ( 
.A1(n_1188),
.A2(n_80),
.B(n_85),
.C(n_88),
.Y(n_1189)
);

XNOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1187),
.B(n_89),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_1190),
.Y(n_1191)
);

XOR2x2_ASAP7_75t_L g1192 ( 
.A(n_1189),
.B(n_90),
.Y(n_1192)
);

XOR2xp5_ASAP7_75t_L g1193 ( 
.A(n_1191),
.B(n_91),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_R g1194 ( 
.A1(n_1192),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1191),
.Y(n_1195)
);

BUFx4f_ASAP7_75t_SL g1196 ( 
.A(n_1195),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1194),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_1193),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1196),
.Y(n_1199)
);

INVxp67_ASAP7_75t_SL g1200 ( 
.A(n_1197),
.Y(n_1200)
);

XNOR2xp5_ASAP7_75t_L g1201 ( 
.A(n_1199),
.B(n_1198),
.Y(n_1201)
);

XNOR2xp5_ASAP7_75t_L g1202 ( 
.A(n_1200),
.B(n_96),
.Y(n_1202)
);

AOI221xp5_ASAP7_75t_L g1203 ( 
.A1(n_1201),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.C(n_100),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1202),
.A2(n_101),
.B(n_102),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1201),
.B(n_103),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1204),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1205),
.A2(n_1005),
.B1(n_993),
.B2(n_1043),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1203),
.A2(n_1005),
.B1(n_993),
.B2(n_566),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1206),
.A2(n_1208),
.B1(n_1207),
.B2(n_113),
.C(n_114),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1206),
.A2(n_111),
.B(n_112),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1206),
.B(n_116),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1211),
.A2(n_117),
.B(n_118),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1209),
.A2(n_1210),
.B(n_120),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1211),
.B(n_1005),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1211),
.B(n_119),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1211),
.A2(n_121),
.B(n_123),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1211),
.A2(n_124),
.B(n_125),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1211),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1210),
.B(n_126),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1211),
.B(n_127),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1211),
.A2(n_128),
.B(n_129),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1211),
.B(n_130),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1211),
.A2(n_131),
.B(n_133),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1211),
.B(n_134),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1218),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_1225)
);

AOI322xp5_ASAP7_75t_L g1226 ( 
.A1(n_1213),
.A2(n_139),
.A3(n_140),
.B1(n_141),
.B2(n_142),
.C1(n_143),
.C2(n_144),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1219),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_1227)
);

OAI221xp5_ASAP7_75t_R g1228 ( 
.A1(n_1224),
.A2(n_150),
.B1(n_153),
.B2(n_155),
.C(n_156),
.Y(n_1228)
);

OAI221xp5_ASAP7_75t_R g1229 ( 
.A1(n_1215),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.C(n_166),
.Y(n_1229)
);

AOI322xp5_ASAP7_75t_L g1230 ( 
.A1(n_1220),
.A2(n_167),
.A3(n_168),
.B1(n_169),
.B2(n_171),
.C1(n_172),
.C2(n_173),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1222),
.A2(n_178),
.B1(n_543),
.B2(n_566),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1212),
.A2(n_566),
.B1(n_543),
.B2(n_390),
.Y(n_1232)
);

AOI222xp33_ASAP7_75t_L g1233 ( 
.A1(n_1214),
.A2(n_390),
.B1(n_566),
.B2(n_543),
.C1(n_415),
.C2(n_457),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1232),
.A2(n_1223),
.B1(n_1221),
.B2(n_1216),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1231),
.A2(n_1217),
.B1(n_467),
.B2(n_480),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1229),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1228),
.A2(n_1008),
.B(n_1011),
.Y(n_1237)
);

OAI321xp33_ASAP7_75t_L g1238 ( 
.A1(n_1227),
.A2(n_996),
.A3(n_457),
.B1(n_491),
.B2(n_486),
.C(n_480),
.Y(n_1238)
);

AO221x2_ASAP7_75t_L g1239 ( 
.A1(n_1226),
.A2(n_1014),
.B1(n_1007),
.B2(n_1013),
.C(n_983),
.Y(n_1239)
);

AOI221xp5_ASAP7_75t_L g1240 ( 
.A1(n_1236),
.A2(n_1233),
.B1(n_1230),
.B2(n_1225),
.C(n_491),
.Y(n_1240)
);

AOI221x1_ASAP7_75t_L g1241 ( 
.A1(n_1234),
.A2(n_1235),
.B1(n_1237),
.B2(n_1239),
.C(n_1238),
.Y(n_1241)
);

AOI221xp5_ASAP7_75t_L g1242 ( 
.A1(n_1236),
.A2(n_479),
.B1(n_467),
.B2(n_486),
.C(n_491),
.Y(n_1242)
);

AOI221xp5_ASAP7_75t_L g1243 ( 
.A1(n_1236),
.A2(n_479),
.B1(n_467),
.B2(n_486),
.C(n_491),
.Y(n_1243)
);

AOI221xp5_ASAP7_75t_L g1244 ( 
.A1(n_1240),
.A2(n_1011),
.B1(n_1012),
.B2(n_1006),
.C(n_981),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1244),
.A2(n_1241),
.B1(n_1242),
.B2(n_1243),
.Y(n_1245)
);

AOI211xp5_ASAP7_75t_L g1246 ( 
.A1(n_1245),
.A2(n_992),
.B(n_983),
.C(n_994),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1246),
.A2(n_1042),
.B1(n_1003),
.B2(n_987),
.Y(n_1247)
);


endmodule