module fake_jpeg_5272_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_60),
.C(n_44),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_32),
.B1(n_16),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_23),
.B1(n_20),
.B2(n_16),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_64),
.B1(n_47),
.B2(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_62),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_18),
.B1(n_34),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_34),
.B1(n_17),
.B2(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_41),
.B1(n_39),
.B2(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_67),
.B1(n_35),
.B2(n_45),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_35),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_81),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_46),
.B1(n_43),
.B2(n_38),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_80),
.B(n_43),
.C(n_70),
.Y(n_133)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_83),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_91),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_46),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_100),
.B1(n_72),
.B2(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_43),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_90),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_60),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_55),
.B1(n_54),
.B2(n_67),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_71),
.B1(n_49),
.B2(n_62),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_17),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_98),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_50),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_108),
.C(n_88),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_112),
.B1(n_115),
.B2(n_92),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_113),
.A2(n_52),
.B(n_29),
.C(n_43),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_69),
.B1(n_61),
.B2(n_65),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_63),
.B1(n_43),
.B2(n_70),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_79),
.B1(n_78),
.B2(n_68),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_69),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_109),
.B(n_116),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_130),
.B(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_74),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_72),
.B(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_141),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_155),
.B(n_159),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_137),
.A2(n_156),
.B1(n_161),
.B2(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_160),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_76),
.B(n_91),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_97),
.A3(n_17),
.B1(n_22),
.B2(n_119),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_152),
.Y(n_194)
);

OR2x6_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_104),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_122),
.B(n_114),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_81),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_77),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_145),
.B(n_153),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_107),
.A2(n_101),
.B1(n_98),
.B2(n_84),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_113),
.B1(n_121),
.B2(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_52),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_125),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_74),
.B1(n_102),
.B2(n_90),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_117),
.A2(n_40),
.B1(n_68),
.B2(n_103),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_168),
.B1(n_147),
.B2(n_148),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_121),
.B1(n_111),
.B2(n_114),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_122),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_171),
.A2(n_173),
.B(n_174),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_111),
.C(n_129),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_176),
.C(n_200),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_97),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_179),
.B1(n_136),
.B2(n_162),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_105),
.B(n_43),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_188),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_123),
.B(n_129),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_125),
.B1(n_105),
.B2(n_123),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_186),
.B1(n_190),
.B2(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_34),
.B1(n_97),
.B2(n_27),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_17),
.B(n_22),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_141),
.B1(n_161),
.B2(n_140),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_0),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_119),
.B1(n_17),
.B2(n_124),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_158),
.B1(n_162),
.B2(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_139),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_22),
.C(n_1),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_224),
.B1(n_171),
.B2(n_173),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_134),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_212),
.CI(n_214),
.CON(n_250),
.SN(n_250)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_208),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_162),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_216),
.C(n_227),
.Y(n_232)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_138),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_150),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_162),
.C(n_155),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_225),
.B1(n_183),
.B2(n_185),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_22),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_180),
.B(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_167),
.A2(n_139),
.B1(n_144),
.B2(n_22),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_186),
.B1(n_182),
.B2(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_15),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_169),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_0),
.C(n_1),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_200),
.C(n_188),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_193),
.B1(n_178),
.B2(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_181),
.B(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_237),
.B1(n_224),
.B2(n_208),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_209),
.C(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_243),
.C(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_194),
.B1(n_196),
.B2(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_217),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_216),
.C(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_191),
.C(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_194),
.B1(n_185),
.B2(n_4),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_15),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_0),
.C(n_3),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_205),
.B(n_14),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_207),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_256),
.B(n_269),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_228),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_218),
.B1(n_229),
.B2(n_202),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_273),
.B1(n_231),
.B2(n_253),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_212),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_265),
.A2(n_255),
.B1(n_250),
.B2(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_221),
.B1(n_225),
.B2(n_5),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_276),
.B1(n_254),
.B2(n_235),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_3),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_248),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_4),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_245),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_236),
.B1(n_230),
.B2(n_241),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_281),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_234),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_291),
.C(n_271),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_239),
.B1(n_233),
.B2(n_249),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_232),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_238),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_297),
.B(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_268),
.C(n_266),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_268),
.C(n_258),
.Y(n_299)
);

OAI221xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_250),
.B1(n_274),
.B2(n_272),
.C(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_267),
.C(n_250),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_5),
.C(n_6),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_277),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_7),
.C(n_8),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_287),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_292),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_314),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_280),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_287),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_304),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_9),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_9),
.C(n_11),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_301),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_299),
.B1(n_297),
.B2(n_301),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_325),
.B(n_327),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_328),
.B(n_319),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_320),
.B(n_324),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_315),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_334),
.B(n_322),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_310),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_321),
.B(n_323),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_333),
.B1(n_329),
.B2(n_331),
.Y(n_339)
);

AOI221xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_11),
.B1(n_12),
.B2(n_337),
.C(n_334),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_11),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_11),
.Y(n_342)
);


endmodule