module real_aes_7049_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_241;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g489 ( .A(n_1), .Y(n_489) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_3), .A2(n_37), .B1(n_175), .B2(n_498), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g214 ( .A1(n_4), .A2(n_132), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_5), .B(n_162), .Y(n_481) );
AND2x6_ASAP7_75t_L g137 ( .A(n_6), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_7), .A2(n_183), .B(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_38), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_9), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g220 ( .A(n_10), .Y(n_220) );
INVx1_ASAP7_75t_L g158 ( .A(n_11), .Y(n_158) );
INVx1_ASAP7_75t_L g485 ( .A(n_12), .Y(n_485) );
INVx1_ASAP7_75t_L g191 ( .A(n_13), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_14), .B(n_206), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_15), .B(n_154), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_16), .A2(n_41), .B1(n_727), .B2(n_728), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_16), .Y(n_728) );
AO32x2_ASAP7_75t_L g495 ( .A1(n_17), .A2(n_153), .A3(n_162), .B1(n_467), .B2(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_18), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_19), .B(n_175), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_20), .B(n_148), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_21), .B(n_154), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_22), .A2(n_49), .B1(n_175), .B2(n_498), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_23), .B(n_132), .Y(n_131) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_24), .A2(n_76), .B1(n_175), .B2(n_206), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_25), .B(n_175), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_26), .B(n_213), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_27), .A2(n_188), .B(n_190), .C(n_192), .Y(n_187) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_29), .B(n_166), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_30), .B(n_173), .Y(n_204) );
INVx1_ASAP7_75t_L g230 ( .A(n_31), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_32), .B(n_166), .Y(n_511) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_34), .B(n_175), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_35), .B(n_166), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_36), .A2(n_137), .B(n_140), .C(n_143), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_38), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g228 ( .A(n_39), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_40), .B(n_173), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_41), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_42), .B(n_175), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_43), .A2(n_86), .B1(n_151), .B2(n_498), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_44), .B(n_175), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_45), .B(n_175), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_46), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_47), .B(n_465), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_48), .B(n_132), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_50), .A2(n_59), .B1(n_175), .B2(n_206), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_51), .A2(n_140), .B1(n_206), .B2(n_227), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_52), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_53), .B(n_175), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_54), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_55), .B(n_175), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_56), .A2(n_218), .B(n_219), .C(n_221), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_57), .Y(n_268) );
INVx1_ASAP7_75t_L g216 ( .A(n_58), .Y(n_216) );
INVx1_ASAP7_75t_L g138 ( .A(n_60), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_61), .B(n_175), .Y(n_490) );
INVx1_ASAP7_75t_L g157 ( .A(n_62), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_63), .Y(n_742) );
AO32x2_ASAP7_75t_L g531 ( .A1(n_64), .A2(n_162), .A3(n_165), .B1(n_467), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g463 ( .A(n_65), .Y(n_463) );
INVx1_ASAP7_75t_L g506 ( .A(n_66), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_67), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_SL g238 ( .A1(n_68), .A2(n_148), .B(n_221), .C(n_239), .Y(n_238) );
INVxp67_ASAP7_75t_L g240 ( .A(n_69), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_70), .B(n_206), .Y(n_507) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_72), .A2(n_102), .B1(n_114), .B2(n_758), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_73), .Y(n_233) );
INVx1_ASAP7_75t_L g261 ( .A(n_74), .Y(n_261) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_75), .A2(n_88), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_75), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_77), .A2(n_137), .B(n_140), .C(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_78), .B(n_498), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_79), .B(n_206), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_80), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g155 ( .A(n_81), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_82), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_83), .B(n_206), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_84), .A2(n_137), .B(n_140), .C(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g110 ( .A(n_85), .Y(n_110) );
OR2x2_ASAP7_75t_L g120 ( .A(n_85), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g751 ( .A(n_85), .B(n_738), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_87), .A2(n_100), .B1(n_206), .B2(n_207), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_88), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_89), .B(n_166), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_90), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_91), .A2(n_137), .B(n_140), .C(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_92), .Y(n_178) );
INVx1_ASAP7_75t_L g237 ( .A(n_93), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_94), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_95), .B(n_145), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_96), .B(n_206), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_97), .B(n_162), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_98), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_99), .A2(n_132), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g758 ( .A(n_104), .Y(n_758) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g450 ( .A(n_110), .B(n_121), .Y(n_450) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_110), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO221x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_740), .B1(n_743), .B2(n_752), .C(n_754), .Y(n_114) );
OAI222xp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_726), .B1(n_729), .B2(n_733), .C1(n_734), .C2(n_739), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B1(n_448), .B2(n_451), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_120), .A2(n_448), .B1(n_731), .B2(n_732), .Y(n_730) );
INVx2_ASAP7_75t_L g738 ( .A(n_121), .Y(n_738) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx2_ASAP7_75t_L g731 ( .A(n_124), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_124), .A2(n_731), .B1(n_746), .B2(n_747), .Y(n_745) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_417), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_310), .C(n_383), .Y(n_125) );
OAI211xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_195), .B(n_242), .C(n_294), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
AND2x2_ASAP7_75t_L g258 ( .A(n_129), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g277 ( .A(n_129), .Y(n_277) );
INVx2_ASAP7_75t_L g292 ( .A(n_129), .Y(n_292) );
INVx1_ASAP7_75t_L g322 ( .A(n_129), .Y(n_322) );
AND2x2_ASAP7_75t_L g372 ( .A(n_129), .B(n_293), .Y(n_372) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_129), .A2(n_327), .A3(n_400), .B1(n_402), .B2(n_403), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_129), .B(n_248), .Y(n_405) );
AND2x2_ASAP7_75t_L g432 ( .A(n_129), .B(n_275), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_129), .B(n_441), .Y(n_440) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_159), .Y(n_129) );
AOI21xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_139), .B(n_152), .Y(n_130) );
BUFx2_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_133), .B(n_137), .Y(n_200) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g465 ( .A(n_134), .Y(n_465) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g207 ( .A(n_135), .Y(n_207) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx3_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
INVx4_ASAP7_75t_SL g193 ( .A(n_137), .Y(n_193) );
BUFx3_ASAP7_75t_L g467 ( .A(n_137), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_137), .A2(n_474), .B(n_477), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_137), .A2(n_484), .B(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_137), .A2(n_505), .B(n_508), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_137), .A2(n_514), .B(n_518), .Y(n_513) );
INVx5_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx3_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx1_ASAP7_75t_L g498 ( .A(n_141), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B(n_149), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_145), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_145), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_145), .A2(n_475), .B(n_476), .Y(n_474) );
INVx2_ASAP7_75t_L g480 ( .A(n_145), .Y(n_480) );
O2A1O1Ixp5_ASAP7_75t_SL g505 ( .A1(n_145), .A2(n_221), .B(n_506), .C(n_507), .Y(n_505) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_146), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_146), .B(n_240), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g532 ( .A1(n_146), .A2(n_173), .B1(n_533), .B2(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g517 ( .A(n_148), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_149), .A2(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
INVx1_ASAP7_75t_L g266 ( .A(n_152), .Y(n_266) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_152), .A2(n_458), .B(n_468), .Y(n_457) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_152), .A2(n_483), .B(n_491), .Y(n_482) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_153), .A2(n_198), .B(n_208), .Y(n_197) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_153), .A2(n_225), .B(n_232), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_153), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_155), .B(n_156), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
AO21x1_ASAP7_75t_L g543 ( .A1(n_161), .A2(n_544), .B(n_547), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_161), .B(n_467), .C(n_544), .Y(n_568) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_162), .A2(n_235), .B(n_241), .Y(n_234) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_162), .A2(n_473), .B(n_481), .Y(n_472) );
AND2x2_ASAP7_75t_L g321 ( .A(n_163), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g343 ( .A(n_163), .Y(n_343) );
AND2x2_ASAP7_75t_L g428 ( .A(n_163), .B(n_258), .Y(n_428) );
AND2x2_ASAP7_75t_L g431 ( .A(n_163), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
INVx2_ASAP7_75t_L g250 ( .A(n_164), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_164), .B(n_275), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_164), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g327 ( .A(n_164), .Y(n_327) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_177), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g179 ( .A(n_166), .Y(n_179) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_166), .A2(n_182), .B(n_194), .Y(n_181) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_166), .A2(n_504), .B(n_511), .Y(n_503) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_166), .A2(n_513), .B(n_521), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_176), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_174), .Y(n_169) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_173), .A2(n_480), .B1(n_497), .B2(n_499), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_173), .A2(n_480), .B1(n_545), .B2(n_546), .Y(n_544) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_179), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_179), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_180), .B(n_250), .Y(n_269) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
AND2x2_ASAP7_75t_L g293 ( .A(n_181), .B(n_275), .Y(n_293) );
AND2x2_ASAP7_75t_L g362 ( .A(n_181), .B(n_259), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_193), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_186), .A2(n_193), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_186), .A2(n_193), .B(n_237), .C(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_188), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g487 ( .A(n_188), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_188), .A2(n_509), .B(n_510), .Y(n_508) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g227 ( .A1(n_189), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_227) );
INVx2_ASAP7_75t_L g229 ( .A(n_189), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_193), .A2(n_200), .B1(n_226), .B2(n_231), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
OR2x2_ASAP7_75t_L g256 ( .A(n_196), .B(n_224), .Y(n_256) );
INVx1_ASAP7_75t_L g335 ( .A(n_196), .Y(n_335) );
AND2x2_ASAP7_75t_L g349 ( .A(n_196), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_196), .B(n_223), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_196), .B(n_347), .Y(n_401) );
AND2x2_ASAP7_75t_L g409 ( .A(n_196), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
AND2x2_ASAP7_75t_L g316 ( .A(n_197), .B(n_224), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_200), .A2(n_261), .B(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_205), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_210), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_210), .Y(n_443) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_223), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_211), .B(n_287), .Y(n_309) );
OR2x2_ASAP7_75t_L g338 ( .A(n_211), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g370 ( .A(n_211), .B(n_350), .Y(n_370) );
INVx1_ASAP7_75t_SL g390 ( .A(n_211), .Y(n_390) );
AND2x2_ASAP7_75t_L g394 ( .A(n_211), .B(n_255), .Y(n_394) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_212), .B(n_223), .Y(n_247) );
AND2x2_ASAP7_75t_L g254 ( .A(n_212), .B(n_234), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_212), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g297 ( .A(n_212), .B(n_279), .Y(n_297) );
INVx1_ASAP7_75t_SL g304 ( .A(n_212), .Y(n_304) );
BUFx2_ASAP7_75t_L g315 ( .A(n_212), .Y(n_315) );
AND2x2_ASAP7_75t_L g331 ( .A(n_212), .B(n_246), .Y(n_331) );
AND2x2_ASAP7_75t_L g346 ( .A(n_212), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g410 ( .A(n_212), .B(n_224), .Y(n_410) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_222), .Y(n_212) );
O2A1O1Ixp5_ASAP7_75t_L g462 ( .A1(n_218), .A2(n_463), .B(n_464), .C(n_466), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_218), .A2(n_519), .B(n_520), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_223), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g334 ( .A(n_223), .B(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_223), .A2(n_352), .B1(n_355), .B2(n_358), .C(n_363), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_223), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_234), .Y(n_223) );
INVx3_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
BUFx2_ASAP7_75t_L g289 ( .A(n_234), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_234), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
OR2x2_ASAP7_75t_L g339 ( .A(n_234), .B(n_279), .Y(n_339) );
INVx3_ASAP7_75t_L g347 ( .A(n_234), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_234), .B(n_279), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B1(n_252), .B2(n_257), .C(n_270), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_245), .B(n_319), .Y(n_444) );
OR2x2_ASAP7_75t_L g447 ( .A(n_245), .B(n_278), .Y(n_447) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OAI221xp5_ASAP7_75t_SL g270 ( .A1(n_246), .A2(n_271), .B1(n_278), .B2(n_280), .C(n_283), .Y(n_270) );
AND2x2_ASAP7_75t_L g287 ( .A(n_246), .B(n_279), .Y(n_287) );
AND2x2_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_246), .B(n_303), .Y(n_302) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_246), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g397 ( .A(n_246), .B(n_339), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_248), .A2(n_357), .B1(n_386), .B2(n_388), .Y(n_385) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI322xp5_ASAP7_75t_L g294 ( .A1(n_249), .A2(n_258), .A3(n_295), .B1(n_298), .B2(n_301), .C1(n_305), .C2(n_308), .Y(n_294) );
OR2x2_ASAP7_75t_L g306 ( .A(n_249), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g285 ( .A(n_250), .B(n_259), .Y(n_285) );
INVx1_ASAP7_75t_L g300 ( .A(n_250), .Y(n_300) );
AND2x2_ASAP7_75t_L g366 ( .A(n_250), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g276 ( .A(n_251), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g367 ( .A(n_251), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_251), .B(n_275), .Y(n_441) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_255), .B(n_390), .Y(n_389) );
INVx3_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g341 ( .A(n_256), .B(n_288), .Y(n_341) );
OR2x2_ASAP7_75t_L g438 ( .A(n_256), .B(n_289), .Y(n_438) );
INVx1_ASAP7_75t_L g419 ( .A(n_257), .Y(n_419) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_269), .Y(n_257) );
INVx4_ASAP7_75t_L g307 ( .A(n_258), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_258), .B(n_326), .Y(n_332) );
INVx2_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_266), .B(n_267), .Y(n_259) );
INVx1_ASAP7_75t_L g357 ( .A(n_269), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_269), .B(n_329), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_271), .A2(n_345), .B(n_348), .Y(n_344) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx1_ASAP7_75t_L g356 ( .A(n_275), .Y(n_356) );
INVx1_ASAP7_75t_L g282 ( .A(n_276), .Y(n_282) );
AND2x2_ASAP7_75t_L g284 ( .A(n_276), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g380 ( .A(n_277), .B(n_366), .Y(n_380) );
AND2x2_ASAP7_75t_L g402 ( .A(n_277), .B(n_362), .Y(n_402) );
BUFx2_ASAP7_75t_L g354 ( .A(n_279), .Y(n_354) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AOI32xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .A3(n_287), .B1(n_288), .B2(n_290), .Y(n_283) );
INVx1_ASAP7_75t_L g364 ( .A(n_284), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_284), .A2(n_412), .B1(n_413), .B2(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_287), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_287), .B(n_346), .Y(n_387) );
AND2x2_ASAP7_75t_L g434 ( .A(n_287), .B(n_319), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_288), .B(n_335), .Y(n_382) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g435 ( .A(n_290), .Y(n_435) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_293), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g407 ( .A(n_293), .B(n_327), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_293), .B(n_322), .Y(n_414) );
INVx1_ASAP7_75t_SL g396 ( .A(n_295), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_296), .B(n_347), .Y(n_374) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_296), .B(n_319), .C(n_421), .D(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_297), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_L g377 ( .A(n_300), .Y(n_377) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_303), .A2(n_394), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g319 ( .A(n_304), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g368 ( .A(n_307), .Y(n_368) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND4xp25_ASAP7_75t_SL g310 ( .A(n_311), .B(n_336), .C(n_351), .D(n_371), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_317), .B(n_321), .C(n_323), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g403 ( .A(n_316), .B(n_346), .Y(n_403) );
AND2x2_ASAP7_75t_L g412 ( .A(n_316), .B(n_390), .Y(n_412) );
INVx3_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_319), .B(n_354), .Y(n_416) );
AND2x2_ASAP7_75t_L g328 ( .A(n_322), .B(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_330), .B1(n_332), .B2(n_333), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g426 ( .A(n_326), .B(n_372), .Y(n_426) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_328), .B(n_377), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_329), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B(n_342), .C(n_344), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_372), .B1(n_373), .B2(n_375), .C(n_378), .Y(n_371) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_345), .A2(n_430), .B1(n_433), .B2(n_435), .C(n_436), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_346), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_354), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_359), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_369), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_368), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_379), .A2(n_405), .B1(n_443), .B2(n_444), .C(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_391), .C(n_411), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_395), .C(n_404), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_398), .C(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g423 ( .A(n_401), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_402), .A2(n_428), .B(n_446), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_414), .A2(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_429), .C(n_442), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_425), .C(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx14_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g732 ( .A(n_451), .Y(n_732) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR3x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_654), .C(n_703), .Y(n_452) );
NAND5xp2_ASAP7_75t_L g453 ( .A(n_454), .B(n_569), .C(n_597), .D(n_627), .E(n_641), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_492), .B1(n_522), .B2(n_527), .C(n_536), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_469), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_456), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
AND2x2_ASAP7_75t_L g557 ( .A(n_457), .B(n_472), .Y(n_557) );
AND2x2_ASAP7_75t_L g580 ( .A(n_457), .B(n_471), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_457), .B(n_482), .Y(n_595) );
OR2x2_ASAP7_75t_L g604 ( .A(n_457), .B(n_543), .Y(n_604) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_457), .Y(n_607) );
AND2x2_ASAP7_75t_L g715 ( .A(n_457), .B(n_543), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_467), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_464), .A2(n_480), .B(n_489), .C(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_469), .B(n_607), .Y(n_663) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OAI311xp33_ASAP7_75t_L g605 ( .A1(n_470), .A2(n_606), .A3(n_607), .B1(n_608), .C1(n_623), .Y(n_605) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_482), .Y(n_470) );
AND2x2_ASAP7_75t_L g566 ( .A(n_471), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g573 ( .A(n_471), .Y(n_573) );
AND2x2_ASAP7_75t_L g694 ( .A(n_471), .B(n_526), .Y(n_694) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_472), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g550 ( .A(n_472), .B(n_482), .Y(n_550) );
AND2x2_ASAP7_75t_L g602 ( .A(n_472), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g616 ( .A(n_472), .B(n_549), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_480), .Y(n_477) );
INVx2_ASAP7_75t_L g526 ( .A(n_482), .Y(n_526) );
AND2x2_ASAP7_75t_L g565 ( .A(n_482), .B(n_549), .Y(n_565) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_500), .Y(n_492) );
OR2x2_ASAP7_75t_L g660 ( .A(n_493), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_493), .B(n_666), .Y(n_677) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_494), .B(n_673), .Y(n_672) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g535 ( .A(n_495), .Y(n_535) );
AND2x2_ASAP7_75t_L g601 ( .A(n_495), .B(n_531), .Y(n_601) );
AND2x2_ASAP7_75t_L g612 ( .A(n_495), .B(n_512), .Y(n_612) );
AND2x2_ASAP7_75t_L g621 ( .A(n_495), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_500), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_500), .B(n_562), .Y(n_606) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g593 ( .A(n_501), .B(n_552), .Y(n_593) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
INVx2_ASAP7_75t_L g529 ( .A(n_502), .Y(n_529) );
AND2x2_ASAP7_75t_L g620 ( .A(n_502), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g539 ( .A(n_503), .Y(n_539) );
OR2x2_ASAP7_75t_L g637 ( .A(n_503), .B(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_503), .Y(n_700) );
AND2x2_ASAP7_75t_L g540 ( .A(n_512), .B(n_535), .Y(n_540) );
INVx1_ASAP7_75t_L g560 ( .A(n_512), .Y(n_560) );
AND2x2_ASAP7_75t_L g581 ( .A(n_512), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g622 ( .A(n_512), .Y(n_622) );
INVx1_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_512), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVxp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_524), .B(n_626), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_524), .A2(n_611), .B1(n_660), .B2(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_525), .A2(n_704), .B(n_706), .C(n_724), .Y(n_703) );
INVx2_ASAP7_75t_L g556 ( .A(n_526), .Y(n_556) );
AND2x2_ASAP7_75t_L g614 ( .A(n_526), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g625 ( .A(n_526), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_527), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
AND2x2_ASAP7_75t_L g598 ( .A(n_528), .B(n_562), .Y(n_598) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g630 ( .A(n_529), .B(n_621), .Y(n_630) );
AND2x2_ASAP7_75t_L g649 ( .A(n_529), .B(n_563), .Y(n_649) );
AND2x4_ASAP7_75t_L g585 ( .A(n_530), .B(n_559), .Y(n_585) );
AND2x2_ASAP7_75t_L g723 ( .A(n_530), .B(n_699), .Y(n_723) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
INVx1_ASAP7_75t_L g563 ( .A(n_531), .Y(n_563) );
INVx1_ASAP7_75t_L g662 ( .A(n_531), .Y(n_662) );
OR2x2_ASAP7_75t_L g553 ( .A(n_535), .B(n_539), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_535), .B(n_563), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g582 ( .A(n_535), .B(n_583), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_541), .B1(n_551), .B2(n_554), .C(n_558), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_538), .A2(n_559), .B(n_561), .C(n_564), .Y(n_558) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g583 ( .A(n_539), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_539), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_539), .B(n_560), .Y(n_666) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_539), .Y(n_673) );
AND2x2_ASAP7_75t_L g591 ( .A(n_540), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g628 ( .A(n_540), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_550), .Y(n_541) );
INVx2_ASAP7_75t_L g619 ( .A(n_542), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_542), .A2(n_552), .B1(n_669), .B2(n_671), .C1(n_672), .C2(n_674), .Y(n_668) );
AND2x2_ASAP7_75t_L g725 ( .A(n_542), .B(n_694), .Y(n_725) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_549), .Y(n_542) );
INVx1_ASAP7_75t_L g615 ( .A(n_543), .Y(n_615) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g567 ( .A(n_548), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g653 ( .A(n_550), .B(n_587), .Y(n_653) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_551), .A2(n_665), .B(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g592 ( .A(n_552), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_552), .B(n_559), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_552), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx3_ASAP7_75t_L g618 ( .A(n_556), .Y(n_618) );
OR2x2_ASAP7_75t_L g670 ( .A(n_556), .B(n_592), .Y(n_670) );
AND2x2_ASAP7_75t_L g586 ( .A(n_557), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g624 ( .A(n_557), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_557), .B(n_618), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_557), .B(n_614), .Y(n_640) );
AND2x2_ASAP7_75t_L g644 ( .A(n_557), .B(n_626), .Y(n_644) );
INVxp67_ASAP7_75t_L g576 ( .A(n_559), .Y(n_576) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_561), .A2(n_634), .B1(n_639), .B2(n_640), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_561), .B(n_666), .Y(n_696) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g682 ( .A(n_562), .B(n_673), .Y(n_682) );
AND2x2_ASAP7_75t_L g711 ( .A(n_562), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g716 ( .A(n_562), .B(n_666), .Y(n_716) );
INVx1_ASAP7_75t_L g629 ( .A(n_563), .Y(n_629) );
BUFx2_ASAP7_75t_L g635 ( .A(n_563), .Y(n_635) );
INVx1_ASAP7_75t_L g720 ( .A(n_564), .Y(n_720) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_565), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_567), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_567), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
INVx3_ASAP7_75t_L g626 ( .A(n_567), .Y(n_626) );
OR2x2_ASAP7_75t_L g692 ( .A(n_567), .B(n_693), .Y(n_692) );
AOI211xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_574), .B(n_577), .C(n_589), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_570), .A2(n_707), .B1(n_714), .B2(n_716), .C(n_717), .Y(n_706) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_578), .B(n_584), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_580), .B(n_618), .Y(n_632) );
AND2x2_ASAP7_75t_L g674 ( .A(n_580), .B(n_614), .Y(n_674) );
INVx1_ASAP7_75t_SL g687 ( .A(n_581), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_581), .B(n_635), .Y(n_690) );
INVx1_ASAP7_75t_L g708 ( .A(n_582), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_586), .A2(n_676), .B1(n_678), .B2(n_682), .C(n_683), .Y(n_675) );
AND2x2_ASAP7_75t_L g702 ( .A(n_587), .B(n_694), .Y(n_702) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g686 ( .A(n_588), .Y(n_686) );
AOI21xp33_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_593), .B(n_594), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g657 ( .A(n_592), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g643 ( .A(n_593), .Y(n_643) );
INVx1_ASAP7_75t_L g671 ( .A(n_594), .Y(n_671) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_602), .C(n_605), .Y(n_597) );
OAI31xp33_ASAP7_75t_L g724 ( .A1(n_598), .A2(n_636), .A3(n_723), .B(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g698 ( .A(n_601), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g719 ( .A(n_601), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_603), .B(n_618), .Y(n_646) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g721 ( .A(n_604), .B(n_618), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_613), .B1(n_617), .B2(n_620), .Y(n_608) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_612), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g648 ( .A(n_612), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_612), .B(n_635), .Y(n_651) );
AND2x2_ASAP7_75t_L g705 ( .A(n_612), .B(n_700), .Y(n_705) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g680 ( .A(n_616), .Y(n_680) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OAI32xp33_ASAP7_75t_L g683 ( .A1(n_618), .A2(n_652), .A3(n_684), .B1(n_686), .B2(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g658 ( .A(n_621), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_621), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g681 ( .A(n_625), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B(n_631), .C(n_633), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_629), .B(n_666), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_630), .A2(n_642), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g642 ( .A(n_640), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_650), .B2(n_652), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_650), .B(n_708), .C(n_709), .D(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NAND4xp25_ASAP7_75t_SL g654 ( .A(n_655), .B(n_668), .C(n_675), .D(n_688), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B(n_663), .C(n_664), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g685 ( .A(n_661), .Y(n_685) );
INVx2_ASAP7_75t_L g709 ( .A(n_666), .Y(n_709) );
OR2x2_ASAP7_75t_L g718 ( .A(n_673), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_695), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g714 ( .A(n_694), .B(n_715), .Y(n_714) );
AOI21xp33_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_697), .B(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
CKINVDCx16_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g733 ( .A(n_726), .Y(n_733) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_SL g753 ( .A(n_741), .Y(n_753) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_745), .B(n_750), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g757 ( .A(n_751), .Y(n_757) );
BUFx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
endmodule