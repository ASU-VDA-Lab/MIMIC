module fake_jpeg_1835_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_12),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_14),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_53),
.B(n_61),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_53),
.Y(n_99)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_96),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_57),
.B1(n_77),
.B2(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_55),
.B1(n_75),
.B2(n_72),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_64),
.B(n_63),
.C(n_59),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_116),
.B1(n_110),
.B2(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_67),
.B1(n_56),
.B2(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_67),
.B1(n_75),
.B2(n_73),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_57),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_59),
.B1(n_56),
.B2(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_124),
.B1(n_131),
.B2(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_129),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_127),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_136),
.B1(n_0),
.B2(n_1),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_132),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_73),
.B1(n_51),
.B2(n_52),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_2),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_51),
.B1(n_54),
.B2(n_66),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_8),
.Y(n_174)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_110),
.C(n_109),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_149),
.C(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_155),
.C(n_7),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_54),
.B(n_68),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_161),
.B(n_6),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_154),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_48),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_0),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_46),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_42),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_41),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_160),
.C(n_6),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_118),
.C(n_128),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_40),
.C(n_37),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_3),
.B(n_5),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_36),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_33),
.B(n_32),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_172),
.B(n_12),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_174),
.B1(n_179),
.B2(n_10),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_31),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_181),
.B(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_188),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_158),
.B(n_139),
.C(n_156),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_184),
.B(n_171),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_159),
.B(n_160),
.C(n_13),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_30),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_178),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_177),
.C(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_194),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_198),
.B1(n_163),
.B2(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_168),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_199),
.B1(n_180),
.B2(n_184),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_174),
.B1(n_166),
.B2(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_189),
.C(n_166),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_204),
.B1(n_193),
.B2(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_205),
.C(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_206),
.A3(n_201),
.B1(n_186),
.B2(n_29),
.C1(n_28),
.C2(n_22),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_211),
.B(n_13),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_16),
.B(n_18),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_19),
.Y(n_215)
);


endmodule