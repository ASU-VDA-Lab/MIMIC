module fake_jpeg_6982_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_41),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_12),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_27),
.B1(n_28),
.B2(n_17),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_50),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_63),
.Y(n_73)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_30),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_31),
.B(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_29),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_45),
.B1(n_65),
.B2(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_33),
.B(n_27),
.C(n_24),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_81),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_87),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_17),
.B(n_39),
.C(n_42),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_39),
.B1(n_24),
.B2(n_32),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_86),
.B1(n_47),
.B2(n_45),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_28),
.B1(n_23),
.B2(n_36),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_39),
.B1(n_32),
.B2(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_68),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_42),
.C(n_31),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_42),
.B1(n_31),
.B2(n_22),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_65),
.B1(n_46),
.B2(n_59),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_26),
.B(n_83),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_56),
.C(n_51),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_103),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_65),
.B1(n_56),
.B2(n_62),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_77),
.B1(n_70),
.B2(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_121),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_113),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_69),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_66),
.B1(n_46),
.B2(n_67),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_19),
.B(n_31),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_67),
.B1(n_20),
.B2(n_21),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_81),
.B1(n_83),
.B2(n_72),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_46),
.B1(n_22),
.B2(n_21),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_82),
.B1(n_88),
.B2(n_78),
.Y(n_138)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_72),
.B(n_57),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_138),
.B1(n_81),
.B2(n_96),
.Y(n_181)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_130),
.Y(n_159)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_132),
.Y(n_167)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_136),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_89),
.B(n_93),
.C(n_94),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_123),
.B(n_119),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_75),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_75),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_137),
.B(n_143),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_82),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_145),
.Y(n_172)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_148),
.Y(n_182)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_151),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_82),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_97),
.C(n_122),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_168),
.C(n_142),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_158),
.B(n_163),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_97),
.C(n_106),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_160),
.B(n_162),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_106),
.B(n_114),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_174),
.B(n_175),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_113),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_111),
.B1(n_101),
.B2(n_120),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_151),
.B1(n_139),
.B2(n_140),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_127),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_126),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_103),
.B1(n_106),
.B2(n_115),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_181),
.B1(n_144),
.B2(n_90),
.Y(n_206)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_107),
.A3(n_116),
.B1(n_96),
.B2(n_98),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_135),
.B(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_90),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_178),
.B(n_124),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_184),
.A2(n_193),
.B(n_183),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_197),
.B(n_187),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_190),
.C(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_202),
.B1(n_208),
.B2(n_157),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_162),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_146),
.C(n_140),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_164),
.A3(n_166),
.B1(n_169),
.B2(n_160),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_209),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_138),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_78),
.C(n_133),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_135),
.C(n_68),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_198),
.C(n_207),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_135),
.B(n_90),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_135),
.C(n_68),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_148),
.B1(n_145),
.B2(n_129),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_76),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_210),
.B1(n_180),
.B2(n_182),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_64),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_94),
.B1(n_20),
.B2(n_21),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_68),
.C(n_64),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_21),
.B1(n_20),
.B2(n_64),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_184),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_177),
.C(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_197),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_177),
.B1(n_180),
.B2(n_154),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_219),
.B1(n_223),
.B2(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_185),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_224),
.B1(n_34),
.B2(n_1),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_155),
.B(n_163),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_153),
.B1(n_172),
.B2(n_176),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_25),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_234),
.B1(n_211),
.B2(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_0),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_34),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_238),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_189),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_186),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_205),
.C(n_190),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_251),
.C(n_233),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_194),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_249),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_216),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_208),
.C(n_34),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_218),
.B1(n_212),
.B2(n_224),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_259),
.B1(n_269),
.B2(n_271),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_9),
.CI(n_15),
.CON(n_280),
.SN(n_280)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_218),
.B1(n_219),
.B2(n_225),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_270),
.C(n_245),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_265),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_233),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_242),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_223),
.C(n_227),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_214),
.B1(n_234),
.B2(n_229),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_259),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_244),
.B(n_236),
.C(n_249),
.D(n_241),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_280),
.C(n_267),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_251),
.B1(n_234),
.B2(n_250),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_284),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_281),
.C(n_10),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_248),
.C(n_1),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_283),
.C(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_0),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_12),
.B(n_16),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_2),
.C(n_3),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_291),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_11),
.C(n_14),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_288),
.B(n_289),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_282),
.B1(n_263),
.B2(n_284),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_260),
.B(n_267),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.C(n_295),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_9),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_9),
.B(n_14),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_276),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_301),
.B(n_303),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_283),
.C(n_274),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_16),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_280),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_7),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_310),
.B(n_13),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_309),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_8),
.B(n_11),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_12),
.B(n_13),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_13),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_311),
.B1(n_6),
.B2(n_308),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_6),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_299),
.Y(n_317)
);


endmodule