module fake_ibex_457_n_907 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_907);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_907;

wire n_151;
wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_141;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_841;
wire n_679;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_148;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_794;
wire n_260;
wire n_620;
wire n_836;
wire n_683;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_895;
wire n_687;
wire n_202;
wire n_231;
wire n_159;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_73),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_41),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_49),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_14),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_48),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_52),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_70),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_29),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_57),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_83),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_42),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_11),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_60),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_22),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_51),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_38),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_67),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_106),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_100),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_56),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_44),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_63),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_43),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_109),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_91),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_75),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_58),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_34),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_50),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_46),
.B(n_77),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_104),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_125),
.Y(n_204)
);

BUFx8_ASAP7_75t_SL g205 ( 
.A(n_40),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_37),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_105),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_47),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_78),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_32),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_11),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_69),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_53),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_6),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_107),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_25),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_82),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_124),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_98),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_80),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_15),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_31),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_22),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_101),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_10),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_66),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_110),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_89),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_118),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_55),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_85),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_147),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_142),
.A2(n_61),
.B(n_137),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_162),
.B(n_3),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_4),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_7),
.Y(n_259)
);

CKINVDCx6p67_ASAP7_75t_R g260 ( 
.A(n_202),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_9),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_142),
.A2(n_62),
.B(n_132),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_173),
.B(n_196),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_165),
.B(n_211),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_9),
.Y(n_267)
);

CKINVDCx11_ASAP7_75t_R g268 ( 
.A(n_143),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_161),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_141),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_155),
.Y(n_275)
);

CKINVDCx11_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_146),
.Y(n_277)
);

BUFx8_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_12),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_151),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_149),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_209),
.B(n_13),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_170),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_172),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_154),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_160),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_224),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_170),
.B(n_39),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_245),
.B(n_145),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_145),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_246),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_155),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_150),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_152),
.A2(n_72),
.B(n_119),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_195),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_205),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_175),
.B(n_16),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_152),
.B(n_16),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_167),
.Y(n_307)
);

BUFx8_ASAP7_75t_SL g308 ( 
.A(n_225),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_167),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_175),
.B(n_17),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_153),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_185),
.B(n_17),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_197),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_185),
.B(n_18),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_157),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_159),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_176),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_197),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_192),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_178),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_166),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_197),
.Y(n_323)
);

CKINVDCx11_ASAP7_75t_R g324 ( 
.A(n_193),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_191),
.B(n_24),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_212),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_218),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_169),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_168),
.B(n_26),
.Y(n_330)
);

AOI22x1_ASAP7_75t_SL g331 ( 
.A1(n_193),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_226),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_250),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_252),
.B(n_235),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_251),
.B(n_174),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_249),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_194),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_251),
.B(n_177),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_194),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_251),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_274),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_256),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_256),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_206),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_299),
.Y(n_364)
);

BUFx6f_ASAP7_75t_SL g365 ( 
.A(n_257),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_261),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_265),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_277),
.B(n_180),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_265),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_265),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_286),
.B(n_280),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_258),
.B(n_215),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_300),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_265),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_300),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_266),
.B(n_181),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_304),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_302),
.B(n_290),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_263),
.B(n_182),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_254),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_296),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_254),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_309),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_271),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_296),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_294),
.B(n_184),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_294),
.B(n_189),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_271),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_298),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_263),
.B(n_183),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_285),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_283),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_302),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_311),
.B(n_315),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_283),
.Y(n_402)
);

AO21x2_ASAP7_75t_L g403 ( 
.A1(n_255),
.A2(n_262),
.B(n_306),
.Y(n_403)
);

NOR2x1p5_ASAP7_75t_L g404 ( 
.A(n_260),
.B(n_200),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_291),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_305),
.Y(n_411)
);

AO21x2_ASAP7_75t_L g412 ( 
.A1(n_330),
.A2(n_222),
.B(n_244),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_314),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

AO22x2_ASAP7_75t_L g418 ( 
.A1(n_331),
.A2(n_241),
.B1(n_240),
.B2(n_239),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_292),
.B(n_188),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_267),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_319),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_303),
.B(n_190),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_325),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_272),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_326),
.B(n_216),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_293),
.B(n_198),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_287),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_293),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_328),
.Y(n_434)
);

AND3x2_ASAP7_75t_L g435 ( 
.A(n_324),
.B(n_223),
.C(n_227),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_272),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_320),
.Y(n_437)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_372),
.B(n_276),
.C(n_268),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_363),
.A2(n_279),
.B1(n_248),
.B2(n_329),
.Y(n_443)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_436),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_374),
.B(n_281),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g446 ( 
.A(n_372),
.B(n_276),
.C(n_268),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_348),
.B(n_281),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_334),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_282),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_344),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_363),
.B(n_282),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_345),
.B(n_322),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_433),
.B(n_329),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_324),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_199),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_374),
.B(n_158),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_301),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_342),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_374),
.B(n_163),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_342),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_373),
.B(n_233),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_207),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_342),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_R g469 ( 
.A(n_381),
.B(n_297),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_340),
.B(n_316),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_347),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_179),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_413),
.B(n_201),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_347),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_396),
.B(n_204),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_344),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_430),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_347),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_333),
.B(n_247),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_SL g482 ( 
.A(n_340),
.B(n_233),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_373),
.B(n_430),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_428),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_344),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_356),
.B(n_208),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_356),
.B(n_210),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_366),
.B(n_213),
.Y(n_488)
);

AOI221xp5_ASAP7_75t_L g489 ( 
.A1(n_337),
.A2(n_392),
.B1(n_393),
.B2(n_401),
.C(n_418),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_339),
.A2(n_367),
.B1(n_402),
.B2(n_398),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_335),
.B(n_219),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_428),
.B(n_308),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_419),
.B(n_424),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_420),
.B(n_220),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_351),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_332),
.B(n_217),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_420),
.B(n_238),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_332),
.B(n_229),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_341),
.B(n_230),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_341),
.B(n_242),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_353),
.B(n_243),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_353),
.B(n_187),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_360),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_436),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_404),
.B(n_418),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_369),
.B(n_387),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_381),
.B(n_308),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_361),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_361),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_351),
.B(n_186),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_352),
.B(n_187),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_364),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_364),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_375),
.Y(n_515)
);

NAND2x1_ASAP7_75t_L g516 ( 
.A(n_377),
.B(n_275),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_377),
.Y(n_517)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_431),
.B(n_30),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_354),
.B(n_87),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_462),
.A2(n_403),
.B(n_354),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_493),
.B(n_378),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_462),
.A2(n_403),
.B(n_379),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_454),
.B(n_365),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_448),
.B(n_365),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_514),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_403),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_483),
.B(n_380),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_478),
.B(n_380),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_466),
.B(n_383),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_448),
.B(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_463),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_465),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_501),
.A2(n_350),
.B(n_338),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_452),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_468),
.Y(n_538)
);

A2O1A1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_489),
.A2(n_422),
.B(n_390),
.C(n_388),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_518),
.A2(n_422),
.B1(n_390),
.B2(n_388),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_461),
.B(n_405),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

NOR3xp33_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_336),
.C(n_346),
.Y(n_543)
);

OR2x6_ASAP7_75t_SL g544 ( 
.A(n_492),
.B(n_405),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_444),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_451),
.B(n_415),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_464),
.B(n_415),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_502),
.B(n_481),
.Y(n_548)
);

NOR2x1p5_ASAP7_75t_L g549 ( 
.A(n_508),
.B(n_33),
.Y(n_549)
);

AO21x1_ASAP7_75t_L g550 ( 
.A1(n_519),
.A2(n_512),
.B(n_503),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_447),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_512),
.A2(n_349),
.B(n_343),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_440),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_471),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_467),
.B(n_432),
.Y(n_555)
);

BUFx4f_ASAP7_75t_L g556 ( 
.A(n_505),
.Y(n_556)
);

NOR2x1_ASAP7_75t_L g557 ( 
.A(n_457),
.B(n_355),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_484),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_441),
.Y(n_560)
);

NOR2x1_ASAP7_75t_L g561 ( 
.A(n_445),
.B(n_355),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_507),
.A2(n_487),
.B(n_486),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_455),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_496),
.A2(n_429),
.B(n_427),
.C(n_426),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_476),
.B(n_358),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_491),
.B(n_35),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_474),
.B(n_479),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_504),
.A2(n_362),
.B(n_427),
.C(n_426),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_506),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_456),
.B(n_36),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_497),
.A2(n_359),
.B1(n_423),
.B2(n_421),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_486),
.A2(n_358),
.B(n_421),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_509),
.A2(n_399),
.B(n_417),
.C(n_416),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_487),
.A2(n_399),
.B(n_417),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_437),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_510),
.Y(n_577)
);

AO21x1_ASAP7_75t_L g578 ( 
.A1(n_497),
.A2(n_395),
.B(n_371),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_513),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_488),
.B(n_36),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_470),
.A2(n_370),
.B1(n_414),
.B2(n_410),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_488),
.B(n_37),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_485),
.B(n_368),
.Y(n_583)
);

A2O1A1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_515),
.A2(n_391),
.B(n_409),
.C(n_408),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_450),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_453),
.B(n_45),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_495),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_517),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_499),
.B(n_500),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_459),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_500),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_480),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_443),
.A2(n_386),
.B1(n_376),
.B2(n_407),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_516),
.Y(n_595)
);

OR2x6_ASAP7_75t_SL g596 ( 
.A(n_469),
.B(n_65),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_438),
.C(n_446),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_523),
.A2(n_589),
.B(n_562),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_522),
.B(n_472),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_576),
.B(n_506),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_591),
.B(n_475),
.Y(n_602)
);

OAI22x1_ASAP7_75t_L g603 ( 
.A1(n_549),
.A2(n_494),
.B1(n_498),
.B2(n_511),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_546),
.B(n_460),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_534),
.A2(n_539),
.B(n_552),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_530),
.B(n_473),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_545),
.B(n_458),
.Y(n_608)
);

INVx3_ASAP7_75t_SL g609 ( 
.A(n_559),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_545),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_556),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_528),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_529),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_579),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_588),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_524),
.A2(n_531),
.B1(n_586),
.B2(n_570),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_544),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_556),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_580),
.A2(n_582),
.B(n_541),
.C(n_547),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_537),
.B(n_434),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_596),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_533),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_537),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_571),
.B(n_567),
.Y(n_625)
);

OA22x2_ASAP7_75t_L g626 ( 
.A1(n_538),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_568),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_555),
.B(n_99),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_554),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_520),
.A2(n_543),
.B1(n_581),
.B2(n_526),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_558),
.B(n_108),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_595),
.B(n_113),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_564),
.B(n_115),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_564),
.B(n_140),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_560),
.B(n_593),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_587),
.B(n_592),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_561),
.B(n_595),
.Y(n_638)
);

AO31x2_ASAP7_75t_L g639 ( 
.A1(n_572),
.A2(n_594),
.A3(n_584),
.B(n_569),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_563),
.Y(n_640)
);

CKINVDCx14_ASAP7_75t_R g641 ( 
.A(n_594),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g642 ( 
.A(n_595),
.B(n_566),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_557),
.Y(n_643)
);

AO31x2_ASAP7_75t_L g644 ( 
.A1(n_565),
.A2(n_574),
.A3(n_575),
.B(n_573),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_585),
.Y(n_645)
);

OAI21xp33_ASAP7_75t_L g646 ( 
.A1(n_583),
.A2(n_548),
.B(n_449),
.Y(n_646)
);

AO31x2_ASAP7_75t_L g647 ( 
.A1(n_550),
.A2(n_578),
.A3(n_527),
.B(n_521),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_542),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_542),
.B(n_545),
.Y(n_649)
);

AND3x1_ASAP7_75t_SL g650 ( 
.A(n_549),
.B(n_489),
.C(n_404),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_536),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_542),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_522),
.B(n_591),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_522),
.B(n_591),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_521),
.A2(n_431),
.B(n_523),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_559),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_522),
.B(n_591),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_577),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_559),
.A2(n_506),
.B1(n_449),
.B2(n_143),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_521),
.A2(n_431),
.B(n_523),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_535),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_521),
.A2(n_431),
.B(n_523),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_542),
.B(n_545),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_577),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_576),
.B(n_483),
.Y(n_665)
);

OAI21xp33_ASAP7_75t_SL g666 ( 
.A1(n_589),
.A2(n_518),
.B(n_540),
.Y(n_666)
);

AO22x1_ASAP7_75t_L g667 ( 
.A1(n_576),
.A2(n_446),
.B1(n_438),
.B2(n_320),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_542),
.B(n_444),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_576),
.B(n_483),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_562),
.A2(n_548),
.B(n_591),
.C(n_589),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_577),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_654),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_612),
.B(n_602),
.Y(n_674)
);

BUFx2_ASAP7_75t_SL g675 ( 
.A(n_656),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_655),
.A2(n_662),
.B(n_660),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_665),
.B(n_670),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_657),
.Y(n_678)
);

BUFx2_ASAP7_75t_R g679 ( 
.A(n_609),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_615),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_669),
.B(n_607),
.Y(n_681)
);

INVx8_ASAP7_75t_L g682 ( 
.A(n_668),
.Y(n_682)
);

BUFx2_ASAP7_75t_SL g683 ( 
.A(n_611),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_627),
.B(n_668),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_613),
.B(n_600),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_SL g686 ( 
.A1(n_626),
.A2(n_627),
.B(n_628),
.Y(n_686)
);

NOR2x1_ASAP7_75t_SL g687 ( 
.A(n_648),
.B(n_652),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_614),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_648),
.B(n_652),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_597),
.B(n_648),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_621),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_649),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_652),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_649),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_619),
.A2(n_671),
.B(n_605),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_663),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_663),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_641),
.A2(n_659),
.B1(n_617),
.B2(n_666),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_625),
.B(n_598),
.C(n_646),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_661),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_610),
.Y(n_702)
);

OAI21x1_ASAP7_75t_SL g703 ( 
.A1(n_604),
.A2(n_634),
.B(n_664),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_658),
.B(n_672),
.Y(n_704)
);

AND2x4_ASAP7_75t_SL g705 ( 
.A(n_618),
.B(n_651),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_664),
.B(n_672),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_606),
.A2(n_630),
.B(n_629),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_629),
.B(n_622),
.Y(n_708)
);

INVxp33_ASAP7_75t_L g709 ( 
.A(n_601),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_616),
.B(n_623),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_632),
.A2(n_635),
.B(n_636),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_667),
.B(n_608),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_645),
.B(n_640),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_647),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_642),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_603),
.B(n_643),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_638),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_637),
.B(n_631),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_647),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_644),
.A2(n_620),
.B(n_639),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_638),
.Y(n_721)
);

OA21x2_ASAP7_75t_L g722 ( 
.A1(n_639),
.A2(n_644),
.B(n_633),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_650),
.B(n_638),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_653),
.B(n_654),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_624),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_653),
.B(n_654),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_653),
.B(n_654),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_597),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_653),
.B(n_654),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_612),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_648),
.B(n_545),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_612),
.B(n_665),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_612),
.B(n_470),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_648),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_671),
.A2(n_599),
.B(n_619),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_612),
.B(n_470),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_671),
.A2(n_599),
.B(n_619),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_688),
.Y(n_738)
);

INVx6_ASAP7_75t_L g739 ( 
.A(n_697),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_688),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_704),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_702),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_698),
.A2(n_727),
.B1(n_724),
.B2(n_729),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_682),
.A2(n_684),
.B1(n_697),
.B2(n_703),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_698),
.A2(n_710),
.B1(n_700),
.B2(n_685),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_727),
.A2(n_673),
.B1(n_729),
.B2(n_724),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_678),
.B(n_673),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_678),
.B(n_726),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_708),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_726),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_708),
.Y(n_752)
);

NOR2x1p5_ASAP7_75t_L g753 ( 
.A(n_693),
.B(n_717),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_706),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_680),
.Y(n_755)
);

AOI221xp5_ASAP7_75t_L g756 ( 
.A1(n_685),
.A2(n_674),
.B1(n_710),
.B2(n_736),
.C(n_733),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_702),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_718),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_714),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_728),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_714),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_707),
.B(n_674),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_707),
.B(n_732),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_719),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_694),
.B(n_701),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_713),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_735),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_735),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_684),
.B(n_677),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_728),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_682),
.Y(n_772)
);

INVx6_ASAP7_75t_L g773 ( 
.A(n_699),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_690),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_737),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_733),
.A2(n_736),
.B1(n_723),
.B2(n_709),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_675),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_730),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_692),
.B(n_696),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_695),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_771),
.B(n_681),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_746),
.A2(n_723),
.B1(n_709),
.B2(n_716),
.Y(n_783)
);

OAI222xp33_ASAP7_75t_L g784 ( 
.A1(n_743),
.A2(n_712),
.B1(n_716),
.B2(n_691),
.C1(n_731),
.C2(n_721),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_749),
.B(n_722),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_742),
.B(n_695),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_742),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_741),
.B(n_745),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_741),
.B(n_686),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_759),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_776),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_767),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_776),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_762),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_757),
.B(n_722),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_SL g796 ( 
.A1(n_744),
.A2(n_689),
.B(n_715),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_759),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_768),
.B(n_720),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_749),
.B(n_722),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_738),
.B(n_740),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_757),
.Y(n_801)
);

BUFx8_ASAP7_75t_L g802 ( 
.A(n_758),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_750),
.B(n_752),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_763),
.B(n_689),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_747),
.A2(n_712),
.B1(n_711),
.B2(n_716),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_771),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_748),
.B(n_693),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_740),
.B(n_676),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_770),
.B(n_691),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_751),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_792),
.B(n_763),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_800),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_800),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_790),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_810),
.B(n_764),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_785),
.B(n_769),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_785),
.B(n_769),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_790),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_799),
.B(n_775),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_787),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_797),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_799),
.B(n_775),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_803),
.B(n_764),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_805),
.A2(n_777),
.B1(n_712),
.B2(n_748),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_808),
.B(n_781),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_803),
.B(n_755),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_794),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_788),
.B(n_755),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_801),
.B(n_781),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_805),
.A2(n_739),
.B1(n_756),
.B2(n_766),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_801),
.B(n_765),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_817),
.B(n_808),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_818),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_827),
.Y(n_834)
);

OAI221xp5_ASAP7_75t_L g835 ( 
.A1(n_830),
.A2(n_783),
.B1(n_796),
.B2(n_782),
.C(n_774),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_815),
.B(n_786),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_820),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_812),
.B(n_789),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_811),
.B(n_786),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_827),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_818),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_813),
.B(n_804),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_821),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_816),
.B(n_798),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_831),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_816),
.B(n_798),
.Y(n_846)
);

INVxp67_ASAP7_75t_SL g847 ( 
.A(n_831),
.Y(n_847)
);

OAI211xp5_ASAP7_75t_L g848 ( 
.A1(n_835),
.A2(n_796),
.B(n_806),
.C(n_772),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_844),
.B(n_822),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_837),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_836),
.B(n_822),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_834),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_836),
.B(n_817),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_839),
.B(n_817),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_839),
.B(n_819),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_841),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_845),
.B(n_819),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_834),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_832),
.B(n_819),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_847),
.B(n_829),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_840),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_850),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_856),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_860),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_848),
.A2(n_784),
.B(n_809),
.Y(n_865)
);

OAI33xp33_ASAP7_75t_L g866 ( 
.A1(n_857),
.A2(n_838),
.A3(n_824),
.B1(n_842),
.B2(n_823),
.B3(n_828),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_849),
.B(n_846),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_851),
.B(n_846),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_848),
.A2(n_832),
.B1(n_844),
.B2(n_825),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_854),
.Y(n_870)
);

NOR3xp33_ASAP7_75t_L g871 ( 
.A(n_856),
.B(n_779),
.C(n_766),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_855),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_859),
.B(n_832),
.Y(n_873)
);

OAI321xp33_ASAP7_75t_L g874 ( 
.A1(n_865),
.A2(n_869),
.A3(n_873),
.B1(n_866),
.B2(n_853),
.C(n_863),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_873),
.A2(n_859),
.B1(n_778),
.B2(n_793),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_862),
.B(n_861),
.C(n_858),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_863),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_864),
.A2(n_825),
.B1(n_833),
.B2(n_861),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_871),
.A2(n_760),
.B(n_789),
.C(n_770),
.Y(n_879)
);

OAI332xp33_ASAP7_75t_L g880 ( 
.A1(n_870),
.A2(n_826),
.A3(n_679),
.B1(n_829),
.B2(n_852),
.B3(n_788),
.C1(n_821),
.C2(n_795),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_SL g881 ( 
.A1(n_875),
.A2(n_868),
.B(n_867),
.C(n_872),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_874),
.B(n_679),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_878),
.B(n_843),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_876),
.Y(n_884)
);

CKINVDCx16_ASAP7_75t_R g885 ( 
.A(n_879),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_877),
.A2(n_843),
.B1(n_841),
.B2(n_802),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_884),
.B(n_880),
.Y(n_887)
);

NAND4xp75_ASAP7_75t_L g888 ( 
.A(n_882),
.B(n_734),
.C(n_791),
.D(n_780),
.Y(n_888)
);

OAI321xp33_ASAP7_75t_L g889 ( 
.A1(n_886),
.A2(n_791),
.A3(n_795),
.B1(n_807),
.B2(n_814),
.C(n_758),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_885),
.B(n_683),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_887),
.B(n_881),
.C(n_883),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_890),
.Y(n_892)
);

NOR3x1_ASAP7_75t_L g893 ( 
.A(n_888),
.B(n_761),
.C(n_772),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_889),
.B(n_802),
.C(n_699),
.Y(n_894)
);

NOR2x1_ASAP7_75t_L g895 ( 
.A(n_892),
.B(n_753),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_893),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_896),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_895),
.B(n_891),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_897),
.Y(n_899)
);

XOR2x1_ASAP7_75t_L g900 ( 
.A(n_899),
.B(n_898),
.Y(n_900)
);

OAI331xp33_ASAP7_75t_L g901 ( 
.A1(n_900),
.A2(n_682),
.A3(n_894),
.B1(n_772),
.B2(n_687),
.B3(n_754),
.C1(n_752),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_SL g902 ( 
.A1(n_901),
.A2(n_773),
.B1(n_772),
.B2(n_739),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_902),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_SL g904 ( 
.A1(n_903),
.A2(n_705),
.B(n_772),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_904),
.B(n_699),
.C(n_725),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_905),
.B(n_773),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_906),
.A2(n_773),
.B1(n_739),
.B2(n_753),
.Y(n_907)
);


endmodule