module fake_jpeg_2220_n_371 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_51),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_52),
.B(n_65),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_67),
.Y(n_103)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_64),
.B(n_71),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_2),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_2),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_85),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_6),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_99),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_90),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_96),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_6),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

NAND2x1_ASAP7_75t_SL g99 ( 
.A(n_46),
.B(n_7),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_41),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_52),
.B1(n_65),
.B2(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_106),
.A2(n_115),
.B1(n_160),
.B2(n_126),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_47),
.A2(n_41),
.B1(n_40),
.B2(n_29),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_128),
.B1(n_155),
.B2(n_136),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_40),
.B1(n_29),
.B2(n_25),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_25),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_120),
.B(n_131),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_148),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_49),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_97),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_8),
.B(n_9),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_158),
.B(n_144),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_59),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_159),
.B1(n_141),
.B2(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_14),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_50),
.A2(n_16),
.B1(n_60),
.B2(n_69),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_89),
.A2(n_99),
.B(n_93),
.C(n_98),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_94),
.A2(n_70),
.B1(n_35),
.B2(n_82),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_76),
.A2(n_64),
.B1(n_71),
.B2(n_96),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_162),
.Y(n_212)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_189),
.B(n_191),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_113),
.A2(n_151),
.B1(n_114),
.B2(n_111),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_192),
.B1(n_174),
.B2(n_179),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_195),
.B1(n_201),
.B2(n_186),
.Y(n_226)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_193),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_147),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_181),
.Y(n_205)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_101),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_104),
.A2(n_119),
.B1(n_129),
.B2(n_158),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_188),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_157),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_202),
.Y(n_220)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_105),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_117),
.A2(n_143),
.B1(n_132),
.B2(n_152),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_108),
.B(n_153),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_124),
.B1(n_146),
.B2(n_137),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_143),
.Y(n_193)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_124),
.B1(n_133),
.B2(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_198),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_190),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_146),
.A2(n_126),
.B1(n_141),
.B2(n_125),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_125),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_185),
.B(n_188),
.C(n_168),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_195),
.B(n_202),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_228),
.B1(n_201),
.B2(n_182),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_199),
.B1(n_181),
.B2(n_163),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_167),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_231),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_181),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_232),
.A2(n_227),
.B(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_237),
.A2(n_205),
.B1(n_223),
.B2(n_213),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_238),
.B(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_164),
.C(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_175),
.Y(n_241)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_170),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_178),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_180),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_187),
.C(n_166),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_202),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_194),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_261),
.B(n_274),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_229),
.B(n_225),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_271),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI221xp5_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_228),
.B1(n_225),
.B2(n_213),
.C(n_208),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_246),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_225),
.B(n_206),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_242),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_229),
.B1(n_227),
.B2(n_205),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_275),
.B1(n_240),
.B2(n_237),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_213),
.B(n_205),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_285),
.B1(n_290),
.B2(n_237),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_239),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_286),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_249),
.B(n_236),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_293),
.B(n_262),
.Y(n_310)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_231),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_239),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_248),
.C(n_268),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_230),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_264),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_240),
.B1(n_271),
.B2(n_255),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_254),
.A2(n_235),
.B(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_304),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_308),
.C(n_272),
.Y(n_314)
);

OAI221xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_269),
.B1(n_270),
.B2(n_268),
.C(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_280),
.B1(n_276),
.B2(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_311),
.B1(n_283),
.B2(n_277),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_265),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_303),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_287),
.B(n_274),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_310),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_248),
.C(n_263),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_276),
.A2(n_271),
.B1(n_275),
.B2(n_255),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_285),
.B1(n_262),
.B2(n_273),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_277),
.A2(n_271),
.B(n_273),
.C(n_259),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_310),
.B1(n_311),
.B2(n_308),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_307),
.C(n_306),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_246),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_324),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_294),
.B1(n_284),
.B2(n_279),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_325),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_217),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_319),
.B(n_244),
.Y(n_332)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_241),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_314),
.B1(n_320),
.B2(n_324),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_316),
.C(n_320),
.Y(n_339)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_313),
.A2(n_302),
.B(n_311),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_334),
.A2(n_311),
.B(n_322),
.Y(n_337)
);

NAND4xp25_ASAP7_75t_SL g335 ( 
.A(n_322),
.B(n_243),
.C(n_259),
.D(n_241),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_330),
.B(n_318),
.CI(n_315),
.CON(n_336),
.SN(n_336)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_337),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_327),
.B1(n_335),
.B2(n_281),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_341),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_312),
.B1(n_296),
.B2(n_305),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_342),
.A2(n_343),
.B1(n_267),
.B2(n_258),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_317),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_341),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_347),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_327),
.C(n_334),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_348),
.B(n_336),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_350),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_343),
.B(n_258),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_351),
.B(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_353),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_337),
.C(n_340),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_356),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_346),
.B(n_336),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_357),
.A2(n_250),
.B(n_234),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g359 ( 
.A(n_358),
.B(n_352),
.CI(n_349),
.CON(n_359),
.SN(n_359)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_361),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_355),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_355),
.B(n_247),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_243),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_363),
.A2(n_245),
.B(n_215),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_360),
.B(n_259),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_367),
.B(n_368),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_369),
.B(n_365),
.C(n_215),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_211),
.Y(n_371)
);


endmodule