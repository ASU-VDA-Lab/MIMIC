module fake_jpeg_18018_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

AND2x6_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_5),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_22),
.C(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_32),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_9),
.C(n_11),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_27),
.C(n_26),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_11),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

AOI322xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_3),
.A3(n_4),
.B1(n_12),
.B2(n_23),
.C1(n_28),
.C2(n_31),
.Y(n_35)
);

BUFx24_ASAP7_75t_SL g42 ( 
.A(n_35),
.Y(n_42)
);

OAI21x1_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_38),
.B(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_39),
.A3(n_38),
.B1(n_36),
.B2(n_26),
.C1(n_33),
.C2(n_34),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_42),
.B(n_43),
.Y(n_45)
);


endmodule