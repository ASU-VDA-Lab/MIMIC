module fake_netlist_5_1731_n_107 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_107);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_107;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx2_ASAP7_75t_SL g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_36),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_25),
.B(n_31),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_32),
.Y(n_54)
);

OR2x6_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_26),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_45),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_47),
.B(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_46),
.B(n_40),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_44),
.B1(n_33),
.B2(n_21),
.Y(n_60)
);

NOR4xp25_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_42),
.C(n_41),
.D(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_39),
.Y(n_62)
);

OA21x2_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_50),
.B(n_53),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_62),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_52),
.B(n_51),
.C(n_56),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_34),
.B1(n_55),
.B2(n_21),
.Y(n_67)
);

AOI21x1_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_52),
.B(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_55),
.B1(n_58),
.B2(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_63),
.B(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_73),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_69),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_63),
.B(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_39),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_76),
.B(n_68),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_86),
.C(n_87),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_37),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_38),
.C(n_37),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_1),
.B(n_3),
.Y(n_98)
);

NAND4xp75_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_1),
.C(n_5),
.D(n_6),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AOI222xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_101),
.B1(n_98),
.B2(n_100),
.C1(n_39),
.C2(n_7),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_103),
.B1(n_16),
.B2(n_68),
.Y(n_107)
);


endmodule