module fake_jpeg_17425_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_3),
.B(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_72),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_48),
.B1(n_43),
.B2(n_50),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_40),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_57),
.B1(n_46),
.B2(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_71),
.B1(n_79),
.B2(n_78),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_91),
.B1(n_96),
.B2(n_7),
.Y(n_103)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_95),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_107),
.B(n_10),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_105),
.B1(n_104),
.B2(n_108),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_85),
.B1(n_91),
.B2(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_114),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_94),
.B(n_92),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_17),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_109),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_12),
.B(n_13),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_19),
.Y(n_120)
);

AO21x2_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_106),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_20),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_124),
.C(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_125),
.B(n_25),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_23),
.B(n_26),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_29),
.B(n_30),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_32),
.B(n_33),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_34),
.Y(n_143)
);


endmodule