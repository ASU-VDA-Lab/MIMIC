module fake_jpeg_25500_n_300 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_12),
.B1(n_24),
.B2(n_14),
.Y(n_47)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_24),
.B1(n_14),
.B2(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_35),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_52),
.B1(n_32),
.B2(n_34),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_31),
.B1(n_47),
.B2(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_58),
.B1(n_63),
.B2(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_31),
.B1(n_33),
.B2(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_65),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_27),
.B1(n_12),
.B2(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_80),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_29),
.B(n_20),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_45),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_40),
.C(n_43),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_86),
.B1(n_87),
.B2(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_50),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_43),
.B1(n_40),
.B2(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_99),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_75),
.B1(n_32),
.B2(n_85),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_63),
.B1(n_48),
.B2(n_64),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_105),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_63),
.B1(n_59),
.B2(n_48),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_62),
.B1(n_60),
.B2(n_43),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_53),
.B1(n_61),
.B2(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_29),
.B1(n_34),
.B2(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_110),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_60),
.B(n_20),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_35),
.B1(n_20),
.B2(n_22),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_79),
.B1(n_71),
.B2(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_135),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_86),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_117),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_81),
.B1(n_69),
.B2(n_67),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_124),
.B1(n_128),
.B2(n_93),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_67),
.B1(n_74),
.B2(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_15),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_139),
.B(n_140),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_75),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_136),
.C(n_137),
.Y(n_147)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_15),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_35),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_89),
.A2(n_22),
.B(n_25),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_104),
.B1(n_94),
.B2(n_99),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_141),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_111),
.C(n_73),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_170),
.C(n_19),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_73),
.B(n_16),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_13),
.B1(n_16),
.B2(n_23),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_23),
.B(n_17),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_32),
.B1(n_22),
.B2(n_17),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_112),
.B1(n_113),
.B2(n_136),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_132),
.B(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_32),
.B1(n_22),
.B2(n_42),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_35),
.B1(n_13),
.B2(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_42),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_42),
.B1(n_35),
.B2(n_36),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_42),
.B1(n_36),
.B2(n_19),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_159),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_114),
.A2(n_13),
.B1(n_16),
.B2(n_23),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_19),
.C(n_21),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_17),
.B1(n_25),
.B2(n_15),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_30),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_199),
.B1(n_18),
.B2(n_7),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_19),
.C(n_21),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_191),
.C(n_197),
.Y(n_208)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_189),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_25),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_7),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_21),
.C(n_30),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_196),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_25),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_21),
.C(n_30),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_21),
.C(n_30),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_168),
.C(n_21),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_143),
.B1(n_160),
.B2(n_171),
.Y(n_199)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_15),
.B(n_6),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_169),
.B1(n_149),
.B2(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_172),
.B1(n_146),
.B2(n_154),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_154),
.B1(n_167),
.B2(n_151),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_170),
.B1(n_164),
.B2(n_165),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_152),
.B(n_156),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_212),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_200),
.B1(n_188),
.B2(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_191),
.C(n_186),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_182),
.C(n_197),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_18),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_224),
.C(n_231),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_208),
.C(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_226),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_181),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_180),
.CI(n_184),
.CON(n_229),
.SN(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_203),
.C(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_202),
.B1(n_209),
.B2(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_200),
.C(n_193),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_240),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_215),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_205),
.C(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_245),
.B1(n_254),
.B2(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_227),
.A2(n_214),
.B1(n_210),
.B2(n_2),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_247),
.Y(n_257)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_5),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_18),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_230),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_240),
.A2(n_238),
.B1(n_232),
.B2(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_225),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_4),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_224),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_266),
.B(n_249),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_223),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_5),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_8),
.B(n_11),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_8),
.B(n_11),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_250),
.C(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_270),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_250),
.C(n_258),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_273),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_8),
.B(n_10),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_4),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_8),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_284),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_3),
.B(n_9),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_0),
.B(n_1),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_18),
.B1(n_3),
.B2(n_9),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_285),
.A2(n_286),
.B(n_0),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_9),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_291),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_269),
.B(n_270),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_289),
.B(n_278),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_292),
.A2(n_287),
.B(n_282),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_271),
.C(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_18),
.C(n_1),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_296),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_18),
.C(n_1),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_0),
.Y(n_300)
);


endmodule