module real_jpeg_28698_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_3),
.A2(n_6),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_5),
.A2(n_6),
.B1(n_22),
.B2(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_7),
.B(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_5),
.A2(n_35),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_5),
.B(n_17),
.Y(n_91)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_7),
.B1(n_19),
.B2(n_22),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_26),
.B(n_45),
.C(n_46),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_22),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_83),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_82),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_56),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_13),
.B(n_56),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_29),
.C(n_43),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_15),
.B1(n_29),
.B2(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B(n_24),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_16),
.A2(n_21),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_18),
.A2(n_20),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_18),
.A2(n_26),
.B(n_37),
.C(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_26),
.B(n_33),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_29),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_29),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B(n_38),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_31),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_34),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_43),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_55),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_76),
.B2(n_77),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_81),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_92),
.C(n_94),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_112),
.B(n_116),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_96),
.B(n_111),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_89),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_108),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B(n_110),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_107),
.B(n_109),
.Y(n_101)
);

INVx5_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);


endmodule