module real_jpeg_17681_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_8),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_49),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_1),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_1),
.B(n_116),
.Y(n_115)
);

NAND2x1_ASAP7_75t_SL g136 ( 
.A(n_1),
.B(n_137),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_5),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_6),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_49),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_92),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_6),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_7),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_7),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_7),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_7),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_7),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_9),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_9),
.B(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_10),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

BUFx8_ASAP7_75t_L g175 ( 
.A(n_13),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_13),
.Y(n_214)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_301),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_268),
.B(n_299),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_226),
.B(n_262),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_191),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_153),
.B(n_190),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_125),
.B(n_152),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_97),
.B(n_124),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_60),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_60),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_45),
.C(n_54),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_27),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_27)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_28),
.A2(n_43),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

O2A1O1Ixp5_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_106),
.B(n_115),
.C(n_143),
.Y(n_160)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_34),
.A2(n_35),
.B1(n_131),
.B2(n_138),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_34),
.B(n_138),
.C(n_198),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_34),
.B(n_143),
.C(n_292),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_35),
.B(n_39),
.C(n_43),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_35),
.B(n_291),
.Y(n_290)
);

OR2x4_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_36),
.Y(n_240)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_52),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_38),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_39),
.A2(n_40),
.B1(n_165),
.B2(n_168),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_40),
.B(n_203),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_40),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_40),
.B(n_82),
.C(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_45),
.A2(n_54),
.B1(n_55),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_45),
.A2(n_46),
.B(n_50),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_50),
.A2(n_51),
.B1(n_64),
.B2(n_65),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_50),
.A2(n_51),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_51),
.B(n_213),
.C(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_56),
.A2(n_57),
.B1(n_103),
.B2(n_104),
.Y(n_257)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_65),
.B(n_76),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_57),
.B(n_103),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_57),
.A2(n_103),
.B(n_253),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_57),
.B(n_64),
.C(n_136),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_79),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_80),
.C(n_96),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_112),
.B(n_117),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_63),
.A2(n_71),
.B(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_64),
.A2(n_65),
.B1(n_114),
.B2(n_115),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_100),
.B(n_102),
.C(n_106),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_77),
.B1(n_100),
.B2(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_75),
.A2(n_78),
.B1(n_135),
.B2(n_136),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_76),
.B(n_131),
.C(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_95),
.B2(n_96),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_94),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_87),
.C(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_82),
.A2(n_94),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

AOI22x1_ASAP7_75t_SL g237 ( 
.A1(n_87),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_87),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_87),
.B(n_236),
.C(n_239),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_87),
.B(n_212),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_87),
.A2(n_173),
.B1(n_174),
.B2(n_238),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_90),
.B(n_164),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_93),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_94),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_110),
.B(n_123),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_100),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_100),
.B(n_114),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_100),
.B(n_115),
.C(n_174),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_100),
.A2(n_121),
.B1(n_202),
.B2(n_206),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_100),
.B(n_204),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_103),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_103),
.A2(n_104),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_103),
.B(n_149),
.C(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_119),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_118),
.B(n_122),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_115),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_121),
.B(n_203),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_127),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_140),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_139),
.C(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_138),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_135),
.A2(n_136),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_147),
.C(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g291 ( 
.A1(n_143),
.A2(n_144),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_155),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_169),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_158),
.C(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_163),
.C(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_162),
.B(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_165),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_189),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_177),
.C(n_189),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_188),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_183),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_183),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_183),
.Y(n_310)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_192),
.B(n_193),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_209),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_210),
.C(n_225),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_207),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_200),
.C(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_225),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_221),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_223),
.C(n_224),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_212),
.B(n_238),
.C(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_261),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_261),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_230),
.C(n_245),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_244),
.B2(n_245),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_242),
.B2(n_243),
.Y(n_233)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_272),
.C(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_258),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_251),
.C(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_298),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_298),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_275),
.C(n_286),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_286),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_283),
.B2(n_284),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_284),
.C(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2x1_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_297),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_290),
.C(n_297),
.Y(n_327)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_328),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_305),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_321),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule