module fake_netlist_6_2236_n_787 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_787);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_787;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g158 ( 
.A(n_40),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_42),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_4),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_13),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_78),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_116),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_44),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_39),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_83),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_23),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_18),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_32),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_65),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_37),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_16),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_80),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_74),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_85),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_27),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_51),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_73),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_92),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_47),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_62),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_49),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_87),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_93),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_22),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_26),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_58),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_53),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_67),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_178),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_20),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_0),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_175),
.A2(n_0),
.B(n_1),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_21),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_1),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_166),
.B(n_2),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_167),
.B(n_2),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_159),
.B(n_3),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_174),
.B(n_203),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_170),
.B(n_24),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_R g258 ( 
.A(n_227),
.B(n_160),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_228),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_201),
.B(n_208),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_227),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_219),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_226),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_213),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_161),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_216),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_216),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_166),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_236),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_236),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_163),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_236),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_220),
.B(n_204),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_233),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_215),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_232),
.B(n_180),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_251),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_256),
.B(n_193),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_251),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_241),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_215),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_246),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_232),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_237),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_283),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_250),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_301),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_250),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_275),
.B(n_193),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_293),
.B(n_250),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_287),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_255),
.B(n_254),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_284),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_221),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_256),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_221),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_255),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_231),
.C(n_229),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_221),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_272),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_292),
.B(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_271),
.B(n_244),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_224),
.C(n_251),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_268),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_251),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_273),
.B(n_240),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_265),
.B(n_212),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_240),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_276),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_266),
.B(n_267),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_257),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_251),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_269),
.B(n_240),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_R g354 ( 
.A(n_260),
.B(n_176),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_281),
.B(n_244),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_259),
.B(n_212),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_270),
.B(n_177),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_264),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_264),
.B(n_240),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_264),
.B(n_224),
.C(n_186),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_300),
.B(n_184),
.Y(n_363)
);

NOR3xp33_ASAP7_75t_L g364 ( 
.A(n_297),
.B(n_187),
.C(n_223),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_300),
.B(n_190),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_300),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_299),
.B(n_240),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_285),
.A2(n_225),
.B1(n_218),
.B2(n_247),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_300),
.B(n_192),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_285),
.A2(n_225),
.B1(n_218),
.B2(n_247),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_258),
.Y(n_371)
);

NOR2x1p5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_321),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_307),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_317),
.A2(n_217),
.B(n_222),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_311),
.B(n_247),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_371),
.B(n_194),
.Y(n_378)
);

NOR2x2_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_3),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_342),
.B(n_195),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_311),
.A2(n_308),
.B1(n_328),
.B2(n_342),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_223),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_199),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_341),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_200),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_336),
.Y(n_390)
);

AND3x1_ASAP7_75t_L g391 ( 
.A(n_308),
.B(n_244),
.C(n_222),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_328),
.B(n_202),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_331),
.B(n_247),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

NOR2x1_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_247),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_331),
.B(n_334),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

NOR3xp33_ASAP7_75t_SL g404 ( 
.A(n_320),
.B(n_207),
.C(n_210),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_306),
.B(n_211),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_310),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_320),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_315),
.B(n_217),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_238),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_238),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_324),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_365),
.A2(n_218),
.B1(n_239),
.B2(n_242),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_358),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_239),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_335),
.B(n_242),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_335),
.B(n_234),
.Y(n_418)
);

AND2x4_ASAP7_75t_SL g419 ( 
.A(n_348),
.B(n_234),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_351),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_367),
.A2(n_234),
.B(n_218),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_327),
.B(n_218),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_234),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_314),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_319),
.A2(n_234),
.B1(n_7),
.B2(n_8),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_354),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_322),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_316),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_329),
.B(n_6),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_323),
.B(n_25),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_354),
.B(n_7),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_355),
.B(n_8),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_326),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_353),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_352),
.B(n_28),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_355),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_438)
);

AND3x1_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_12),
.C(n_14),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_363),
.B(n_15),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_369),
.Y(n_441)
);

OA22x2_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_344),
.B1(n_349),
.B2(n_357),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_374),
.A2(n_360),
.B(n_352),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_407),
.A2(n_359),
.B(n_16),
.C(n_17),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_405),
.A2(n_15),
.B1(n_17),
.B2(n_29),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_30),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_426),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_427),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_390),
.B(n_31),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_383),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

AOI22x1_ASAP7_75t_L g457 ( 
.A1(n_372),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_417),
.B(n_43),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_380),
.B(n_45),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_46),
.B(n_48),
.C(n_50),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_392),
.A2(n_52),
.B(n_54),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_391),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_SL g464 ( 
.A(n_433),
.B(n_59),
.C(n_60),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_392),
.A2(n_63),
.B(n_64),
.Y(n_465)
);

O2A1O1Ixp5_ASAP7_75t_L g466 ( 
.A1(n_374),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_408),
.B(n_71),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_408),
.B(n_72),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

O2A1O1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_430),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_392),
.A2(n_79),
.B(n_81),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_418),
.B(n_394),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_394),
.B(n_84),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_377),
.B(n_86),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_88),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_439),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_419),
.B(n_96),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

OAI22x1_ASAP7_75t_L g482 ( 
.A1(n_387),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_392),
.A2(n_101),
.B(n_102),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_440),
.A2(n_432),
.B(n_436),
.C(n_411),
.Y(n_484)
);

O2A1O1Ixp33_ASAP7_75t_L g485 ( 
.A1(n_411),
.A2(n_103),
.B(n_104),
.C(n_105),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_378),
.B(n_106),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_L g487 ( 
.A1(n_412),
.A2(n_107),
.B(n_108),
.C(n_109),
.Y(n_487)
);

NAND3xp33_ASAP7_75t_SL g488 ( 
.A(n_385),
.B(n_110),
.C(n_111),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

O2A1O1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_412),
.A2(n_416),
.B(n_393),
.C(n_423),
.Y(n_490)
);

O2A1O1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_431),
.A2(n_112),
.B(n_113),
.C(n_114),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_381),
.B(n_117),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_416),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_398),
.A2(n_375),
.B(n_402),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_409),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_405),
.A2(n_123),
.B(n_124),
.C(n_125),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_375),
.A2(n_404),
.B(n_423),
.C(n_403),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_446),
.B(n_413),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_444),
.B(n_389),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_494),
.A2(n_431),
.B(n_421),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_490),
.A2(n_422),
.B(n_437),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_479),
.B(n_386),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_389),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_453),
.B(n_386),
.Y(n_505)
);

NAND2x1p5_ASAP7_75t_L g506 ( 
.A(n_446),
.B(n_415),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_456),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_498),
.A2(n_437),
.B(n_414),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_459),
.B(n_434),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_467),
.B(n_429),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

CKINVDCx11_ASAP7_75t_R g518 ( 
.A(n_446),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_449),
.B(n_428),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_474),
.A2(n_399),
.B(n_382),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_441),
.B(n_398),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_489),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_470),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_475),
.B(n_438),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_476),
.B(n_425),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g532 ( 
.A(n_455),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_455),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_473),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_442),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_SL g536 ( 
.A(n_462),
.B(n_415),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_478),
.B(n_379),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_482),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_468),
.A2(n_415),
.B(n_127),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_484),
.B(n_157),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_478),
.Y(n_541)
);

INVx3_ASAP7_75t_SL g542 ( 
.A(n_458),
.Y(n_542)
);

BUFx8_ASAP7_75t_L g543 ( 
.A(n_448),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_492),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_486),
.B(n_126),
.Y(n_545)
);

BUFx8_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_522),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_539),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_507),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_518),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_508),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_508),
.Y(n_553)
);

CKINVDCx11_ASAP7_75t_R g554 ( 
.A(n_515),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_541),
.A2(n_454),
.B1(n_493),
.B2(n_469),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_512),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_512),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_531),
.A2(n_463),
.B1(n_464),
.B2(n_496),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_524),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_525),
.A2(n_463),
.B1(n_443),
.B2(n_457),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_524),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_517),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g565 ( 
.A1(n_540),
.A2(n_443),
.B(n_465),
.Y(n_565)
);

NAND2x1p5_ASAP7_75t_L g566 ( 
.A(n_536),
.B(n_472),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_500),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_534),
.B(n_466),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_543),
.A2(n_483),
.B1(n_471),
.B2(n_460),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_543),
.A2(n_487),
.B1(n_485),
.B2(n_491),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_500),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

CKINVDCx6p67_ASAP7_75t_R g573 ( 
.A(n_532),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_529),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_546),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_529),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_503),
.B(n_132),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_546),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_535),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_527),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_522),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_528),
.Y(n_586)
);

BUFx8_ASAP7_75t_L g587 ( 
.A(n_514),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_519),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_571),
.B(n_588),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_550),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_SL g591 ( 
.A(n_558),
.B(n_530),
.C(n_538),
.Y(n_591)
);

NOR3xp33_ASAP7_75t_SL g592 ( 
.A(n_562),
.B(n_545),
.C(n_533),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_554),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_588),
.B(n_505),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_559),
.B(n_562),
.Y(n_595)
);

BUFx4f_ASAP7_75t_SL g596 ( 
.A(n_573),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_574),
.Y(n_597)
);

AND2x4_ASAP7_75t_SL g598 ( 
.A(n_573),
.B(n_505),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_556),
.B(n_557),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_571),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_587),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

AOI221xp5_ASAP7_75t_L g603 ( 
.A1(n_558),
.A2(n_511),
.B1(n_504),
.B2(n_544),
.C(n_523),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_537),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_557),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_551),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_567),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_587),
.Y(n_608)
);

NOR2x1_ASAP7_75t_SL g609 ( 
.A(n_550),
.B(n_521),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_580),
.A2(n_537),
.B1(n_542),
.B2(n_547),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

AO31x2_ASAP7_75t_L g612 ( 
.A1(n_561),
.A2(n_502),
.A3(n_533),
.B(n_501),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_548),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_570),
.B(n_513),
.C(n_519),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_564),
.B(n_516),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_R g616 ( 
.A(n_578),
.B(n_547),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_564),
.B(n_516),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_588),
.A2(n_513),
.B1(n_520),
.B2(n_148),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_568),
.B(n_144),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_548),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_552),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_578),
.B(n_146),
.Y(n_623)
);

NAND2x1p5_ASAP7_75t_L g624 ( 
.A(n_574),
.B(n_149),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_553),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_575),
.B(n_154),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_553),
.B(n_155),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_575),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_582),
.A2(n_569),
.B1(n_577),
.B2(n_581),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_560),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_585),
.B(n_586),
.Y(n_631)
);

AND2x2_ASAP7_75t_SL g632 ( 
.A(n_568),
.B(n_579),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_579),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_585),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_560),
.B(n_572),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_SL g636 ( 
.A(n_584),
.B(n_555),
.C(n_566),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_605),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_572),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_636),
.B(n_576),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_635),
.B(n_576),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_589),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_600),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_600),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_612),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_591),
.B(n_584),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_605),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

AND2x4_ASAP7_75t_SL g648 ( 
.A(n_636),
.B(n_549),
.Y(n_648)
);

NOR4xp25_ASAP7_75t_SL g649 ( 
.A(n_620),
.B(n_555),
.C(n_566),
.D(n_549),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_602),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_563),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_628),
.Y(n_652)
);

AND2x2_ASAP7_75t_SL g653 ( 
.A(n_629),
.B(n_549),
.Y(n_653)
);

AO21x2_ASAP7_75t_L g654 ( 
.A1(n_609),
.A2(n_565),
.B(n_592),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_595),
.Y(n_655)
);

NOR4xp25_ASAP7_75t_SL g656 ( 
.A(n_603),
.B(n_566),
.C(n_565),
.D(n_586),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_622),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_633),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_612),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_591),
.B(n_583),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_599),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_589),
.B(n_583),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_599),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_630),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_589),
.Y(n_665)
);

AO21x2_ASAP7_75t_L g666 ( 
.A1(n_618),
.A2(n_586),
.B(n_614),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_603),
.A2(n_610),
.B1(n_604),
.B2(n_594),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_627),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_627),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_653),
.A2(n_594),
.B1(n_625),
.B2(n_608),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_652),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_641),
.B(n_619),
.Y(n_672)
);

AOI221xp5_ASAP7_75t_L g673 ( 
.A1(n_667),
.A2(n_625),
.B1(n_617),
.B2(n_615),
.C(n_621),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_641),
.B(n_619),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_652),
.B(n_626),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_653),
.A2(n_607),
.B1(n_606),
.B2(n_601),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_647),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_647),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_658),
.B(n_613),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_658),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_657),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_638),
.B(n_624),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_638),
.B(n_624),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_655),
.B(n_634),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_650),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_642),
.B(n_631),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_665),
.B(n_662),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_646),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_640),
.B(n_597),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_650),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_640),
.B(n_597),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_643),
.B(n_593),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_668),
.B(n_616),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_668),
.B(n_598),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_645),
.B(n_659),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_651),
.B(n_611),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_651),
.B(n_623),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_685),
.B(n_660),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_690),
.B(n_646),
.Y(n_699)
);

INVx6_ASAP7_75t_L g700 ( 
.A(n_672),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_677),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_678),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_680),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_688),
.B(n_639),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_687),
.B(n_665),
.Y(n_705)
);

INVxp33_ASAP7_75t_SL g706 ( 
.A(n_692),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_671),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_681),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_687),
.B(n_662),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_687),
.B(n_662),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_688),
.B(n_660),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_698),
.B(n_695),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

OAI211xp5_ASAP7_75t_SL g714 ( 
.A1(n_699),
.A2(n_693),
.B(n_676),
.C(n_686),
.Y(n_714)
);

O2A1O1Ixp5_ASAP7_75t_R g715 ( 
.A1(n_699),
.A2(n_684),
.B(n_694),
.C(n_649),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_711),
.B(n_679),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_701),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_706),
.B(n_697),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_702),
.Y(n_719)
);

OA222x2_ASAP7_75t_L g720 ( 
.A1(n_703),
.A2(n_695),
.B1(n_645),
.B2(n_644),
.C1(n_669),
.C2(n_671),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_715),
.A2(n_670),
.B1(n_704),
.B2(n_648),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_714),
.A2(n_697),
.B(n_679),
.C(n_696),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_718),
.A2(n_704),
.B(n_696),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_716),
.B(n_708),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_717),
.A2(n_653),
.B(n_682),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_722),
.B(n_719),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_721),
.B(n_596),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_724),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_673),
.C(n_712),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_723),
.B(n_712),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_724),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_731),
.B(n_713),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_730),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_727),
.Y(n_734)
);

NOR3x1_ASAP7_75t_L g735 ( 
.A(n_733),
.B(n_729),
.C(n_728),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_734),
.B(n_710),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_736),
.A2(n_732),
.B(n_648),
.Y(n_737)
);

NAND4xp25_ASAP7_75t_L g738 ( 
.A(n_735),
.B(n_682),
.C(n_683),
.D(n_691),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_735),
.A2(n_720),
.B(n_666),
.C(n_669),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_738),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_739),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_737),
.B(n_654),
.Y(n_742)
);

NOR2x1_ASAP7_75t_L g743 ( 
.A(n_738),
.B(n_654),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_738),
.B(n_689),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_738),
.Y(n_745)
);

NAND3x1_ASAP7_75t_L g746 ( 
.A(n_741),
.B(n_683),
.C(n_709),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_745),
.B(n_705),
.Y(n_747)
);

INVxp33_ASAP7_75t_SL g748 ( 
.A(n_740),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_744),
.B(n_705),
.Y(n_749)
);

NAND4xp75_ASAP7_75t_L g750 ( 
.A(n_743),
.B(n_691),
.C(n_689),
.D(n_675),
.Y(n_750)
);

NOR4xp75_ASAP7_75t_SL g751 ( 
.A(n_742),
.B(n_700),
.C(n_648),
.D(n_656),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_740),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_747),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_748),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_752),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_749),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_746),
.Y(n_757)
);

XNOR2xp5_ASAP7_75t_L g758 ( 
.A(n_750),
.B(n_751),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_748),
.Y(n_759)
);

XNOR2x2_ASAP7_75t_L g760 ( 
.A(n_754),
.B(n_675),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_753),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_756),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_758),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_759),
.A2(n_700),
.B1(n_672),
.B2(n_674),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_757),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_755),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_755),
.Y(n_768)
);

OAI31xp33_ASAP7_75t_L g769 ( 
.A1(n_766),
.A2(n_768),
.A3(n_761),
.B(n_767),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_762),
.B(n_700),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_764),
.A2(n_674),
.B1(n_672),
.B2(n_639),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_765),
.A2(n_674),
.B1(n_639),
.B2(n_669),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_763),
.A2(n_639),
.B1(n_666),
.B2(n_662),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_760),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_762),
.Y(n_775)
);

OAI31xp33_ASAP7_75t_L g776 ( 
.A1(n_766),
.A2(n_664),
.A3(n_663),
.B(n_661),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_775),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_769),
.A2(n_664),
.B(n_654),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_SL g779 ( 
.A1(n_774),
.A2(n_637),
.B1(n_657),
.B2(n_663),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_770),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_772),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_780),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_777),
.Y(n_783)
);

AO22x2_ASAP7_75t_L g784 ( 
.A1(n_783),
.A2(n_781),
.B1(n_778),
.B2(n_779),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_784),
.A2(n_782),
.B1(n_771),
.B2(n_773),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_785),
.B(n_776),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_786),
.A2(n_666),
.B1(n_644),
.B2(n_681),
.Y(n_787)
);


endmodule