module real_jpeg_32924_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_715, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_715;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_620;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_605;
wire n_216;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_634;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_704;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_195;
wire n_110;
wire n_703;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_712;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_711;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_667;
wire n_375;
wire n_708;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_713;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_0),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_0),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_1),
.A2(n_217),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_1),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_1),
.A2(n_288),
.B1(n_365),
.B2(n_368),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_1),
.A2(n_288),
.B1(n_543),
.B2(n_546),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_1),
.A2(n_288),
.B1(n_607),
.B2(n_608),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22x1_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_213),
.B1(n_214),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_3),
.Y(n_213)
);

AOI22x1_ASAP7_75t_SL g295 ( 
.A1(n_3),
.A2(n_213),
.B1(n_296),
.B2(n_300),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_3),
.A2(n_213),
.B1(n_353),
.B2(n_357),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_3),
.A2(n_213),
.B1(n_407),
.B2(n_412),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_4),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_128),
.B1(n_131),
.B2(n_133),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_5),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_133),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_5),
.A2(n_133),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_5),
.A2(n_133),
.B1(n_444),
.B2(n_448),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_6),
.A2(n_123),
.B1(n_215),
.B2(n_387),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_6),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_6),
.A2(n_387),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_6),
.A2(n_387),
.B1(n_582),
.B2(n_584),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_6),
.A2(n_387),
.B1(n_589),
.B2(n_630),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_66),
.B1(n_70),
.B2(n_75),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_75),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_7),
.A2(n_75),
.B1(n_167),
.B2(n_170),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_7),
.A2(n_75),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_8),
.A2(n_378),
.B(n_382),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_8),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_8),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g549 ( 
.A1(n_8),
.A2(n_422),
.A3(n_550),
.B1(n_553),
.B2(n_554),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_8),
.B(n_165),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_8),
.A2(n_195),
.B1(n_629),
.B2(n_645),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_8),
.A2(n_418),
.B1(n_670),
.B2(n_674),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_63),
.B1(n_156),
.B2(n_160),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_9),
.A2(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_238),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_9),
.A2(n_63),
.B1(n_206),
.B2(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_11),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_12),
.Y(n_447)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_13),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_14),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_14),
.Y(n_124)
);

OAI22x1_ASAP7_75t_SL g249 ( 
.A1(n_14),
.A2(n_124),
.B1(n_250),
.B2(n_256),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_14),
.A2(n_124),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_14),
.A2(n_124),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_15),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_15),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_15),
.A2(n_225),
.B1(n_347),
.B2(n_350),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_15),
.A2(n_225),
.B1(n_468),
.B2(n_470),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_15),
.A2(n_225),
.B1(n_468),
.B2(n_470),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_15),
.A2(n_225),
.B1(n_558),
.B2(n_560),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_16),
.A2(n_368),
.B1(n_371),
.B2(n_374),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_16),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_16),
.A2(n_67),
.B1(n_374),
.B2(n_477),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_16),
.A2(n_374),
.B1(n_617),
.B2(n_620),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_16),
.A2(n_374),
.B1(n_634),
.B2(n_637),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_17),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_18),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_18),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_19),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_19),
.Y(n_169)
);

OAI31xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_180),
.A3(n_704),
.B(n_710),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_22),
.B(n_704),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_179),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_77),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_25),
.B(n_77),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND4xp25_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_52),
.C(n_64),
.D(n_76),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_R g27 ( 
.A(n_28),
.B(n_51),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_28),
.A2(n_51),
.B1(n_121),
.B2(n_127),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_28),
.A2(n_51),
.B1(n_53),
.B2(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_29),
.A2(n_122),
.B1(n_211),
.B2(n_212),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_29),
.A2(n_211),
.B1(n_475),
.B2(n_480),
.Y(n_474)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_30),
.A2(n_51),
.B1(n_377),
.B2(n_386),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_30),
.A2(n_51),
.B1(n_287),
.B2(n_476),
.Y(n_494)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_31),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_31),
.A2(n_211),
.B1(n_221),
.B2(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_42),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_35),
.Y(n_291)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_36),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_36),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_37),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_38),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_39),
.Y(n_132)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_45),
.Y(n_163)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_45),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_46),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_46),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_47),
.Y(n_159)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_47),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_47),
.Y(n_436)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_51),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_51),
.B(n_418),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_62),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g226 ( 
.A(n_68),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_73),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_74),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_175),
.C(n_176),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_78),
.A2(n_79),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_120),
.C(n_134),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_80),
.A2(n_312),
.B1(n_313),
.B2(n_315),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_80),
.A2(n_135),
.B1(n_315),
.B2(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_109),
.B(n_112),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_81),
.B(n_268),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_81),
.A2(n_109),
.B(n_112),
.Y(n_315)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_82),
.A2(n_110),
.B1(n_229),
.B2(n_234),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_82),
.Y(n_246)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_82),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_82),
.A2(n_269),
.B1(n_352),
.B2(n_361),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_82),
.A2(n_361),
.B1(n_616),
.B2(n_622),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_91),
.B(n_99),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_89),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_90),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_90),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_90),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_91),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_96),
.Y(n_359)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_97),
.Y(n_231)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_97),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_98),
.Y(n_274)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_107),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_101),
.Y(n_404)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_101),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_101),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_101),
.Y(n_651)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_106),
.Y(n_415)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_109),
.A2(n_112),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_109),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_109),
.B(n_276),
.Y(n_501)
);

AO22x1_ASAP7_75t_L g541 ( 
.A1(n_109),
.A2(n_345),
.B1(n_346),
.B2(n_542),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_109),
.A2(n_246),
.B1(n_542),
.B2(n_667),
.Y(n_666)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_110),
.B(n_418),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_111),
.Y(n_362)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_118),
.Y(n_233)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_119),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_119),
.Y(n_580)
);

XOR2x2_ASAP7_75t_L g325 ( 
.A(n_120),
.B(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_135),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_155),
.B1(n_164),
.B2(n_166),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_136),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_136),
.A2(n_155),
.B1(n_164),
.B2(n_314),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g363 ( 
.A1(n_136),
.A2(n_164),
.B1(n_364),
.B2(n_370),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_136),
.A2(n_164),
.B1(n_370),
.B2(n_391),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_136),
.A2(n_164),
.B1(n_364),
.B2(n_467),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_136),
.A2(n_164),
.B1(n_295),
.B2(n_496),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_136),
.A2(n_164),
.B1(n_391),
.B2(n_669),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_142),
.B(n_148),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_142),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_143),
.Y(n_300)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_144),
.Y(n_396)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_144),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_149),
.Y(n_585)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_159),
.Y(n_675)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_165),
.A2(n_177),
.B1(n_249),
.B2(n_260),
.Y(n_248)
);

AOI22x1_ASAP7_75t_L g293 ( 
.A1(n_165),
.A2(n_177),
.B1(n_249),
.B2(n_294),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

INVx8_ASAP7_75t_L g367 ( 
.A(n_169),
.Y(n_367)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_174),
.Y(n_673)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_175),
.B(n_176),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_180),
.A2(n_711),
.B(n_712),
.Y(n_710)
);

OAI21x1_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_330),
.B(n_697),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_316),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_301),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_184),
.B(n_301),
.Y(n_700)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_243),
.C(n_265),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_186),
.A2(n_243),
.B1(n_244),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_186),
.Y(n_524)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_227),
.B2(n_242),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_210),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_189),
.A2(n_303),
.B1(n_305),
.B2(n_715),
.Y(n_302)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_189),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_194),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_195),
.A2(n_202),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_195),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_195),
.A2(n_282),
.B1(n_440),
.B2(n_443),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_195),
.A2(n_603),
.B1(n_605),
.B2(n_606),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_195),
.A2(n_629),
.B1(n_633),
.B2(n_640),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

BUFx2_ASAP7_75t_R g405 ( 
.A(n_196),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_196),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_197),
.Y(n_641)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_197),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_206),
.Y(n_607)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_209),
.Y(n_411)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_209),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_210),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B(n_220),
.Y(n_210)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_224),
.Y(n_428)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_228),
.Y(n_514)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_230),
.Y(n_546)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_240),
.Y(n_583)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_248),
.B(n_264),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_248),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_246),
.A2(n_360),
.B1(n_573),
.B2(n_581),
.Y(n_572)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_259),
.Y(n_369)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_265),
.B(n_523),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_284),
.C(n_292),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_266),
.B(n_518),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_275),
.B(n_277),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_267),
.B(n_501),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx4f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_274),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_277),
.B(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_279),
.B(n_418),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx8_ASAP7_75t_L g604 ( 
.A(n_281),
.Y(n_604)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_283),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_285),
.B(n_293),
.Y(n_518)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_308),
.C(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_320),
.C(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_317),
.B(n_700),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_328),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_SL g702 ( 
.A(n_318),
.B(n_328),
.Y(n_702)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_320),
.C(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_337),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g697 ( 
.A1(n_331),
.A2(n_698),
.B(n_703),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_336),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_332),
.B(n_336),
.Y(n_703)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AO21x2_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_525),
.B(n_690),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_504),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_484),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_458),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_341),
.B(n_458),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_388),
.C(n_419),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_342),
.B(n_529),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_375),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_363),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_344),
.B(n_363),
.C(n_375),
.Y(n_463)
);

AOI22x1_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_351),
.B2(n_360),
.Y(n_344)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_357),
.B(n_418),
.Y(n_554)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_382),
.Y(n_437)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_389),
.B(n_419),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_397),
.C(n_417),
.Y(n_389)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_390),
.Y(n_533)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_397),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_397),
.A2(n_534),
.B(n_535),
.Y(n_539)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_398),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_405),
.B1(n_406),
.B2(n_416),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_399),
.A2(n_416),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_406),
.A2(n_416),
.B1(n_557),
.B2(n_564),
.Y(n_556)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_411),
.Y(n_559)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_411),
.Y(n_599)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_411),
.Y(n_632)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_415),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_416),
.A2(n_655),
.B1(n_656),
.B2(n_657),
.Y(n_654)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_417),
.B(n_538),
.Y(n_537)
);

OAI21xp33_ASAP7_75t_SL g573 ( 
.A1(n_418),
.A2(n_574),
.B(n_577),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_418),
.B(n_578),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_438),
.B1(n_452),
.B2(n_457),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_420),
.B(n_457),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_424),
.A3(n_427),
.B1(n_429),
.B2(n_437),
.Y(n_420)
);

OAI32xp33_ASAP7_75t_L g453 ( 
.A1(n_421),
.A2(n_424),
.A3(n_429),
.B1(n_437),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_447),
.Y(n_612)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_464),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_460),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_461),
.B(n_462),
.Y(n_491)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

MAJx2_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_486),
.C(n_487),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_483),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_474),
.B1(n_481),
.B2(n_482),
.Y(n_465)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_466),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_481),
.C(n_483),
.Y(n_503)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx8_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NAND2xp67_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_488),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g692 ( 
.A(n_485),
.B(n_488),
.C(n_693),
.Y(n_692)
);

XOR2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_503),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_498),
.B1(n_499),
.B2(n_502),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_490),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_493),
.C(n_510),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_494),
.B1(n_495),
.B2(n_497),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_495),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_497),
.Y(n_510)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_503),
.C(n_507),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g690 ( 
.A1(n_504),
.A2(n_691),
.B(n_694),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_519),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_506),
.B(n_508),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_511),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_512),
.C(n_521),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_517),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_515),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_517),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_519),
.A2(n_695),
.B(n_696),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_522),
.Y(n_696)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_566),
.B(n_689),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_528),
.B(n_530),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_SL g689 ( 
.A(n_528),
.B(n_530),
.Y(n_689)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_541),
.C(n_547),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_531),
.B(n_684),
.Y(n_683)
);

AOI22x1_ASAP7_75t_L g531 ( 
.A1(n_532),
.A2(n_537),
.B1(n_539),
.B2(n_540),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_536),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_541),
.A2(n_685),
.B(n_686),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_541),
.B(n_548),
.Y(n_686)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_547),
.Y(n_685)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_555),
.Y(n_548)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_549),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_549),
.B(n_556),
.Y(n_680)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_555),
.Y(n_679)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_557),
.Y(n_605)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_567),
.A2(n_682),
.B(n_688),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g567 ( 
.A1(n_568),
.A2(n_661),
.B(n_681),
.Y(n_567)
);

OAI21x1_ASAP7_75t_SL g568 ( 
.A1(n_569),
.A2(n_625),
.B(n_660),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_601),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_570),
.B(n_601),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_571),
.B(n_586),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_571),
.A2(n_572),
.B1(n_586),
.B2(n_587),
.Y(n_658)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_577),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_581),
.Y(n_622)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_588),
.A2(n_595),
.B1(n_596),
.B2(n_600),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_SL g588 ( 
.A(n_589),
.B(n_591),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_602),
.B(n_613),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_602),
.B(n_615),
.C(n_623),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_606),
.Y(n_656)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_614),
.A2(n_615),
.B1(n_623),
.B2(n_624),
.Y(n_613)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_614),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_615),
.Y(n_624)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_616),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

AOI21x1_ASAP7_75t_SL g625 ( 
.A1(n_626),
.A2(n_653),
.B(n_659),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_627),
.A2(n_643),
.B(n_652),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_628),
.B(n_642),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_628),
.B(n_642),
.Y(n_652)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_633),
.Y(n_655)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_644),
.B(n_646),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_647),
.B(n_648),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

BUFx2_ASAP7_75t_SL g650 ( 
.A(n_651),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_654),
.B(n_658),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g659 ( 
.A(n_654),
.B(n_658),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_663),
.Y(n_661)
);

NOR2x1_ASAP7_75t_L g681 ( 
.A(n_662),
.B(n_663),
.Y(n_681)
);

XNOR2x1_ASAP7_75t_L g663 ( 
.A(n_664),
.B(n_677),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_665),
.A2(n_666),
.B1(n_668),
.B2(n_676),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_666),
.B(n_676),
.C(n_677),
.Y(n_687)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_668),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_671),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_673),
.Y(n_672)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_675),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g677 ( 
.A1(n_678),
.A2(n_679),
.B(n_680),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_SL g682 ( 
.A(n_683),
.B(n_687),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_683),
.B(n_687),
.Y(n_688)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_692),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g698 ( 
.A(n_699),
.B(n_701),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g701 ( 
.A(n_702),
.Y(n_701)
);

NOR2x1_ASAP7_75t_R g712 ( 
.A(n_704),
.B(n_713),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_705),
.B(n_709),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_706),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_707),
.Y(n_706)
);

BUFx12f_ASAP7_75t_SL g707 ( 
.A(n_708),
.Y(n_707)
);

INVx6_ASAP7_75t_L g713 ( 
.A(n_708),
.Y(n_713)
);


endmodule