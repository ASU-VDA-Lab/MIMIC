module fake_aes_111_n_23 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_23;
wire n_20;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_5), .Y(n_8) );
NOR2xp67_ASAP7_75t_L g9 ( .A(n_3), .B(n_7), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_13), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_10), .B1(n_9), .B2(n_8), .Y(n_17) );
O2A1O1Ixp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_15), .B(n_14), .C(n_9), .Y(n_18) );
OAI221xp5_ASAP7_75t_SL g19 ( .A1(n_17), .A2(n_15), .B1(n_14), .B2(n_2), .C(n_3), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
BUFx8_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_20), .B(n_0), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_21), .B1(n_1), .B2(n_6), .Y(n_23) );
endmodule