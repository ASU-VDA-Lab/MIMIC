module real_jpeg_5868_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_2),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_3),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_3),
.B(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_5),
.B(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_8),
.B(n_37),
.Y(n_114)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_11),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_102),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_67),
.B(n_101),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_49),
.B(n_66),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_39),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_39),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_25),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_22),
.C(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_20),
.Y(n_120)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_33),
.B(n_38),
.Y(n_90)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_60),
.B(n_65),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_64),
.Y(n_65)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_69),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_88),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_89),
.C(n_92),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_82),
.C(n_87),
.Y(n_116)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_83),
.B2(n_87),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_133),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_132),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_132),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);


endmodule