module fake_jpeg_6010_n_80 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_42),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_45),
.B1(n_47),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_41),
.B1(n_58),
.B2(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_72),
.B(n_2),
.C(n_9),
.D(n_10),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_44),
.B1(n_3),
.B2(n_8),
.Y(n_72)
);

AO221x1_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.C(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_20),
.Y(n_77)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_24),
.A3(n_25),
.B1(n_26),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_78)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_30),
.B(n_31),
.C(n_33),
.D(n_34),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_35),
.Y(n_80)
);


endmodule