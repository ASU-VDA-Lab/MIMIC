module fake_jpeg_8915_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_51),
.Y(n_78)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_36),
.B(n_38),
.C(n_31),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_28),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_18),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_0),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_0),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_27),
.A3(n_21),
.B1(n_30),
.B2(n_17),
.Y(n_107)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_66),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_45),
.B1(n_49),
.B2(n_43),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_79),
.A3(n_88),
.B1(n_30),
.B2(n_21),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_77),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_19),
.B1(n_34),
.B2(n_20),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_19),
.B1(n_34),
.B2(n_20),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_19),
.B1(n_34),
.B2(n_20),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_75),
.B1(n_26),
.B2(n_28),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_27),
.B1(n_38),
.B2(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_18),
.B1(n_21),
.B2(n_30),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_39),
.B1(n_23),
.B2(n_37),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_39),
.C(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_51),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_30),
.B1(n_18),
.B2(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_94),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_88),
.B1(n_65),
.B2(n_59),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_104),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_110),
.B1(n_67),
.B2(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_88),
.B1(n_62),
.B2(n_80),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_47),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_29),
.C(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_86),
.Y(n_104)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_67),
.B1(n_79),
.B2(n_71),
.Y(n_131)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_119),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_40),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_61),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_22),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_40),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_134),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_130),
.B(n_136),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_154),
.B1(n_92),
.B2(n_89),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_68),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_148),
.B(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_135),
.B(n_146),
.Y(n_196)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_59),
.A3(n_68),
.B1(n_79),
.B2(n_88),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_147),
.B1(n_112),
.B2(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_85),
.B1(n_22),
.B2(n_17),
.Y(n_147)
);

AO21x2_ASAP7_75t_SL g148 ( 
.A1(n_98),
.A2(n_50),
.B(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_153),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_17),
.B(n_22),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_155),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_50),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

AO21x2_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_50),
.B(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_1),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_40),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_100),
.B1(n_89),
.B2(n_121),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_9),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_1),
.C(n_2),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_177),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_93),
.B1(n_97),
.B2(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_179),
.B1(n_185),
.B2(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_170),
.B(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_126),
.B(n_13),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_120),
.B1(n_105),
.B2(n_111),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_123),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_189),
.B1(n_192),
.B2(n_175),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_188),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_154),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_3),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_145),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_12),
.B1(n_15),
.B2(n_6),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_135),
.B1(n_160),
.B2(n_134),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_7),
.B1(n_9),
.B2(n_13),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_149),
.B(n_153),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_7),
.B1(n_14),
.B2(n_16),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_183),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_200),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_201),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_140),
.C(n_150),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_209),
.Y(n_235)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_130),
.B(n_136),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_211),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_159),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_138),
.B1(n_158),
.B2(n_129),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

XOR2x2_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_226),
.B1(n_227),
.B2(n_181),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_128),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_166),
.A2(n_151),
.B1(n_126),
.B2(n_137),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_174),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_16),
.B(n_5),
.C(n_4),
.D(n_158),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_162),
.A2(n_132),
.B(n_129),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_162),
.C(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_163),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_196),
.A2(n_179),
.B1(n_164),
.B2(n_167),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_196),
.A2(n_192),
.B1(n_188),
.B2(n_191),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_199),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_198),
.B1(n_227),
.B2(n_211),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_189),
.B1(n_182),
.B2(n_170),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_244),
.C(n_225),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_176),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_228),
.B(n_246),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_218),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_174),
.B1(n_194),
.B2(n_221),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_201),
.B1(n_215),
.B2(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_255),
.B(n_270),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_232),
.B(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_261),
.C(n_265),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_205),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_209),
.C(n_204),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_270),
.B(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_213),
.C(n_219),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_212),
.A3(n_220),
.B1(n_208),
.B2(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_202),
.B1(n_222),
.B2(n_208),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_249),
.B(n_236),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_SL g271 ( 
.A(n_231),
.B(n_252),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_233),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g273 ( 
.A(n_239),
.B(n_248),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_229),
.B1(n_243),
.B2(n_260),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_250),
.B1(n_239),
.B2(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_282),
.B1(n_283),
.B2(n_265),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_250),
.B1(n_237),
.B2(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_229),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_258),
.B(n_253),
.C(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_279),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_290),
.Y(n_298)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_268),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.C(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_261),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_258),
.B(n_257),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_259),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_281),
.C(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_280),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_275),
.C(n_293),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_303),
.C(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_302),
.C(n_282),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_286),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_279),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_298),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_316),
.B1(n_305),
.B2(n_296),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_292),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_288),
.B1(n_284),
.B2(n_280),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_294),
.B(n_296),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_304),
.B(n_314),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_312),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_304),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_309),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_328),
.C(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_276),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_328),
.B(n_321),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_325),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_332),
.C(n_324),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_307),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_306),
.C(n_318),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);


endmodule