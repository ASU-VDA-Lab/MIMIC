module real_jpeg_6223_n_30 (n_17, n_8, n_0, n_21, n_168, n_2, n_29, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_28, n_171, n_169, n_167, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_164, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_29;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_28;
input n_171;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_1),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_56),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_2),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_50),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_5),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_6),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_7),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_8),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_8),
.B(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_9),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_143),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_10),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_10),
.B(n_147),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_33),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_13),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_105),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_14),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_15),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_16),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_17),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_18),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_18),
.B(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_20),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_21),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_22),
.B(n_44),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_28),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_28),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_153),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_152),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_38),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_141),
.B(n_149),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_120),
.B(n_135),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_63),
.B(n_108),
.C(n_117),
.Y(n_41)
);

NOR4xp25_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.C(n_55),
.D(n_58),
.Y(n_42)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_54),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_104),
.B(n_107),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_97),
.B(n_103),
.Y(n_64)
);

AO221x1_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_74),
.B1(n_94),
.B2(n_95),
.C(n_96),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_91),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B(n_93),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_78),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_92),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_88),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_102),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_130),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B(n_114),
.C(n_115),
.D(n_116),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.C(n_131),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_131),
.B(n_136),
.C(n_139),
.D(n_140),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_123),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_161),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_164),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_165),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_166),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_167),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_168),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_169),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_170),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_171),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_172),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_173),
.Y(n_106)
);


endmodule