module real_jpeg_24022_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_288;
wire n_300;
wire n_166;
wire n_221;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_285;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_244;
wire n_167;
wire n_128;
wire n_179;
wire n_295;
wire n_133;
wire n_202;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_40),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_2),
.A2(n_40),
.B1(n_62),
.B2(n_64),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_40),
.B1(n_82),
.B2(n_83),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_302),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_303),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_20),
.B1(n_29),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_20),
.B1(n_62),
.B2(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_20),
.B1(n_82),
.B2(n_83),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_69),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_7),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_7),
.A2(n_69),
.B1(n_82),
.B2(n_83),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_22),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_52),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_52),
.B1(n_82),
.B2(n_83),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_9),
.B(n_28),
.C(n_31),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_9),
.B(n_27),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_59),
.C(n_62),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_79),
.C(n_82),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_9),
.B(n_217),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_9),
.B(n_110),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_9),
.B(n_72),
.Y(n_259)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_22),
.B1(n_28),
.B2(n_32),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_43),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_41),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_19),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_21),
.B(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_26),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_27),
.A2(n_33),
.B1(n_50),
.B2(n_67),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_29),
.A2(n_31),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_31),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_36),
.B(n_45),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_48),
.B(n_49),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_85),
.B(n_301),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_46),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_46),
.B(n_299),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_53),
.CI(n_65),
.CON(n_46),
.SN(n_46)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_48),
.A2(n_49),
.B(n_68),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_57),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_56),
.A2(n_61),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_72),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_57),
.B(n_115),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_61),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_61),
.A2(n_114),
.B(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_64),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_62),
.B(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.C(n_73),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_66),
.B(n_133),
.C(n_141),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_66),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_66),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_66),
.A2(n_141),
.B1(n_142),
.B2(n_155),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_66),
.A2(n_112),
.B1(n_155),
.B2(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_66),
.B(n_112),
.C(n_193),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_70),
.A2(n_73),
.B1(n_122),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_70),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_71),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_122),
.B1(n_123),
.B2(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_118),
.C(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_101),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_77),
.A2(n_101),
.B1(n_110),
.B2(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_81),
.A2(n_100),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_82),
.B(n_249),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_298),
.B(n_300),
.Y(n_85)
);

OAI211xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_143),
.B(n_157),
.C(n_297),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_127),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_127),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_105),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_107),
.C(n_116),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_97),
.B(n_102),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_90),
.A2(n_102),
.B1(n_103),
.B2(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_90),
.A2(n_98),
.B1(n_130),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_92),
.B(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_96),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_93),
.B(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_95),
.A2(n_135),
.B(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_95),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_98),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_116),
.B2(n_117),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_108),
.B(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_112),
.B(n_215),
.C(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_112),
.A2(n_205),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_119),
.B1(n_151),
.B2(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_118),
.B(n_141),
.C(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_118),
.A2(n_119),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_118),
.A2(n_119),
.B1(n_175),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_167),
.C(n_175),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_119),
.B(n_147),
.C(n_151),
.Y(n_299)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_132),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_131),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_134),
.Y(n_288)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_138),
.A2(n_139),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_138),
.A2(n_139),
.B1(n_228),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_222),
.C(n_228),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_139),
.B(n_198),
.C(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_141),
.A2(n_142),
.B1(n_189),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_141),
.A2(n_142),
.B1(n_173),
.B2(n_186),
.Y(n_265)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_142),
.B(n_173),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_158),
.C(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_145),
.B(n_146),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_179),
.B(n_296),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_177),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_161),
.B(n_177),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_162),
.B(n_164),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_166),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_167),
.A2(n_168),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_173),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_200),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_173),
.A2(n_186),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_173),
.B(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_291),
.B(n_295),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_218),
.B(n_277),
.C(n_290),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_207),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_182),
.B(n_207),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_192),
.B2(n_206),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_185),
.B(n_191),
.C(n_206),
.Y(n_278)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_204),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_197),
.A2(n_198),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_251),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_198)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.C(n_214),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_209),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_214),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_216),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_276),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_237),
.B(n_275),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_234),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_221),
.B(n_234),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_222),
.A2(n_223),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_268),
.B(n_274),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_262),
.B(n_267),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_254),
.B(n_261),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_246),
.B(n_253),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_243),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_250),
.B(n_252),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_256),
.Y(n_261)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_289),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_287),
.C(n_289),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);


endmodule