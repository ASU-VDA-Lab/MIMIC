module fake_aes_10419_n_29 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_5), .Y(n_14) );
BUFx8_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
AND3x1_ASAP7_75t_SL g20 ( .A(n_17), .B(n_0), .C(n_1), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx2_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
AO21x2_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_16), .B(n_20), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND4xp25_ASAP7_75t_L g25 ( .A(n_24), .B(n_18), .C(n_15), .D(n_14), .Y(n_25) );
NOR3xp33_ASAP7_75t_SL g26 ( .A(n_25), .B(n_15), .C(n_3), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_26), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_2), .A3(n_4), .B1(n_6), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_29) );
endmodule