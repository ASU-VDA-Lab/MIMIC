module fake_jpeg_13874_n_498 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_498);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_498;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_53),
.Y(n_123)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_54),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_55),
.B(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_15),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_13),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_59),
.B(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_13),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_65),
.Y(n_122)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_67),
.B(n_71),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_29),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_77),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx2_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_81),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_89),
.Y(n_119)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_34),
.B(n_0),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx16f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx11_ASAP7_75t_SL g95 ( 
.A(n_46),
.Y(n_95)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_102),
.B(n_103),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_67),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_35),
.B1(n_25),
.B2(n_23),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_124),
.B1(n_155),
.B2(n_39),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_47),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_36),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_29),
.B(n_39),
.C(n_40),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_66),
.B(n_38),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_150),
.Y(n_189)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_38),
.Y(n_150)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_95),
.A2(n_45),
.B(n_44),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_93),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_72),
.A2(n_25),
.B1(n_35),
.B2(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_74),
.B(n_34),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_36),
.Y(n_199)
);

CKINVDCx12_ASAP7_75t_R g158 ( 
.A(n_109),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g253 ( 
.A(n_158),
.Y(n_253)
);

CKINVDCx12_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_159),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_160),
.Y(n_224)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_161),
.Y(n_257)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_25),
.B1(n_35),
.B2(n_44),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_164),
.A2(n_172),
.B1(n_205),
.B2(n_30),
.Y(n_229)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_201),
.B1(n_133),
.B2(n_137),
.Y(n_228)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_47),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_191),
.Y(n_220)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_105),
.A2(n_58),
.B1(n_52),
.B2(n_40),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_202),
.B1(n_212),
.B2(n_213),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_171),
.B(n_183),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_25),
.B1(n_35),
.B2(n_45),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_99),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_175),
.B(n_188),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g182 ( 
.A(n_101),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx9p33_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_120),
.B(n_99),
.Y(n_188)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_91),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_193),
.Y(n_221)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_117),
.A2(n_30),
.B(n_62),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_203),
.B(n_128),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_144),
.B(n_32),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_125),
.B(n_91),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_204),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_108),
.A2(n_76),
.B1(n_86),
.B2(n_85),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_122),
.A2(n_30),
.B(n_93),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_18),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_114),
.A2(n_79),
.B1(n_40),
.B2(n_18),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_129),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_208),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_210),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_132),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_139),
.Y(n_233)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_146),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_215),
.B(n_219),
.C(n_249),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_216),
.B(n_228),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_136),
.C(n_111),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_229),
.A2(n_244),
.B1(n_213),
.B2(n_202),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_233),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_166),
.A2(n_106),
.B1(n_139),
.B2(n_137),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_235),
.A2(n_236),
.B1(n_177),
.B2(n_167),
.Y(n_290)
);

AO21x2_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_106),
.B(n_133),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_168),
.B(n_126),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_248),
.Y(n_271)
);

OAI22x1_ASAP7_75t_SL g244 ( 
.A1(n_170),
.A2(n_105),
.B1(n_68),
.B2(n_50),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_151),
.B1(n_104),
.B2(n_149),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_180),
.B1(n_190),
.B2(n_161),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_104),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_112),
.C(n_151),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_112),
.B1(n_191),
.B2(n_165),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_203),
.A2(n_96),
.B1(n_65),
.B2(n_107),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_42),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_207),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_178),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_249),
.C(n_242),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_261),
.A2(n_301),
.B1(n_252),
.B2(n_234),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_220),
.B(n_42),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_262),
.B(n_263),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_32),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_186),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_270),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_160),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_268),
.B(n_269),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_240),
.B(n_24),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_226),
.B(n_179),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_169),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_273),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_222),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_275),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_162),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_278),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_255),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_24),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_280),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_247),
.B(n_233),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_283),
.A2(n_292),
.B1(n_214),
.B2(n_224),
.Y(n_322)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

OR2x2_ASAP7_75t_SL g288 ( 
.A(n_216),
.B(n_163),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_231),
.B1(n_244),
.B2(n_236),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_206),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_299),
.A3(n_224),
.B1(n_243),
.B2(n_236),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_184),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_194),
.B(n_253),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_227),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_238),
.B(n_212),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_209),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_217),
.B(n_174),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_229),
.A2(n_185),
.B1(n_176),
.B2(n_107),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_320),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_246),
.Y(n_305)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_271),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_308),
.A2(n_332),
.B1(n_276),
.B2(n_293),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_251),
.C(n_230),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_318),
.C(n_320),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_264),
.A2(n_218),
.B1(n_236),
.B2(n_243),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_321),
.B1(n_324),
.B2(n_336),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_326),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_223),
.C(n_230),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_254),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_287),
.A2(n_236),
.B1(n_254),
.B2(n_214),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

OAI22x1_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_227),
.B1(n_252),
.B2(n_245),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_223),
.B1(n_234),
.B2(n_65),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_274),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_287),
.A2(n_75),
.B1(n_69),
.B2(n_194),
.Y(n_336)
);

AO22x1_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_253),
.B1(n_225),
.B2(n_4),
.Y(n_337)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_337),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_286),
.A2(n_75),
.B1(n_69),
.B2(n_4),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_339),
.A2(n_276),
.B1(n_290),
.B2(n_284),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_323),
.B(n_269),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_340),
.B(n_346),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_267),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_343),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_310),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_345),
.B(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_315),
.B(n_262),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_347),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_263),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_348),
.B(n_349),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_312),
.B(n_279),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_299),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_313),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_L g391 ( 
.A1(n_351),
.A2(n_330),
.B(n_328),
.Y(n_391)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_356),
.A2(n_313),
.B1(n_319),
.B2(n_285),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_364),
.C(n_369),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_283),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_306),
.A2(n_284),
.B(n_271),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_361),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_275),
.Y(n_361)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

NOR2x1_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_305),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_319),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_295),
.C(n_265),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_307),
.B(n_281),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_367),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_306),
.A2(n_326),
.B1(n_332),
.B2(n_318),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_366),
.A2(n_324),
.B1(n_321),
.B2(n_317),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_303),
.B(n_266),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_305),
.B(n_289),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_370),
.B(n_336),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_371),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_366),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_387),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_354),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_381),
.B(n_353),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_358),
.C(n_364),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_386),
.C(n_388),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_357),
.B(n_370),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_368),
.C(n_356),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_329),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_342),
.A2(n_338),
.B1(n_316),
.B2(n_329),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_316),
.C(n_314),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_344),
.B1(n_368),
.B2(n_352),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_342),
.A2(n_319),
.B1(n_328),
.B2(n_330),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_282),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_393),
.A2(n_351),
.B(n_362),
.Y(n_413)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_396),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_397),
.A2(n_344),
.B(n_371),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_343),
.Y(n_400)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_374),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_406),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_385),
.Y(n_424)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_414),
.B1(n_416),
.B2(n_420),
.Y(n_429)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_409),
.A2(n_417),
.B1(n_380),
.B2(n_398),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_389),
.B(n_362),
.CI(n_363),
.CON(n_410),
.SN(n_410)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_410),
.A2(n_413),
.B1(n_421),
.B2(n_4),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_399),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_412),
.B(n_395),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_389),
.A2(n_397),
.B1(n_382),
.B2(n_373),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_372),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_415),
.Y(n_431)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_419),
.B(n_2),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_382),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_350),
.B1(n_341),
.B2(n_355),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_422),
.A2(n_2),
.B(n_3),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_296),
.C(n_225),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_375),
.C(n_386),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_427),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_377),
.B1(n_396),
.B2(n_379),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_425),
.A2(n_403),
.B1(n_401),
.B2(n_410),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_379),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_434),
.C(n_435),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_430),
.A2(n_434),
.B(n_438),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_423),
.C(n_405),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_432),
.B(n_433),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_392),
.C(n_387),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_376),
.C(n_378),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_376),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_441),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_2),
.C(n_3),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_440),
.C(n_442),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_5),
.C(n_7),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_437),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_448),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_431),
.B(n_411),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_446),
.B(n_450),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_407),
.C(n_412),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_408),
.C(n_422),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_456),
.C(n_5),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_429),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_455),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_11),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_439),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_406),
.C(n_402),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_457),
.A2(n_425),
.B1(n_433),
.B2(n_435),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_458),
.A2(n_461),
.B1(n_467),
.B2(n_447),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_442),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_463),
.Y(n_478)
);

FAx1_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_410),
.CI(n_424),
.CON(n_461),
.SN(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_457),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_468),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_448),
.A2(n_440),
.B(n_436),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_466),
.A2(n_470),
.B(n_447),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_452),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_445),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_7),
.C(n_8),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_464),
.A2(n_450),
.B(n_449),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_476),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_474),
.Y(n_485)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_462),
.A2(n_445),
.B(n_444),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_479),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_461),
.B(n_10),
.CI(n_8),
.CON(n_479),
.SN(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_466),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_480),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_478),
.B(n_459),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_486),
.A2(n_467),
.B1(n_470),
.B2(n_468),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_483),
.B(n_473),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_487),
.B(n_488),
.Y(n_492)
);

AOI31xp33_ASAP7_75t_L g488 ( 
.A1(n_482),
.A2(n_480),
.A3(n_461),
.B(n_474),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_477),
.C(n_475),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_490),
.Y(n_491)
);

AOI322xp5_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_481),
.A3(n_485),
.B1(n_489),
.B2(n_479),
.C1(n_484),
.C2(n_469),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_493),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_491),
.C(n_9),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_9),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_496),
.B(n_9),
.Y(n_497)
);

AO21x1_ASAP7_75t_L g498 ( 
.A1(n_497),
.A2(n_9),
.B(n_10),
.Y(n_498)
);


endmodule