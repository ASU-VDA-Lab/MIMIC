module fake_jpeg_2575_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_SL g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_5),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_27)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_9),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_21),
.B1(n_13),
.B2(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_11),
.B1(n_18),
.B2(n_14),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_36),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_29),
.Y(n_48)
);

AOI222xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_13),
.B1(n_21),
.B2(n_20),
.C1(n_16),
.C2(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_39)
);

OAI22x1_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_44),
.B1(n_32),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_54),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_29),
.B1(n_28),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_43),
.B1(n_32),
.B2(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_39),
.B1(n_44),
.B2(n_30),
.Y(n_68)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_30),
.C(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_67),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_57),
.B1(n_47),
.B2(n_45),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_68),
.B1(n_53),
.B2(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_65),
.B1(n_61),
.B2(n_60),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_55),
.C(n_54),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_72),
.C(n_74),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_51),
.C(n_52),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_38),
.B(n_51),
.C(n_56),
.D(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_77),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_30),
.C(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_84),
.B1(n_76),
.B2(n_32),
.C(n_5),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_67),
.C(n_63),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_32),
.C(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_72),
.B1(n_68),
.B2(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_88),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_81),
.C(n_78),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_78),
.C(n_3),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_2),
.B(n_5),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_93),
.C(n_94),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_98),
.B1(n_6),
.B2(n_7),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_6),
.C(n_8),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_6),
.Y(n_101)
);


endmodule