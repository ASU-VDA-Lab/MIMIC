module fake_jpeg_3402_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_7),
.Y(n_23)
);

AO22x1_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_20),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_18),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_12),
.B1(n_11),
.B2(n_23),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_35),
.B(n_37),
.C(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_19),
.B1(n_22),
.B2(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_24),
.B(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_36),
.B(n_38),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_36),
.B(n_35),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_32),
.B1(n_37),
.B2(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_52),
.B(n_42),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_35),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_31),
.B1(n_17),
.B2(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_54),
.C(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_44),
.B(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_66),
.Y(n_67)
);

AO221x1_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_53),
.B1(n_48),
.B2(n_2),
.C(n_3),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_7),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_8),
.B(n_64),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_70),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_64),
.B(n_8),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_0),
.B(n_1),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.C(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_1),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_2),
.CI(n_75),
.CON(n_77),
.SN(n_77)
);


endmodule