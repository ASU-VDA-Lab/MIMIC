module fake_jpeg_6309_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_20),
.B1(n_46),
.B2(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_39),
.B1(n_38),
.B2(n_40),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_62),
.B1(n_69),
.B2(n_71),
.Y(n_83)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_30),
.C(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_55),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_33),
.B1(n_21),
.B2(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_64),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_20),
.B1(n_31),
.B2(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_19),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_22),
.B(n_28),
.C(n_18),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_72),
.Y(n_97)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx2_ASAP7_75t_SL g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_59),
.B1(n_53),
.B2(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_43),
.B(n_25),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_59),
.B1(n_53),
.B2(n_79),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_47),
.C(n_61),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_115),
.C(n_35),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_54),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_108),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_72),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_121),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_62),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_113),
.B(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_37),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_66),
.C(n_45),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_66),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_45),
.B(n_32),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_93),
.B(n_89),
.C(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_134),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_60),
.B1(n_63),
.B2(n_52),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_136),
.B1(n_153),
.B2(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_90),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_115),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_105),
.B(n_110),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_58),
.B1(n_64),
.B2(n_73),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_140),
.B1(n_143),
.B2(n_145),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_99),
.B1(n_56),
.B2(n_79),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_74),
.B1(n_95),
.B2(n_94),
.Y(n_143)
);

OAI211xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_36),
.B(n_35),
.C(n_37),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_74),
.B1(n_97),
.B2(n_41),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_147),
.B1(n_103),
.B2(n_102),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_39),
.B1(n_46),
.B2(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_17),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_17),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_124),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_104),
.A2(n_46),
.B1(n_39),
.B2(n_37),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_108),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_124),
.B1(n_119),
.B2(n_117),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_176),
.B1(n_177),
.B2(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_162),
.C(n_164),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_126),
.C(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_127),
.B(n_116),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_170),
.B(n_162),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_122),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_174),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_128),
.B(n_125),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_137),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_172),
.C(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_111),
.C(n_35),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_119),
.B1(n_103),
.B2(n_102),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_175),
.B1(n_155),
.B2(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_120),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_36),
.B1(n_33),
.B2(n_21),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_17),
.C(n_25),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_33),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_132),
.Y(n_186)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_154),
.B1(n_141),
.B2(n_149),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_24),
.B1(n_28),
.B2(n_17),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_185),
.B(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_203),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_199),
.B1(n_156),
.B2(n_183),
.Y(n_218)
);

XOR2x2_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_129),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_198),
.C(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_200),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_202),
.B(n_207),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_24),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_163),
.B1(n_157),
.B2(n_158),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_144),
.B(n_130),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_130),
.B(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_181),
.B1(n_154),
.B2(n_177),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_146),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_206),
.C(n_208),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_145),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_141),
.B(n_143),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_131),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_166),
.B1(n_169),
.B2(n_158),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_32),
.B(n_26),
.Y(n_224)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_231),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_161),
.B1(n_175),
.B2(n_156),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_230),
.B1(n_202),
.B2(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_216),
.Y(n_256)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_224),
.B1(n_191),
.B2(n_184),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_17),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_229),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_225),
.B(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_28),
.B1(n_32),
.B2(n_25),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_248),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_249),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_252),
.B1(n_0),
.B2(n_1),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_220),
.B1(n_224),
.B2(n_215),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_226),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_194),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_201),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_213),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_211),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_238),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_187),
.B1(n_190),
.B2(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_233),
.B(n_222),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_257),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_225),
.B(n_207),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_190),
.C(n_192),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_223),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_260),
.A2(n_274),
.B(n_271),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_228),
.B1(n_235),
.B2(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_239),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_211),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_269),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_246),
.B1(n_242),
.B2(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_273),
.C(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_230),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_192),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_256),
.B1(n_254),
.B2(n_239),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_15),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_15),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_14),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_14),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_242),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_275),
.A2(n_240),
.B1(n_238),
.B2(n_243),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_281),
.B1(n_265),
.B2(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_252),
.C(n_244),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_0),
.C(n_1),
.Y(n_289)
);

OAI221xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.C(n_11),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_1),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_13),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_299),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_262),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_303),
.C(n_306),
.Y(n_310)
);

OAI321xp33_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_262),
.A3(n_273),
.B1(n_13),
.B2(n_12),
.C(n_10),
.Y(n_300)
);

AOI31xp33_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_302),
.A3(n_4),
.B(n_5),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_1),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_304),
.B(n_3),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_10),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_2),
.C(n_3),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_2),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_3),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_2),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_280),
.C(n_289),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_314),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_308),
.A2(n_286),
.B1(n_294),
.B2(n_280),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_303),
.B(n_297),
.C(n_8),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_298),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_6),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_4),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_6),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_4),
.C(n_5),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_310),
.B(n_312),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_331),
.B(n_332),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_316),
.B(n_319),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_6),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_6),
.B(n_7),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_320),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_330),
.B(n_329),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_334),
.B(n_8),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_7),
.B(n_9),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_9),
.Y(n_340)
);


endmodule