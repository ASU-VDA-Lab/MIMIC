module fake_jpeg_3727_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_23),
.C(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_31),
.B1(n_18),
.B2(n_28),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_58),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_27),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_47),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_41),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_57),
.B1(n_53),
.B2(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_69),
.B1(n_79),
.B2(n_83),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_74),
.B(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_24),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_32),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_91),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_50),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_55),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_110),
.B(n_68),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_103),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_40),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_82),
.C(n_77),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_49),
.B1(n_56),
.B2(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_71),
.B1(n_85),
.B2(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_49),
.Y(n_103)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_73),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_75),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_0),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_56),
.B1(n_55),
.B2(n_32),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_76),
.B1(n_63),
.B2(n_86),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_120),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_76),
.B1(n_72),
.B2(n_63),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_119),
.B1(n_125),
.B2(n_135),
.Y(n_141)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_124),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_129),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_127),
.B(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_75),
.B(n_74),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_65),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_97),
.B1(n_100),
.B2(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_98),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_66),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_1),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_96),
.B(n_87),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_79),
.B1(n_69),
.B2(n_56),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_104),
.B1(n_97),
.B2(n_100),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_32),
.B1(n_21),
.B2(n_20),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_109),
.C(n_105),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_95),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_105),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_156),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_110),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_159),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_160),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_111),
.A2(n_133),
.B(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_38),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_119),
.C(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_1),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_93),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_165),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_89),
.B1(n_130),
.B2(n_113),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_158),
.B1(n_146),
.B2(n_141),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_130),
.B(n_93),
.C(n_135),
.D(n_94),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_41),
.A3(n_40),
.B1(n_38),
.B2(n_94),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2x1_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_90),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_159),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_156),
.C(n_142),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_41),
.B(n_40),
.C(n_38),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_21),
.Y(n_183)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_138),
.C(n_145),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_191),
.C(n_175),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_138),
.C(n_153),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_197),
.B1(n_202),
.B2(n_182),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_174),
.A2(n_15),
.B1(n_12),
.B2(n_5),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_2),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_12),
.B1(n_4),
.B2(n_6),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_169),
.B1(n_179),
.B2(n_164),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_212),
.Y(n_220)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_166),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_170),
.B(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_191),
.C(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_170),
.B1(n_176),
.B2(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_204),
.B1(n_210),
.B2(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_187),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_225),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.C(n_227),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_192),
.B1(n_196),
.B2(n_201),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_216),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_193),
.C(n_201),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_234),
.C(n_236),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_219),
.B(n_212),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_233),
.B(n_221),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_223),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_215),
.C(n_211),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_241),
.C(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_229),
.B(n_220),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_206),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_209),
.B(n_6),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_2),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_250)
);

NOR3xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_11),
.C(n_246),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_11),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_249),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_251),
.Y(n_256)
);


endmodule