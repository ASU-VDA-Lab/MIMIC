module fake_jpeg_1535_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_12),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_34),
.B(n_37),
.C(n_38),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_35),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_56),
.Y(n_66)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_44),
.B1(n_49),
.B2(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_45),
.B1(n_44),
.B2(n_33),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_67),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_1),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_34),
.CI(n_38),
.CON(n_67),
.SN(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_3),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_1),
.B(n_2),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_55),
.CON(n_79),
.SN(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_2),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_84),
.Y(n_94)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_20),
.C(n_30),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_62),
.C(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_64),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_67),
.C(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_61),
.B1(n_51),
.B2(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_93),
.B1(n_8),
.B2(n_9),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_17),
.C(n_29),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_60),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_4),
.B(n_5),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_106),
.B1(n_96),
.B2(n_10),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_103),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_96),
.C(n_15),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_100),
.B1(n_107),
.B2(n_111),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_114),
.B(n_113),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_106),
.B(n_101),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_116),
.B(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_25),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_26),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_28),
.Y(n_121)
);


endmodule