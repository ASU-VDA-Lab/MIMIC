module fake_jpeg_1201_n_607 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_607);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_607;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_75),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_65),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_67),
.B(n_72),
.Y(n_158)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_28),
.B(n_10),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_19),
.C(n_2),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g154 ( 
.A(n_77),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_93),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_88),
.Y(n_117)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_31),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_54),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_99),
.Y(n_119)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_20),
.B(n_11),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_11),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_101),
.B(n_104),
.Y(n_149)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_11),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_22),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_109),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_39),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_111),
.B(n_0),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_115),
.B(n_170),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_54),
.B1(n_20),
.B2(n_29),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_123),
.A2(n_131),
.B1(n_135),
.B2(n_138),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_77),
.A2(n_52),
.B1(n_53),
.B2(n_44),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_23),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_142),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_77),
.A2(n_52),
.B1(n_53),
.B2(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_52),
.B1(n_53),
.B2(n_44),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_65),
.A2(n_32),
.B1(n_54),
.B2(n_47),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_146),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_32),
.B1(n_54),
.B2(n_47),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_60),
.B(n_29),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_72),
.A2(n_50),
.B1(n_47),
.B2(n_37),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_32),
.B1(n_50),
.B2(n_27),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_50),
.B1(n_37),
.B2(n_25),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_150),
.A2(n_66),
.B1(n_63),
.B2(n_97),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_61),
.B(n_25),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_159),
.B(n_168),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_62),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_162),
.A2(n_176),
.B1(n_4),
.B2(n_7),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_76),
.B(n_23),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_21),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_169),
.B(n_177),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_73),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_106),
.B(n_19),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_67),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_190),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_179),
.B(n_185),
.Y(n_249)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_120),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_209),
.Y(n_246)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_182),
.Y(n_298)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_187),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_68),
.B1(n_70),
.B2(n_56),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_212),
.B1(n_216),
.B2(n_230),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_149),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_55),
.Y(n_190)
);

OR2x4_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_86),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_191),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_105),
.C(n_102),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_192),
.B(n_229),
.C(n_239),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_98),
.B1(n_87),
.B2(n_89),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_194),
.Y(n_285)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_160),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_131),
.A2(n_86),
.B(n_74),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_197),
.A2(n_235),
.B(n_12),
.Y(n_274)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_112),
.B(n_84),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_215),
.Y(n_266)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

OR2x2_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_92),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_204),
.Y(n_297)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_205),
.Y(n_279)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_59),
.B1(n_103),
.B2(n_100),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_79),
.B1(n_64),
.B2(n_111),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_214),
.B(n_219),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_118),
.B(n_91),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_141),
.A2(n_85),
.B1(n_82),
.B2(n_69),
.Y(n_216)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_217),
.Y(n_294)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_221),
.Y(n_251)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_223),
.Y(n_270)
);

INVx4_ASAP7_75t_SL g223 ( 
.A(n_121),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_225),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_226),
.B(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_227),
.B(n_228),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_117),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_137),
.B(n_2),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_144),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_136),
.B(n_153),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_166),
.Y(n_268)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_233),
.Y(n_281)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_135),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_174),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_237),
.Y(n_282)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_151),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_234),
.B(n_197),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_129),
.B(n_7),
.C(n_8),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_140),
.A2(n_139),
.B1(n_146),
.B2(n_138),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_176),
.B1(n_166),
.B2(n_163),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_174),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_13),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_164),
.B(n_12),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_242),
.B(n_171),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_162),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_244),
.B(n_259),
.C(n_263),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_188),
.A2(n_163),
.B1(n_153),
.B2(n_133),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_245),
.A2(n_260),
.B1(n_284),
.B2(n_291),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_256),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_129),
.C(n_164),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_161),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_261),
.B(n_265),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_161),
.C(n_113),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_191),
.B(n_184),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_268),
.B(n_213),
.Y(n_339)
);

AOI32xp33_ASAP7_75t_L g269 ( 
.A1(n_198),
.A2(n_113),
.A3(n_171),
.B1(n_130),
.B2(n_157),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_273),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_274),
.A2(n_16),
.B(n_194),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_202),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_278),
.Y(n_312)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_211),
.A2(n_157),
.A3(n_152),
.B1(n_133),
.B2(n_15),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_211),
.A2(n_152),
.B1(n_13),
.B2(n_14),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_200),
.B(n_12),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_296),
.Y(n_309)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_192),
.B(n_12),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_229),
.C(n_242),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_209),
.A2(n_18),
.B1(n_14),
.B2(n_15),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_236),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_206),
.A2(n_18),
.B(n_15),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_242),
.B(n_239),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_228),
.B(n_215),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_231),
.B(n_16),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_179),
.Y(n_317)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_300),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_186),
.B(n_204),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_301),
.A2(n_331),
.B(n_337),
.Y(n_373)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_304),
.B(n_313),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_324),
.Y(n_367)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_264),
.A2(n_226),
.B1(n_229),
.B2(n_238),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_314),
.A2(n_316),
.B1(n_284),
.B2(n_291),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_275),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_315),
.B(n_317),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_264),
.A2(n_199),
.B1(n_217),
.B2(n_214),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_225),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_324),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_250),
.B(n_263),
.C(n_247),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_323),
.C(n_334),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_224),
.C(n_219),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_288),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_257),
.A2(n_233),
.B1(n_180),
.B2(n_201),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_325),
.A2(n_336),
.B1(n_341),
.B2(n_346),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_275),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_326),
.B(n_340),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_222),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_327),
.B(n_330),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_254),
.B(n_261),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_244),
.A2(n_181),
.B(n_221),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_227),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_333),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_187),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_247),
.B(n_237),
.C(n_183),
.Y(n_334)
);

NOR2x1p5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_182),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_338),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_257),
.A2(n_208),
.B1(n_203),
.B2(n_195),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_256),
.A2(n_297),
.B(n_274),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_223),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_243),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_218),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_253),
.A2(n_232),
.B1(n_210),
.B2(n_207),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_342),
.A2(n_292),
.B1(n_251),
.B2(n_290),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_265),
.B(n_16),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_343),
.B(n_344),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_205),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_260),
.A2(n_252),
.B1(n_295),
.B2(n_246),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_299),
.B(n_259),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_348),
.B(n_349),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_270),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_249),
.C(n_246),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_243),
.C(n_262),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_249),
.B(n_282),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_351),
.B(n_303),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_252),
.A2(n_246),
.B1(n_269),
.B2(n_278),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_352),
.A2(n_290),
.B1(n_289),
.B2(n_292),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_273),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_354),
.B(n_385),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_310),
.A2(n_273),
.B1(n_294),
.B2(n_245),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_356),
.A2(n_357),
.B1(n_366),
.B2(n_371),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_294),
.B1(n_282),
.B2(n_270),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_358),
.A2(n_378),
.B1(n_392),
.B2(n_325),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_310),
.A2(n_267),
.B1(n_271),
.B2(n_255),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_379),
.C(n_391),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_346),
.A2(n_322),
.B1(n_319),
.B2(n_333),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_332),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_381),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_251),
.B(n_283),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_374),
.A2(n_335),
.B(n_337),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_322),
.A2(n_271),
.B1(n_267),
.B2(n_255),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_384),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_320),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_301),
.A2(n_289),
.B1(n_285),
.B2(n_262),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_283),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_398),
.Y(n_412)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_305),
.B(n_272),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_314),
.A2(n_279),
.B1(n_285),
.B2(n_336),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_334),
.B(n_285),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_396),
.C(n_351),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_323),
.C(n_331),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_330),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_343),
.Y(n_432)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_403),
.A2(n_410),
.B(n_433),
.Y(n_448)
);

AOI22x1_ASAP7_75t_L g405 ( 
.A1(n_371),
.A2(n_318),
.B1(n_311),
.B2(n_302),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_405),
.A2(n_419),
.B1(n_432),
.B2(n_368),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_408),
.B(n_413),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_409),
.A2(n_423),
.B1(n_400),
.B2(n_366),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_397),
.A2(n_335),
.B(n_303),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_386),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_350),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_428),
.C(n_439),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_370),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_422),
.Y(n_458)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

AOI22x1_ASAP7_75t_L g419 ( 
.A1(n_397),
.A2(n_307),
.B1(n_316),
.B2(n_335),
.Y(n_419)
);

AO22x2_ASAP7_75t_L g420 ( 
.A1(n_362),
.A2(n_349),
.B1(n_304),
.B2(n_326),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_388),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_358),
.A2(n_327),
.B1(n_312),
.B2(n_306),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_382),
.Y(n_425)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_395),
.B(n_309),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_426),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_309),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_435),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_373),
.B(n_308),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_396),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_313),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_431),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g433 ( 
.A(n_373),
.B(n_315),
.CI(n_312),
.CON(n_433),
.SN(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_340),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_389),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_438),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_359),
.B(n_339),
.C(n_338),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_363),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g506 ( 
.A(n_440),
.B(n_444),
.C(n_461),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_375),
.B(n_374),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_442),
.A2(n_468),
.B(n_471),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_328),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_405),
.A2(n_378),
.B1(n_357),
.B2(n_376),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_400),
.A2(n_375),
.B1(n_364),
.B2(n_376),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_453),
.A2(n_475),
.B1(n_409),
.B2(n_411),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_385),
.C(n_379),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_460),
.C(n_465),
.Y(n_481)
);

OAI31xp33_ASAP7_75t_L g487 ( 
.A1(n_456),
.A2(n_419),
.A3(n_424),
.B(n_433),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_354),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_459),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_393),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_428),
.B(n_394),
.C(n_364),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_363),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_394),
.C(n_355),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_406),
.A2(n_392),
.B(n_355),
.Y(n_468)
);

OAI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_406),
.A2(n_353),
.B1(n_390),
.B2(n_317),
.Y(n_469)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_469),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_410),
.A2(n_384),
.B(n_356),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_473),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_407),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_474),
.B(n_383),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_411),
.A2(n_405),
.B1(n_420),
.B2(n_412),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_478),
.A2(n_480),
.B1(n_501),
.B2(n_471),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_439),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_479),
.B(n_495),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_456),
.A2(n_423),
.B1(n_435),
.B2(n_420),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_463),
.A2(n_420),
.B(n_419),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_483),
.A2(n_446),
.B(n_449),
.C(n_470),
.Y(n_527)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_485),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_429),
.C(n_434),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_493),
.C(n_500),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_487),
.B(n_490),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_402),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_488),
.B(n_497),
.Y(n_512)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_436),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_492),
.Y(n_511)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_473),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_451),
.B(n_401),
.C(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_498),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_433),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_344),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_447),
.B(n_300),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_458),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_505),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_459),
.B(n_328),
.C(n_444),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_467),
.B(n_460),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_502),
.B(n_503),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_466),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_482),
.A2(n_448),
.B(n_463),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_509),
.A2(n_510),
.B(n_532),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_482),
.A2(n_448),
.B(n_442),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_455),
.C(n_465),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_516),
.C(n_528),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_455),
.C(n_461),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_453),
.Y(n_517)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_517),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_441),
.Y(n_518)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_518),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_520),
.A2(n_523),
.B1(n_486),
.B2(n_481),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_476),
.A2(n_475),
.B1(n_468),
.B2(n_446),
.Y(n_523)
);

OAI322xp33_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_495),
.A3(n_506),
.B1(n_440),
.B2(n_477),
.C1(n_487),
.C2(n_479),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_506),
.Y(n_542)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_493),
.B(n_441),
.C(n_449),
.Y(n_528)
);

OA21x2_ASAP7_75t_SL g529 ( 
.A1(n_480),
.A2(n_470),
.B(n_466),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_529),
.B(n_531),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_505),
.Y(n_530)
);

CKINVDCx14_ASAP7_75t_R g543 ( 
.A(n_530),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_484),
.B(n_496),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_483),
.A2(n_501),
.B(n_478),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_514),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_533),
.B(n_539),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_500),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_512),
.B(n_522),
.Y(n_540)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_540),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_542),
.A2(n_526),
.B(n_519),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_519),
.A2(n_517),
.B1(n_509),
.B2(n_508),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_544),
.A2(n_523),
.B1(n_517),
.B2(n_532),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_515),
.B(n_492),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_545),
.B(n_551),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_510),
.A2(n_489),
.B(n_491),
.Y(n_546)
);

NAND2x1_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_548),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_547),
.A2(n_524),
.B1(n_530),
.B2(n_513),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_507),
.B(n_481),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_550),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_521),
.B(n_525),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_512),
.B(n_522),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_528),
.B(n_507),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_552),
.B(n_553),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_514),
.C(n_525),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_554),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_518),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_555),
.B(n_562),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_520),
.C(n_529),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_SL g581 ( 
.A(n_558),
.B(n_569),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_559),
.A2(n_560),
.B1(n_534),
.B2(n_547),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_535),
.B(n_515),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_517),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_564),
.B(n_536),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_544),
.A2(n_531),
.B1(n_511),
.B2(n_527),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_565),
.B(n_566),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_524),
.C(n_513),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_548),
.Y(n_570)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_570),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_527),
.C(n_533),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_571),
.B(n_539),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_554),
.A2(n_541),
.B1(n_543),
.B2(n_537),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_575),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_556),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_577),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_564),
.A2(n_538),
.B1(n_549),
.B2(n_536),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_580),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_565),
.A2(n_534),
.B(n_538),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_579),
.B(n_583),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_571),
.B(n_545),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_585),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_542),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_573),
.B(n_561),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_587),
.B(n_591),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_582),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_585),
.B(n_563),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_592),
.B(n_593),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_574),
.B(n_557),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_594),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_595),
.B(n_581),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_586),
.B(n_572),
.Y(n_596)
);

OAI21xp33_ASAP7_75t_L g600 ( 
.A1(n_596),
.A2(n_598),
.B(n_567),
.Y(n_600)
);

AOI221xp5_ASAP7_75t_L g598 ( 
.A1(n_588),
.A2(n_575),
.B1(n_579),
.B2(n_577),
.C(n_558),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_600),
.A2(n_601),
.B(n_602),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_599),
.B(n_590),
.C(n_589),
.Y(n_602)
);

AOI221xp5_ASAP7_75t_L g603 ( 
.A1(n_600),
.A2(n_588),
.B1(n_597),
.B2(n_564),
.C(n_567),
.Y(n_603)
);

OA21x2_ASAP7_75t_SL g605 ( 
.A1(n_603),
.A2(n_589),
.B(n_578),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_605),
.A2(n_604),
.B(n_560),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_606),
.B(n_568),
.Y(n_607)
);


endmodule