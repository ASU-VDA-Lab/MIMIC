module fake_jpeg_12372_n_557 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_557);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_124),
.Y(n_139)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_8),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_65),
.B(n_121),
.Y(n_177)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_22),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g161 ( 
.A(n_68),
.Y(n_161)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_73),
.Y(n_147)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_76),
.Y(n_163)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_77),
.Y(n_181)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_79),
.B(n_116),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_39),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_89),
.A2(n_34),
.B1(n_52),
.B2(n_49),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_8),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_92),
.B(n_100),
.Y(n_169)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_7),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_29),
.B(n_7),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_30),
.B(n_9),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_36),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_55),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_29),
.B(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_123),
.B(n_13),
.Y(n_202)
);

BUFx4f_ASAP7_75t_SL g124 ( 
.A(n_44),
.Y(n_124)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_57),
.CON(n_125),
.SN(n_125)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_125),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_65),
.A2(n_22),
.B1(n_41),
.B2(n_54),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_SL g129 ( 
.A(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_129),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_70),
.A2(n_22),
.B1(n_42),
.B2(n_36),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_70),
.A2(n_36),
.B1(n_42),
.B2(n_50),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_57),
.B1(n_43),
.B2(n_54),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_135),
.A2(n_154),
.B1(n_189),
.B2(n_200),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_42),
.B1(n_36),
.B2(n_55),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_34),
.B(n_43),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_187),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_69),
.A2(n_71),
.B1(n_86),
.B2(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_155),
.A2(n_166),
.B1(n_179),
.B2(n_118),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_52),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_156),
.B(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_49),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_68),
.B(n_37),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_162),
.B(n_27),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_120),
.A2(n_42),
.B1(n_50),
.B2(n_48),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_168),
.B(n_183),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_61),
.A2(n_26),
.B1(n_48),
.B2(n_47),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_64),
.B(n_37),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_89),
.A2(n_47),
.B1(n_46),
.B2(n_35),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_72),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_80),
.A2(n_46),
.B1(n_35),
.B2(n_32),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_202),
.B(n_13),
.Y(n_245)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_205),
.Y(n_313)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_207),
.Y(n_314)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_211),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_229),
.Y(n_291)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_219),
.Y(n_306)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_221),
.Y(n_298)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_223),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_224),
.A2(n_236),
.B1(n_265),
.B2(n_269),
.Y(n_311)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_160),
.A2(n_117),
.B1(n_115),
.B2(n_113),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_226),
.A2(n_175),
.B1(n_182),
.B2(n_188),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_141),
.C(n_165),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_235),
.C(n_246),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_131),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_242),
.Y(n_300)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_233),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_234),
.B(n_237),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_177),
.B(n_27),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_32),
.B1(n_181),
.B2(n_126),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_16),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_16),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_238),
.B(n_240),
.Y(n_293)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_139),
.B(n_16),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g241 ( 
.A(n_181),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_241),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_131),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_171),
.B(n_105),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_243),
.A2(n_161),
.B(n_176),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_104),
.B1(n_98),
.B2(n_97),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_266),
.B1(n_155),
.B2(n_179),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_245),
.B(n_249),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_148),
.B(n_0),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_194),
.A2(n_15),
.B(n_1),
.C(n_2),
.Y(n_248)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_158),
.A3(n_146),
.B1(n_161),
.B2(n_142),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_192),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_133),
.Y(n_250)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_147),
.Y(n_251)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_257),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_164),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_255),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_130),
.A2(n_94),
.B1(n_88),
.B2(n_87),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_256),
.A2(n_0),
.B1(n_203),
.B2(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_140),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_259),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_197),
.B(n_4),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_260),
.Y(n_297)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_262),
.B(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_172),
.B(n_4),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_149),
.A2(n_44),
.B1(n_6),
.B2(n_11),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_167),
.A2(n_44),
.B1(n_6),
.B2(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_159),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_267),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_192),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_216),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_270),
.A2(n_272),
.B1(n_0),
.B2(n_209),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_132),
.B(n_16),
.C(n_15),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_164),
.CI(n_192),
.CON(n_284),
.SN(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_163),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_244),
.A2(n_176),
.B1(n_130),
.B2(n_174),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_274),
.A2(n_289),
.B1(n_292),
.B2(n_295),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_296),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_212),
.A2(n_166),
.B1(n_136),
.B2(n_134),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_255),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_212),
.A2(n_161),
.B1(n_184),
.B2(n_167),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_205),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_208),
.A2(n_174),
.B1(n_146),
.B2(n_142),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_318),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_294),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_214),
.A2(n_175),
.B1(n_182),
.B2(n_188),
.Y(n_295)
);

FAx1_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_0),
.CI(n_203),
.CON(n_308),
.SN(n_308)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_248),
.B(n_271),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_0),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_230),
.B(n_235),
.CI(n_208),
.CON(n_327),
.SN(n_327)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_327),
.B(n_275),
.CI(n_318),
.CON(n_341),
.SN(n_341)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_332),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_341),
.Y(n_380)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_309),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_307),
.B(n_303),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_285),
.A2(n_277),
.B1(n_295),
.B2(n_290),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_342),
.A2(n_359),
.B1(n_362),
.B2(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_311),
.A2(n_273),
.B1(n_261),
.B2(n_243),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_368),
.B1(n_279),
.B2(n_323),
.Y(n_373)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_286),
.A2(n_222),
.B(n_252),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_348),
.A2(n_355),
.B(n_291),
.Y(n_375)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_293),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_350),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_315),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_215),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_353),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_218),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_275),
.B(n_228),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_357),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_308),
.A2(n_264),
.B(n_250),
.Y(n_355)
);

INVx3_ASAP7_75t_SL g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_320),
.A2(n_206),
.A3(n_217),
.B1(n_225),
.B2(n_262),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_254),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_358),
.B(n_364),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_308),
.A2(n_284),
.B1(n_292),
.B2(n_287),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_360),
.Y(n_386)
);

NOR3xp33_ASAP7_75t_SL g361 ( 
.A(n_282),
.B(n_209),
.C(n_241),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_361),
.B(n_365),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_310),
.A2(n_223),
.B1(n_233),
.B2(n_207),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_284),
.A2(n_232),
.B1(n_239),
.B2(n_213),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_247),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_227),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_304),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_368),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_298),
.B(n_229),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_367),
.B(n_288),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_322),
.A2(n_227),
.B1(n_324),
.B2(n_323),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_322),
.C(n_324),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_372),
.B(n_400),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_373),
.A2(n_389),
.B(n_332),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_342),
.A2(n_313),
.B1(n_314),
.B2(n_304),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_374),
.A2(n_382),
.B1(n_384),
.B2(n_393),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_375),
.A2(n_366),
.B(n_299),
.Y(n_429)
);

OAI211xp5_ASAP7_75t_SL g378 ( 
.A1(n_346),
.A2(n_297),
.B(n_313),
.C(n_314),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g425 ( 
.A1(n_378),
.A2(n_330),
.A3(n_329),
.B1(n_316),
.B2(n_288),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_339),
.A2(n_305),
.B1(n_297),
.B2(n_283),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_339),
.A2(n_302),
.B1(n_280),
.B2(n_283),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_359),
.A2(n_306),
.B1(n_317),
.B2(n_281),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_346),
.A2(n_307),
.B1(n_303),
.B2(n_306),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_394),
.A2(n_328),
.B1(n_363),
.B2(n_353),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_403),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_317),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_399),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_299),
.C(n_312),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_281),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_405),
.A2(n_409),
.B1(n_413),
.B2(n_420),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_398),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_416),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_332),
.B(n_355),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_392),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_408),
.A2(n_410),
.B(n_415),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_394),
.A2(n_347),
.B1(n_338),
.B2(n_348),
.Y(n_409)
);

A2O1A1O1Ixp25_ASAP7_75t_L g411 ( 
.A1(n_380),
.A2(n_341),
.B(n_351),
.C(n_361),
.D(n_344),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_417),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_402),
.A2(n_340),
.B1(n_334),
.B2(n_341),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_392),
.A2(n_345),
.B(n_343),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_379),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_379),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_395),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_419),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_369),
.A2(n_340),
.B1(n_356),
.B2(n_357),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_382),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_386),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_423),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_386),
.Y(n_423)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

A2O1A1O1Ixp25_ASAP7_75t_L g426 ( 
.A1(n_380),
.A2(n_366),
.B(n_356),
.C(n_335),
.D(n_316),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_432),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_399),
.Y(n_427)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_427),
.Y(n_451)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_393),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_373),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_430),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_276),
.B(n_312),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_372),
.C(n_403),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_437),
.C(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_413),
.C(n_424),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_402),
.C(n_390),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_433),
.A2(n_376),
.B1(n_370),
.B2(n_369),
.Y(n_442)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_390),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_454),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_400),
.C(n_381),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_453),
.C(n_455),
.Y(n_483)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_381),
.C(n_396),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_410),
.B(n_405),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_396),
.C(n_378),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_418),
.A2(n_420),
.B1(n_421),
.B2(n_374),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_456),
.A2(n_433),
.B1(n_427),
.B2(n_406),
.Y(n_461)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_449),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_463),
.Y(n_495)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_449),
.Y(n_467)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_467),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_408),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_475),
.Y(n_486)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_437),
.B(n_411),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_472),
.B(n_478),
.Y(n_499)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_452),
.Y(n_473)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_473),
.Y(n_497)
);

OAI31xp33_ASAP7_75t_L g474 ( 
.A1(n_444),
.A2(n_416),
.A3(n_417),
.B(n_425),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_474),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_448),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_423),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_480),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_439),
.A2(n_454),
.B1(n_453),
.B2(n_446),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_477),
.A2(n_438),
.B1(n_446),
.B2(n_412),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_415),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_479),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_422),
.Y(n_480)
);

OA22x2_ASAP7_75t_L g481 ( 
.A1(n_456),
.A2(n_432),
.B1(n_426),
.B2(n_384),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_481),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_412),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_482),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_391),
.C(n_436),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_370),
.Y(n_503)
);

FAx1_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_455),
.CI(n_443),
.CON(n_492),
.SN(n_492)
);

AO21x1_ASAP7_75t_L g515 ( 
.A1(n_492),
.A2(n_466),
.B(n_481),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_445),
.C(n_443),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_494),
.B(n_501),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g500 ( 
.A1(n_480),
.A2(n_467),
.B(n_445),
.Y(n_500)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_500),
.Y(n_506)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_483),
.C(n_464),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_505),
.C(n_510),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_483),
.C(n_464),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_481),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_481),
.Y(n_526)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_508),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_484),
.A2(n_462),
.B1(n_466),
.B2(n_468),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_509),
.A2(n_515),
.B1(n_488),
.B2(n_500),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_468),
.C(n_475),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_469),
.C(n_472),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_499),
.C(n_484),
.Y(n_522)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_513),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_391),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_438),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_514),
.A2(n_493),
.B1(n_485),
.B2(n_489),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_517),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_499),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_522),
.B(n_523),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_506),
.A2(n_485),
.B(n_488),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_525),
.Y(n_534)
);

O2A1O1Ixp33_ASAP7_75t_SL g525 ( 
.A1(n_507),
.A2(n_474),
.B(n_482),
.C(n_492),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_516),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_504),
.B(n_492),
.C(n_447),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_505),
.C(n_458),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_515),
.B1(n_509),
.B2(n_502),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_528),
.B(n_530),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_521),
.A2(n_497),
.B1(n_511),
.B2(n_507),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_537),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_523),
.A2(n_497),
.B1(n_465),
.B2(n_498),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_532),
.B(n_533),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_525),
.A2(n_457),
.B1(n_426),
.B2(n_428),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_526),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_377),
.C(n_419),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_537),
.B(n_519),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_539),
.B(n_542),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_531),
.A2(n_527),
.B(n_522),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_540),
.A2(n_544),
.B(n_536),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_529),
.A2(n_517),
.B(n_526),
.Y(n_544)
);

AO21x1_ASAP7_75t_L g550 ( 
.A1(n_545),
.A2(n_547),
.B(n_538),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_543),
.B(n_520),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_SL g548 ( 
.A(n_541),
.B(n_534),
.C(n_536),
.Y(n_548)
);

NOR2x1_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_388),
.Y(n_551)
);

O2A1O1Ixp33_ASAP7_75t_SL g549 ( 
.A1(n_546),
.A2(n_538),
.B(n_533),
.C(n_387),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_550),
.Y(n_553)
);

AOI321xp33_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_383),
.A3(n_385),
.B1(n_377),
.B2(n_401),
.C(n_431),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_552),
.A2(n_385),
.B(n_401),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_553),
.C(n_387),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_388),
.C(n_397),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_556),
.A2(n_337),
.B(n_276),
.Y(n_557)
);


endmodule