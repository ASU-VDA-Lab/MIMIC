module fake_jpeg_723_n_496 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_496);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_496;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_56),
.Y(n_170)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_60),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_86),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_62),
.Y(n_185)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_30),
.B1(n_43),
.B2(n_29),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_79),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_87),
.B(n_116),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

BUFx12f_ASAP7_75t_SL g99 ( 
.A(n_32),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_29),
.B(n_8),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_110),
.Y(n_151)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_20),
.B(n_8),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_114),
.B(n_4),
.Y(n_176)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_112),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_19),
.B(n_8),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_4),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_0),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_24),
.B1(n_47),
.B2(n_40),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_120),
.A2(n_128),
.B1(n_129),
.B2(n_134),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_18),
.B1(n_47),
.B2(n_34),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_124),
.A2(n_138),
.B1(n_147),
.B2(n_154),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_60),
.A2(n_18),
.B1(n_34),
.B2(n_40),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_66),
.A2(n_18),
.B1(n_52),
.B2(n_49),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_114),
.B(n_112),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_0),
.C(n_1),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_56),
.A2(n_19),
.B1(n_43),
.B2(n_36),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_133),
.A2(n_150),
.B1(n_155),
.B2(n_1),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_52),
.B1(n_38),
.B2(n_49),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_39),
.B1(n_38),
.B2(n_50),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_141),
.A2(n_146),
.B(n_185),
.C(n_128),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_144),
.B(n_176),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_39),
.B1(n_46),
.B2(n_50),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_72),
.A2(n_36),
.B1(n_35),
.B2(n_50),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_76),
.A2(n_35),
.B1(n_25),
.B2(n_2),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_78),
.A2(n_46),
.B1(n_25),
.B2(n_11),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_79),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_80),
.A2(n_5),
.B1(n_12),
.B2(n_11),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_166),
.B(n_137),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_77),
.B(n_4),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_188),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_68),
.A2(n_85),
.B1(n_110),
.B2(n_106),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_186),
.B1(n_191),
.B2(n_0),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_82),
.A2(n_91),
.B1(n_88),
.B2(n_113),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_101),
.B(n_5),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_102),
.A2(n_10),
.B1(n_12),
.B2(n_16),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_107),
.B(n_12),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_111),
.B(n_16),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_197),
.A2(n_232),
.B1(n_251),
.B2(n_254),
.Y(n_264)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_198),
.Y(n_279)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_132),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_200),
.B(n_215),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_203),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_204),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_0),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_205),
.B(n_207),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_137),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_206),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_270)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_211),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_213),
.Y(n_299)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_160),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_139),
.Y(n_219)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_225),
.A2(n_229),
.B1(n_233),
.B2(n_242),
.Y(n_292)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_142),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_120),
.A2(n_150),
.B1(n_186),
.B2(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_234),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_142),
.A2(n_124),
.B1(n_146),
.B2(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_238),
.Y(n_293)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_143),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_135),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_239),
.B(n_240),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_241),
.B(n_243),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_141),
.A2(n_119),
.B1(n_134),
.B2(n_191),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_143),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_141),
.A2(n_130),
.B1(n_160),
.B2(n_173),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_250),
.B1(n_260),
.B2(n_223),
.Y(n_291)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_153),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_195),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_252),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_127),
.B(n_175),
.C(n_163),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_165),
.C(n_183),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_129),
.A2(n_172),
.B1(n_122),
.B2(n_183),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_162),
.A2(n_184),
.B1(n_182),
.B2(n_172),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_148),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_145),
.A2(n_164),
.B(n_169),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_253),
.A2(n_226),
.B(n_257),
.Y(n_297)
);

AOI22x1_ASAP7_75t_L g254 ( 
.A1(n_168),
.A2(n_187),
.B1(n_196),
.B2(n_195),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_148),
.A2(n_189),
.B1(n_122),
.B2(n_161),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_253),
.B1(n_220),
.B2(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_257),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_126),
.B(n_161),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_259),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_126),
.B(n_196),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_263),
.B(n_265),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_196),
.C(n_189),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_228),
.B1(n_233),
.B2(n_201),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_266),
.A2(n_275),
.B1(n_296),
.B2(n_288),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g339 ( 
.A1(n_267),
.A2(n_282),
.B1(n_301),
.B2(n_284),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_174),
.B1(n_235),
.B2(n_207),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_280),
.B1(n_291),
.B2(n_302),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_174),
.CI(n_216),
.CON(n_273),
.SN(n_273)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_273),
.B(n_261),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_212),
.A2(n_202),
.B1(n_254),
.B2(n_231),
.Y(n_275)
);

AOI32xp33_ASAP7_75t_L g276 ( 
.A1(n_211),
.A2(n_218),
.A3(n_238),
.B1(n_243),
.B2(n_217),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_263),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_214),
.B1(n_199),
.B2(n_208),
.Y(n_280)
);

AO22x1_ASAP7_75t_L g296 ( 
.A1(n_209),
.A2(n_210),
.B1(n_221),
.B2(n_204),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_297),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_241),
.B1(n_227),
.B2(n_240),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_224),
.A2(n_201),
.B(n_207),
.C(n_131),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_303),
.B(n_307),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_308),
.A2(n_266),
.B1(n_264),
.B2(n_275),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_309),
.A2(n_329),
.B1(n_343),
.B2(n_310),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_277),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_321),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_271),
.B1(n_308),
.B2(n_273),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_313),
.A2(n_315),
.B1(n_325),
.B2(n_326),
.Y(n_352)
);

NOR3xp33_ASAP7_75t_SL g346 ( 
.A(n_314),
.B(n_327),
.C(n_316),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_273),
.B1(n_267),
.B2(n_297),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_262),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_316),
.B(n_340),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_303),
.B(n_298),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_317),
.A2(n_319),
.B(n_345),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_304),
.A2(n_298),
.B(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_322),
.Y(n_350)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_265),
.A2(n_280),
.B1(n_307),
.B2(n_269),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_324),
.A2(n_335),
.B1(n_337),
.B2(n_333),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_262),
.A2(n_276),
.B1(n_300),
.B2(n_299),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_299),
.B1(n_302),
.B2(n_272),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_331),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_295),
.A2(n_281),
.B1(n_294),
.B2(n_290),
.Y(n_329)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_334),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_261),
.A2(n_268),
.B1(n_272),
.B2(n_283),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_282),
.A2(n_295),
.B1(n_294),
.B2(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_339),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_286),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_281),
.B(n_279),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_289),
.A2(n_286),
.B1(n_285),
.B2(n_287),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_289),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_318),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_285),
.A2(n_292),
.B(n_297),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_318),
.C(n_340),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_344),
.Y(n_384)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_310),
.B(n_345),
.C(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_357),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_342),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_356),
.B(n_368),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_309),
.A2(n_314),
.B1(n_331),
.B2(n_324),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_320),
.B1(n_330),
.B2(n_313),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_360),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_310),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_310),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_369),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g365 ( 
.A1(n_325),
.A2(n_311),
.B(n_326),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_311),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_317),
.A3(n_330),
.B1(n_328),
.B2(n_319),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_312),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_370),
.B(n_372),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_337),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_373),
.B(n_374),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_318),
.B(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_385),
.Y(n_404)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_398),
.B1(n_365),
.B2(n_368),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_391),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_394),
.C(n_395),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_355),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_363),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_392),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_360),
.A2(n_329),
.B(n_343),
.Y(n_389)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_389),
.A2(n_351),
.B(n_361),
.C(n_353),
.Y(n_420)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_358),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_338),
.C(n_341),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_367),
.C(n_374),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_364),
.C(n_348),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_323),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_397),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_354),
.A2(n_323),
.B1(n_332),
.B2(n_363),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_365),
.B1(n_386),
.B2(n_387),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_401),
.A2(n_406),
.B1(n_398),
.B2(n_376),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_397),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_414),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_352),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_408),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_382),
.A2(n_365),
.B1(n_372),
.B2(n_352),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_407),
.A2(n_379),
.B1(n_381),
.B2(n_388),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_367),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_413),
.C(n_415),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_348),
.C(n_350),
.Y(n_413)
);

XOR2x2_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_369),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_396),
.C(n_395),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_375),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_420),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_382),
.A2(n_359),
.B1(n_373),
.B2(n_356),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_377),
.B1(n_375),
.B2(n_385),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_350),
.C(n_353),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_399),
.C(n_393),
.Y(n_440)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_422),
.Y(n_425)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_427),
.A2(n_418),
.B1(n_406),
.B2(n_401),
.Y(n_443)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_422),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_419),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_435),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_430),
.A2(n_433),
.B1(n_426),
.B2(n_425),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_404),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_408),
.B(n_415),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_440),
.Y(n_442)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_392),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_438),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_399),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_439),
.Y(n_447)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_380),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_443),
.A2(n_448),
.B1(n_411),
.B2(n_420),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_452),
.B1(n_453),
.B2(n_439),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_427),
.A2(n_410),
.B1(n_404),
.B2(n_405),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_400),
.C(n_412),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_451),
.C(n_434),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_413),
.C(n_414),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_430),
.A2(n_433),
.B1(n_426),
.B2(n_436),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_424),
.A2(n_388),
.B1(n_393),
.B2(n_409),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_440),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_455),
.B(n_464),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_463),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_457),
.Y(n_468)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_452),
.A2(n_383),
.B1(n_421),
.B2(n_409),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_461),
.B1(n_444),
.B2(n_448),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_460),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_445),
.A2(n_411),
.B1(n_378),
.B2(n_437),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_423),
.C(n_403),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_465),
.C(n_442),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_443),
.A2(n_346),
.B1(n_351),
.B2(n_389),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_429),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_423),
.C(n_419),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_471),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_442),
.C(n_447),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_456),
.C(n_462),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_459),
.A2(n_453),
.B(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_474),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_475),
.B(n_481),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_463),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_479),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_457),
.C(n_461),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_458),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g485 ( 
.A(n_480),
.B(n_464),
.C(n_441),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_460),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_L g482 ( 
.A1(n_476),
.A2(n_467),
.B(n_469),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_482),
.B(n_486),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_474),
.B(n_466),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_484),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_485),
.B(n_446),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_487),
.A2(n_488),
.B(n_480),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_483),
.C(n_477),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_490),
.A2(n_491),
.B(n_468),
.Y(n_492)
);

OAI321xp33_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_441),
.A3(n_468),
.B1(n_481),
.B2(n_390),
.C(n_378),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_391),
.C(n_361),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_361),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_361),
.C(n_391),
.Y(n_496)
);


endmodule