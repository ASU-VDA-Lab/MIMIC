module fake_jpeg_22209_n_282 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_25),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_20),
.B1(n_25),
.B2(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_20),
.B1(n_34),
.B2(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_64),
.B1(n_29),
.B2(n_26),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_31),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_34),
.B1(n_19),
.B2(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_33),
.B1(n_21),
.B2(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_50),
.C(n_49),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_66),
.A2(n_23),
.B(n_65),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_75),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_R g70 ( 
.A(n_48),
.B(n_23),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_70),
.B(n_99),
.C(n_101),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_60),
.B1(n_51),
.B2(n_23),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_76),
.B(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_81),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_94),
.B1(n_97),
.B2(n_60),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_30),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_93),
.B1(n_85),
.B2(n_88),
.Y(n_109)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_21),
.B1(n_31),
.B2(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_29),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_38),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_100),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_21),
.Y(n_100)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_58),
.B(n_23),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_42),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_121),
.C(n_122),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_71),
.B1(n_90),
.B2(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_114),
.B1(n_117),
.B2(n_93),
.Y(n_145)
);

XOR2x1_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_78),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_118),
.B(n_73),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_60),
.B1(n_54),
.B2(n_5),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_23),
.B(n_4),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_3),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_127),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_53),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_4),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_130),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_67),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_91),
.B1(n_79),
.B2(n_74),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_141),
.B1(n_145),
.B2(n_113),
.Y(n_172)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_140),
.Y(n_176)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_74),
.B1(n_72),
.B2(n_99),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_68),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_111),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_154),
.B(n_97),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_68),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_158),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_155),
.B1(n_122),
.B2(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_128),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_92),
.B(n_86),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_86),
.B1(n_81),
.B2(n_84),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_98),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_138),
.B1(n_150),
.B2(n_136),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_104),
.C(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_167),
.C(n_171),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_121),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_164),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_127),
.B(n_112),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_172),
.B(n_177),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_113),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_129),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_128),
.C(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_98),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_65),
.B(n_53),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_5),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_186),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_6),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_131),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_193),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_144),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_162),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_201),
.B1(n_191),
.B2(n_159),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_143),
.B(n_146),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_202),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_155),
.B1(n_139),
.B2(n_8),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_203),
.B1(n_185),
.B2(n_182),
.Y(n_215)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_172),
.B1(n_161),
.B2(n_170),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_16),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_186),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_178),
.B1(n_174),
.B2(n_170),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_215),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_216),
.B1(n_219),
.B2(n_200),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_223),
.B(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_164),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.C(n_227),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_168),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_168),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_227),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_224),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_189),
.A3(n_192),
.B1(n_209),
.B2(n_195),
.C1(n_203),
.C2(n_194),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_175),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_192),
.B1(n_220),
.B2(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_197),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_226),
.B(n_10),
.Y(n_248)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_171),
.B1(n_208),
.B2(n_11),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_189),
.C(n_209),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_8),
.C(n_10),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_254),
.C(n_14),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_242),
.C(n_231),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_236),
.C(n_230),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_13),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_260),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_261),
.C(n_249),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_235),
.C(n_228),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_228),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_261),
.B(n_263),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_246),
.C(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_244),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_258),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_256),
.B(n_257),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_274),
.B(n_272),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_258),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_267),
.B(n_245),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_15),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_278),
.C(n_15),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_15),
.Y(n_282)
);


endmodule