module fake_jpeg_29744_n_366 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_366);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_366;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_48),
.B(n_49),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_55),
.Y(n_99)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g56 ( 
.A(n_16),
.B(n_14),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_58),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_59),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_24),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_74),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_0),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_4),
.C(n_5),
.Y(n_116)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_32),
.Y(n_83)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_9),
.B1(n_10),
.B2(n_74),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_80),
.B1(n_62),
.B2(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_84),
.A2(n_90),
.B1(n_71),
.B2(n_48),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_15),
.B1(n_29),
.B2(n_34),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_15),
.B1(n_29),
.B2(n_34),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_97),
.B1(n_106),
.B2(n_108),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_35),
.B1(n_29),
.B2(n_15),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_35),
.B1(n_29),
.B2(n_15),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_32),
.B1(n_37),
.B2(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_38),
.B1(n_23),
.B2(n_28),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_102),
.A2(n_105),
.B1(n_110),
.B2(n_112),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_38),
.B(n_23),
.C(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_81),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_21),
.B1(n_36),
.B2(n_33),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_21),
.B1(n_33),
.B2(n_30),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_37),
.B1(n_30),
.B2(n_11),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_9),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_122),
.B1(n_104),
.B2(n_113),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_47),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_110),
.B1(n_102),
.B2(n_107),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_10),
.B(n_68),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_65),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_128),
.C(n_109),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_53),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_57),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_57),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_149),
.Y(n_185)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_143),
.Y(n_189)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_115),
.B1(n_119),
.B2(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_60),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_107),
.B(n_77),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_164),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_87),
.A2(n_50),
.B1(n_63),
.B2(n_54),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_160),
.B1(n_114),
.B2(n_128),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_163),
.B(n_131),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_166),
.B1(n_171),
.B2(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_52),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_48),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_126),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_162),
.B(n_168),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_97),
.A2(n_124),
.B(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_167),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_92),
.A2(n_112),
.B1(n_87),
.B2(n_93),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_100),
.B(n_99),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_103),
.B(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_89),
.B(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_173),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_93),
.A2(n_123),
.B1(n_91),
.B2(n_114),
.Y(n_171)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_141),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_133),
.Y(n_215)
);

AO21x1_ASAP7_75t_SL g226 ( 
.A1(n_180),
.A2(n_201),
.B(n_144),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_198),
.B1(n_199),
.B2(n_177),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_196),
.B1(n_184),
.B2(n_179),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_89),
.B1(n_119),
.B2(n_115),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_109),
.A3(n_114),
.B1(n_128),
.B2(n_137),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_212),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_161),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_141),
.A2(n_158),
.B1(n_163),
.B2(n_160),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_158),
.A2(n_150),
.B1(n_164),
.B2(n_130),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_130),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_151),
.B(n_156),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_206),
.B(n_197),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_138),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_140),
.B(n_149),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_212),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_154),
.A2(n_153),
.B1(n_173),
.B2(n_143),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_174),
.B1(n_167),
.B2(n_145),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_135),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_191),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_226),
.B(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_134),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

AO21x2_ASAP7_75t_L g221 ( 
.A1(n_180),
.A2(n_167),
.B(n_172),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_231),
.B1(n_187),
.B2(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_175),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_228),
.A2(n_232),
.B1(n_204),
.B2(n_189),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_197),
.B(n_206),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_185),
.Y(n_260)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_244),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_198),
.C(n_177),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_245),
.C(n_185),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_175),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_201),
.B(n_186),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_177),
.B(n_178),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_194),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_231),
.A2(n_178),
.B1(n_192),
.B2(n_186),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_270),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_221),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_193),
.C(n_204),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_269),
.C(n_271),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_239),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_221),
.A2(n_194),
.B1(n_208),
.B2(n_193),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_239),
.B1(n_230),
.B2(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_176),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_210),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_283),
.B1(n_292),
.B2(n_260),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_226),
.C(n_227),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_278),
.B(n_246),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_235),
.B(n_215),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_257),
.B(n_246),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_262),
.A2(n_235),
.B1(n_221),
.B2(n_189),
.Y(n_278)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_248),
.B(n_214),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_228),
.B1(n_247),
.B2(n_254),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_215),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_286),
.C(n_289),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_223),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_210),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_287),
.Y(n_306)
);

INVx3_ASAP7_75t_SL g288 ( 
.A(n_262),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_293),
.B1(n_255),
.B2(n_253),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_222),
.C(n_216),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_271),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_221),
.B1(n_225),
.B2(n_189),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_295),
.A2(n_299),
.B(n_288),
.Y(n_323)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_302),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_248),
.B(n_272),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_294),
.B(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_294),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_250),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_258),
.B1(n_253),
.B2(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_258),
.B1(n_256),
.B2(n_255),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_312),
.B1(n_281),
.B2(n_280),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_251),
.B1(n_252),
.B2(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_265),
.B1(n_264),
.B2(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_265),
.B1(n_224),
.B2(n_188),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

BUFx12_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_327),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_284),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_322),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_275),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_295),
.B(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_330),
.A2(n_305),
.B(n_312),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_335),
.Y(n_340)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_302),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_321),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_337),
.A2(n_304),
.B(n_315),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_339),
.B(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_330),
.A2(n_326),
.B(n_325),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_346),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_320),
.B(n_323),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_306),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_347),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_306),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_325),
.B1(n_326),
.B2(n_332),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_349),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_310),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_351),
.A2(n_354),
.B(n_341),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_311),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_358),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_348),
.A2(n_307),
.B1(n_320),
.B2(n_303),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_356),
.A2(n_348),
.B1(n_357),
.B2(n_350),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_334),
.C(n_322),
.Y(n_358)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_359),
.A2(n_303),
.A3(n_349),
.B1(n_300),
.B2(n_319),
.C1(n_285),
.C2(n_297),
.Y(n_362)
);

AOI321xp33_ASAP7_75t_L g361 ( 
.A1(n_358),
.A2(n_353),
.A3(n_334),
.B1(n_346),
.B2(n_336),
.C(n_289),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_361),
.B(n_275),
.C(n_286),
.Y(n_363)
);

AOI321xp33_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_363),
.A3(n_360),
.B1(n_224),
.B2(n_205),
.C(n_188),
.Y(n_364)
);

AOI221xp5_ASAP7_75t_L g365 ( 
.A1(n_364),
.A2(n_175),
.B1(n_176),
.B2(n_182),
.C(n_353),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_182),
.Y(n_366)
);


endmodule