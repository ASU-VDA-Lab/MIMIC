module fake_jpeg_21748_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_54),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_43),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_60),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_15),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_67),
.A2(n_84),
.B1(n_95),
.B2(n_52),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_17),
.B1(n_29),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_97),
.B1(n_15),
.B2(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_82),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_78),
.B(n_81),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_42),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_18),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_41),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_38),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_32),
.B1(n_29),
.B2(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_43),
.B(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_16),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_115),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_47),
.B1(n_53),
.B2(n_49),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_105),
.A2(n_109),
.B1(n_114),
.B2(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_66),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_124),
.B1(n_141),
.B2(n_127),
.Y(n_151)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_111),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_125),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_63),
.B1(n_39),
.B2(n_51),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_126),
.B1(n_135),
.B2(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_129),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_65),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_46),
.B1(n_45),
.B2(n_36),
.Y(n_126)
);

FAx1_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_55),
.CI(n_18),
.CON(n_127),
.SN(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_132),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_137),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_37),
.B1(n_44),
.B2(n_17),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_21),
.Y(n_160)
);

BUFx2_ASAP7_75t_SL g140 ( 
.A(n_103),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_68),
.B(n_60),
.C(n_58),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_103),
.C(n_101),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_21),
.B1(n_16),
.B2(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_169),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_103),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_77),
.B(n_11),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_163),
.B(n_177),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_18),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_170),
.B(n_174),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_129),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_119),
.B(n_131),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_113),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_106),
.B1(n_110),
.B2(n_125),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_107),
.A2(n_73),
.B1(n_90),
.B2(n_70),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_101),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_178),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_100),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_179),
.B(n_181),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_109),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_208),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_112),
.B1(n_133),
.B2(n_76),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_186),
.B1(n_191),
.B2(n_196),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_164),
.B1(n_157),
.B2(n_112),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_214),
.B1(n_168),
.B2(n_176),
.Y(n_218)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_165),
.B1(n_167),
.B2(n_161),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_132),
.B1(n_120),
.B2(n_70),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_104),
.B1(n_116),
.B2(n_115),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_202),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_173),
.B1(n_151),
.B2(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_100),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_211),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_199),
.A2(n_203),
.B(n_210),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_21),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_200),
.B(n_2),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_108),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_160),
.B(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_33),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_148),
.B(n_122),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_205),
.B(n_163),
.Y(n_219)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_122),
.C(n_33),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_178),
.B1(n_153),
.B2(n_174),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_153),
.B1(n_174),
.B2(n_143),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_128),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_213),
.Y(n_233)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_168),
.B1(n_143),
.B2(n_150),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_96),
.C(n_103),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_96),
.C(n_150),
.Y(n_232)
);

INVxp33_ASAP7_75t_SL g216 ( 
.A(n_154),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_72),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_219),
.B(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_210),
.B1(n_182),
.B2(n_191),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_181),
.B1(n_209),
.B2(n_210),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_180),
.B(n_144),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_236),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_199),
.A2(n_23),
.B1(n_17),
.B2(n_156),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_128),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_33),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_187),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_118),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_72),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_118),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_96),
.Y(n_246)
);

NAND4xp25_ASAP7_75t_SL g247 ( 
.A(n_190),
.B(n_31),
.C(n_96),
.D(n_4),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_189),
.B(n_14),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_2),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_190),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_196),
.C(n_188),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_257),
.C(n_264),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_199),
.B(n_206),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_254),
.A2(n_246),
.B(n_233),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_226),
.B1(n_244),
.B2(n_236),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_206),
.C(n_192),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_265),
.Y(n_285)
);

OAI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_221),
.A2(n_195),
.B(n_213),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_SL g301 ( 
.A1(n_260),
.A2(n_263),
.B(n_280),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_195),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_262),
.B(n_243),
.Y(n_304)
);

AOI32xp33_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_185),
.A3(n_207),
.B1(n_13),
.B2(n_12),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_13),
.C(n_3),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_224),
.C(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_279),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_270),
.B(n_276),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_3),
.C(n_5),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_235),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_225),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_5),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_229),
.A2(n_234),
.B1(n_226),
.B2(n_223),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_241),
.A2(n_6),
.B(n_7),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_237),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_282),
.A2(n_287),
.B(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_298),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_288),
.A2(n_294),
.B1(n_296),
.B2(n_275),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_295),
.B(n_299),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_220),
.B1(n_233),
.B2(n_248),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_231),
.B(n_222),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_231),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_253),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_238),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_222),
.Y(n_302)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_279),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_310),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_267),
.B1(n_281),
.B2(n_258),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_311),
.A2(n_328),
.B1(n_282),
.B2(n_301),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_321),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_316),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_285),
.B(n_252),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_321),
.C(n_326),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_271),
.B1(n_228),
.B2(n_275),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_294),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_265),
.C(n_262),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_307),
.B1(n_298),
.B2(n_282),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_264),
.Y(n_324)
);

AOI21x1_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_295),
.B(n_304),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_283),
.B(n_266),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_228),
.B1(n_272),
.B2(n_255),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_337),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_300),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_283),
.C(n_297),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_343),
.C(n_323),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_312),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_341),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_313),
.Y(n_351)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_344),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_288),
.C(n_296),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_346),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_358),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_351),
.B(n_330),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_336),
.B(n_324),
.CI(n_311),
.CON(n_353),
.SN(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_354),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_314),
.B1(n_320),
.B2(n_308),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_345),
.A2(n_328),
.B(n_315),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_333),
.B(n_335),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_329),
.C(n_291),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_330),
.C(n_341),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_329),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_369),
.C(n_358),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_366),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_SL g365 ( 
.A(n_356),
.B(n_346),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_365),
.A2(n_357),
.B(n_352),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_332),
.C(n_331),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_332),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_368),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_306),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_337),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_370),
.A2(n_348),
.B(n_347),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_353),
.B(n_344),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_371),
.B(n_335),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_363),
.B(n_250),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_376),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_342),
.C(n_349),
.Y(n_374)
);

NOR3xp33_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_6),
.C(n_7),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g384 ( 
.A1(n_377),
.A2(n_247),
.B(n_250),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_364),
.A2(n_366),
.B1(n_360),
.B2(n_353),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_369),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_351),
.C(n_250),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_378),
.C(n_8),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_382),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_375),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_384),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_387),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_385),
.A2(n_6),
.B(n_8),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_389),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_388),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_392),
.A2(n_393),
.B1(n_391),
.B2(n_8),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_10),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_10),
.Y(n_396)
);


endmodule