module fake_jpeg_13975_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_51),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_61),
.Y(n_104)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_8),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_71),
.B(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_84),
.Y(n_143)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_35),
.Y(n_84)
);

INVx11_ASAP7_75t_SL g85 ( 
.A(n_29),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_89),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_26),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

OR2x4_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_43),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_38),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_15),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_99),
.C(n_60),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_38),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_21),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_25),
.B1(n_30),
.B2(n_37),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_41),
.B1(n_37),
.B2(n_30),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_106),
.A2(n_110),
.B1(n_112),
.B2(n_118),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_41),
.B1(n_30),
.B2(n_34),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_34),
.B1(n_36),
.B2(n_32),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_25),
.B1(n_32),
.B2(n_28),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_116),
.A2(n_117),
.B1(n_131),
.B2(n_122),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_36),
.B1(n_28),
.B2(n_23),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_91),
.B1(n_86),
.B2(n_80),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_127),
.A2(n_142),
.B1(n_149),
.B2(n_138),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_50),
.A2(n_56),
.B1(n_59),
.B2(n_52),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_102),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_49),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_150),
.B1(n_151),
.B2(n_128),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_67),
.A2(n_3),
.B1(n_6),
.B2(n_9),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_88),
.A2(n_12),
.B1(n_15),
.B2(n_97),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_85),
.A2(n_15),
.B1(n_62),
.B2(n_71),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_163),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_147),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_130),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_182),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_166),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_101),
.A3(n_124),
.B1(n_132),
.B2(n_109),
.Y(n_166)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_169),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_171),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_101),
.B(n_114),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_129),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_186),
.C(n_145),
.Y(n_206)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_123),
.B(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_183),
.Y(n_189)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_146),
.B1(n_120),
.B2(n_144),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_102),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_125),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_125),
.C(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_173),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_110),
.B1(n_127),
.B2(n_106),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_194),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_103),
.B(n_121),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_201),
.B(n_212),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_148),
.B(n_146),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_162),
.B1(n_174),
.B2(n_183),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_120),
.B(n_144),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_211),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_164),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_163),
.A2(n_162),
.B(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_218),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_194),
.B1(n_158),
.B2(n_168),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_180),
.B1(n_173),
.B2(n_177),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_191),
.B1(n_196),
.B2(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_190),
.B(n_160),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_179),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_232),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_210),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_204),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_170),
.B(n_167),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_233),
.B(n_188),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_182),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_200),
.B1(n_202),
.B2(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_243),
.B1(n_244),
.B2(n_248),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_250),
.B1(n_217),
.B2(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_214),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_199),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_196),
.B1(n_193),
.B2(n_204),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_218),
.B1(n_226),
.B2(n_233),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_203),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_222),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_203),
.B(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_231),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_233),
.B1(n_229),
.B2(n_232),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_267),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_263),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_227),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_265),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_216),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_234),
.C(n_243),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_273),
.C(n_276),
.Y(n_287)
);

XNOR2x2_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_239),
.B1(n_250),
.B2(n_240),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_253),
.B1(n_216),
.B2(n_255),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_244),
.C(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_239),
.C(n_249),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_250),
.B1(n_245),
.B2(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_245),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_288),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_259),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_286),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_254),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_277),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_257),
.C(n_254),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_270),
.C(n_237),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_255),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_271),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_272),
.B1(n_268),
.B2(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_296),
.A2(n_301),
.B1(n_230),
.B2(n_251),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_298),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_287),
.B(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_304),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_269),
.B1(n_268),
.B2(n_275),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_252),
.C(n_256),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_302),
.B(n_296),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_303),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_313),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_291),
.C(n_285),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.C(n_311),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_286),
.C(n_271),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_290),
.C(n_280),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_280),
.C(n_261),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_228),
.C(n_205),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_318),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_321),
.B(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_230),
.C(n_223),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_232),
.B(n_224),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_224),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_213),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_327),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_223),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_325),
.A2(n_223),
.B(n_215),
.C(n_195),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_223),
.C(n_205),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_331),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_195),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_213),
.Y(n_331)
);

OAI321xp33_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_324),
.A3(n_215),
.B1(n_194),
.B2(n_195),
.C(n_192),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_334),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_333),
.B(n_192),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_192),
.B(n_207),
.C(n_155),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_335),
.B(n_207),
.C(n_159),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_197),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_197),
.Y(n_340)
);


endmodule