module fake_jpeg_6124_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_13;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_28),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_21),
.B1(n_30),
.B2(n_17),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_57),
.B1(n_65),
.B2(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_30),
.B2(n_37),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_58),
.B(n_66),
.C(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_17),
.B1(n_30),
.B2(n_14),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_45),
.B1(n_14),
.B2(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_37),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_51),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_35),
.Y(n_102)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_86),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_49),
.C(n_50),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_49),
.C(n_31),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_29),
.B1(n_43),
.B2(n_40),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_59),
.B1(n_63),
.B2(n_56),
.Y(n_108)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_62),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_68),
.B(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_R g90 ( 
.A(n_76),
.B(n_66),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_92),
.B(n_95),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_58),
.CI(n_66),
.CON(n_91),
.SN(n_91)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_91),
.B(n_103),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_66),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_54),
.B1(n_57),
.B2(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_81),
.B1(n_70),
.B2(n_59),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_31),
.C(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_105),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_46),
.B1(n_48),
.B2(n_39),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_118),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_85),
.B(n_86),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_111),
.A2(n_115),
.B(n_130),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_95),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_120),
.B1(n_125),
.B2(n_98),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_35),
.B(n_46),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_129),
.C(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_121),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_52),
.B1(n_80),
.B2(n_46),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_98),
.B1(n_107),
.B2(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_48),
.B1(n_87),
.B2(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVxp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_82),
.C(n_72),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_88),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_102),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_138),
.C(n_145),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_152),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_88),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_117),
.B1(n_130),
.B2(n_113),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_98),
.B1(n_92),
.B2(n_91),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_144),
.B1(n_150),
.B2(n_22),
.Y(n_174)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_146),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_149),
.B1(n_130),
.B2(n_110),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_91),
.B(n_92),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_115),
.B(n_112),
.Y(n_155)
);

OAI22x1_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_91),
.B1(n_97),
.B2(n_83),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_94),
.C(n_96),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_94),
.B1(n_87),
.B2(n_89),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_96),
.B1(n_73),
.B2(n_78),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_142),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_165),
.Y(n_197)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_140),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_158),
.B(n_160),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_154),
.A2(n_145),
.B(n_148),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_129),
.B(n_118),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_129),
.B(n_127),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_163),
.B(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_16),
.B1(n_26),
.B2(n_33),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_136),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_109),
.C(n_87),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_170),
.C(n_173),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_137),
.C(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_174),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_109),
.B(n_25),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

BUFx4f_ASAP7_75t_SL g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_142),
.C(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_181),
.B(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_67),
.C(n_36),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_25),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_67),
.C(n_36),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_18),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_11),
.B(n_1),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_160),
.B(n_159),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_165),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_15),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_174),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_187),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_176),
.B1(n_178),
.B2(n_163),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_206),
.B1(n_213),
.B2(n_180),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_185),
.B(n_187),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_158),
.B1(n_170),
.B2(n_155),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_188),
.B(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_159),
.B1(n_167),
.B2(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_10),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_16),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_36),
.B1(n_33),
.B2(n_27),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_219),
.A2(n_194),
.B1(n_185),
.B2(n_200),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_223),
.B1(n_217),
.B2(n_1),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_180),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_226),
.C(n_228),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_197),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_189),
.C(n_199),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_233),
.C(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_27),
.C(n_26),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_27),
.C(n_19),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_218),
.C(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_230),
.Y(n_252)
);

AOI31xp33_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_204),
.A3(n_203),
.B(n_215),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_240),
.B(n_243),
.Y(n_261)
);

AO21x2_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_203),
.B(n_219),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_249),
.B1(n_220),
.B2(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_234),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_7),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_19),
.B1(n_23),
.B2(n_13),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_248),
.B1(n_6),
.B2(n_1),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_19),
.B1(n_23),
.B2(n_13),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_253),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_254),
.B(n_256),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_260),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_242),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_0),
.C(n_2),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_6),
.B(n_3),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_8),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_241),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_266),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_9),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_9),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_257),
.B(n_9),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_274),
.B(n_278),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_251),
.B(n_3),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_263),
.B(n_265),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_279),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_9),
.B(n_3),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_282),
.Y(n_284)
);

A2O1A1O1Ixp25_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_12),
.B(n_5),
.C(n_10),
.D(n_11),
.Y(n_283)
);

AOI321xp33_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_279),
.A3(n_5),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_280),
.B(n_5),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_284),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_12),
.B(n_0),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_12),
.CI(n_274),
.CON(n_289),
.SN(n_289)
);


endmodule