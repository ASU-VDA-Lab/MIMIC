module fake_netlist_6_3286_n_752 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_752);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_752;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_671;
wire n_726;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_43),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_24),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_87),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_18),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_63),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_39),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_72),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_76),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_50),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_93),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_15),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_14),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_44),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_69),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_55),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_38),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_51),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_78),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_45),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_34),
.Y(n_194)
);

INVxp33_ASAP7_75t_SL g195 ( 
.A(n_145),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_66),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_94),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_46),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_49),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_0),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_0),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_1),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_2),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_19),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_2),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_3),
.B(n_4),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_191),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_21),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_3),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_4),
.B(n_5),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_5),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_175),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_173),
.B1(n_172),
.B2(n_195),
.Y(n_237)
);

CKINVDCx11_ASAP7_75t_R g238 ( 
.A(n_187),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_9),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_187),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_167),
.B(n_9),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_10),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_10),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_156),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_186),
.B(n_11),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_11),
.Y(n_246)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_198),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_206),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_158),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_163),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_233),
.B(n_164),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_169),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

AO21x2_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_180),
.B(n_199),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_233),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_170),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_203),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_171),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_215),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_237),
.B(n_174),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_207),
.B(n_179),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_L g289 ( 
.A(n_226),
.B(n_181),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_240),
.B(n_185),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

CKINVDCx6p67_ASAP7_75t_R g293 ( 
.A(n_238),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_220),
.Y(n_294)
);

AND2x6_ASAP7_75t_SL g295 ( 
.A(n_252),
.B(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_232),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_255),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_285),
.B(n_207),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_243),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_214),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_214),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_282),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_216),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_242),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_188),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_253),
.B(n_189),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_253),
.B(n_193),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_253),
.B(n_194),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_285),
.B(n_208),
.Y(n_317)
);

CKINVDCx8_ASAP7_75t_R g318 ( 
.A(n_272),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_197),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_245),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_285),
.B(n_211),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_236),
.B1(n_246),
.B2(n_192),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_285),
.B(n_225),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_215),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_290),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_285),
.B(n_235),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_218),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_263),
.B(n_218),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_263),
.B(n_218),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_231),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_249),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_249),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_269),
.B(n_231),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_251),
.B(n_231),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_250),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_260),
.B(n_12),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

NOR2x1_ASAP7_75t_R g349 ( 
.A(n_293),
.B(n_224),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_254),
.B(n_22),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_277),
.B(n_23),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_277),
.B(n_25),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_254),
.B(n_26),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_289),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_355)
);

INVx8_ASAP7_75t_L g356 ( 
.A(n_247),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_269),
.B(n_15),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

BUFx4f_ASAP7_75t_L g359 ( 
.A(n_347),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_303),
.A2(n_300),
.B(n_301),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_301),
.A2(n_321),
.B(n_317),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_296),
.A2(n_291),
.B1(n_277),
.B2(n_272),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_269),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_317),
.A2(n_247),
.B(n_291),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_324),
.A2(n_311),
.B1(n_294),
.B2(n_304),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_256),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

O2A1O1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_266),
.B(n_288),
.C(n_284),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_283),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_294),
.Y(n_373)
);

AO21x1_ASAP7_75t_L g374 ( 
.A1(n_342),
.A2(n_291),
.B(n_277),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_321),
.A2(n_247),
.B(n_291),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_357),
.A2(n_288),
.B(n_284),
.C(n_259),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_L g377 ( 
.A1(n_342),
.A2(n_247),
.B(n_262),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_247),
.B(n_262),
.Y(n_378)
);

O2A1O1Ixp5_ASAP7_75t_L g379 ( 
.A1(n_330),
.A2(n_261),
.B(n_257),
.C(n_248),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_306),
.B(n_248),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_334),
.B(n_356),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_261),
.B(n_257),
.Y(n_383)
);

AOI21x1_ASAP7_75t_L g384 ( 
.A1(n_325),
.A2(n_259),
.B(n_256),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_274),
.B(n_97),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_318),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_327),
.B(n_274),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_16),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_27),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_224),
.C(n_17),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_329),
.A2(n_96),
.B1(n_152),
.B2(n_28),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_297),
.B(n_29),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_295),
.B(n_16),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_345),
.A2(n_355),
.B1(n_316),
.B2(n_315),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_319),
.B(n_30),
.Y(n_397)
);

BUFx12f_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_325),
.A2(n_99),
.B(n_31),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_314),
.B(n_17),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g401 ( 
.A1(n_351),
.A2(n_32),
.B(n_33),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_326),
.A2(n_36),
.B(n_37),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_313),
.A2(n_40),
.B1(n_41),
.B2(n_47),
.Y(n_404)
);

OAI21xp33_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_48),
.B(n_52),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_309),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_297),
.B(n_53),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_353),
.A2(n_56),
.B(n_58),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_299),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_299),
.Y(n_412)
);

BUFx4f_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_59),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_309),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_312),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_328),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_302),
.B(n_60),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_61),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_353),
.A2(n_62),
.B(n_65),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_302),
.Y(n_423)
);

O2A1O1Ixp5_ASAP7_75t_L g424 ( 
.A1(n_298),
.A2(n_67),
.B(n_68),
.C(n_70),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g425 ( 
.A1(n_384),
.A2(n_354),
.B(n_350),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_411),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_352),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_367),
.B(n_352),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_380),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_348),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_382),
.A2(n_348),
.B(n_343),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_379),
.A2(n_343),
.B(n_332),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_332),
.B(n_331),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_364),
.A2(n_71),
.B(n_73),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_362),
.A2(n_74),
.B(n_75),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_387),
.B(n_349),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g437 ( 
.A(n_366),
.B(n_77),
.C(n_80),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_372),
.A2(n_81),
.B(n_82),
.Y(n_438)
);

OAI22xp33_ASAP7_75t_L g439 ( 
.A1(n_359),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_439)
);

AO21x1_ASAP7_75t_L g440 ( 
.A1(n_364),
.A2(n_390),
.B(n_396),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_365),
.A2(n_153),
.B(n_90),
.Y(n_441)
);

AO31x2_ASAP7_75t_L g442 ( 
.A1(n_374),
.A2(n_88),
.A3(n_95),
.B(n_98),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_412),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_390),
.B(n_393),
.Y(n_444)
);

OR2x6_ASAP7_75t_L g445 ( 
.A(n_398),
.B(n_100),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_372),
.A2(n_101),
.B(n_102),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_359),
.B(n_103),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_375),
.A2(n_104),
.B(n_105),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_377),
.A2(n_106),
.B(n_108),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_383),
.A2(n_109),
.B(n_111),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_388),
.A2(n_113),
.B(n_114),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_396),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_376),
.A2(n_120),
.B(n_121),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_377),
.A2(n_122),
.B(n_125),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_369),
.A2(n_150),
.B(n_128),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_368),
.B(n_127),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_381),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_371),
.A2(n_129),
.B(n_130),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_369),
.A2(n_131),
.B(n_132),
.Y(n_462)
);

AO31x2_ASAP7_75t_L g463 ( 
.A1(n_401),
.A2(n_134),
.A3(n_135),
.B(n_137),
.Y(n_463)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_138),
.Y(n_464)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_406),
.A2(n_140),
.B(n_141),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_397),
.A2(n_143),
.B(n_147),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_419),
.A2(n_148),
.B(n_149),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_370),
.B(n_400),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_392),
.A2(n_402),
.B(n_413),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_410),
.B(n_414),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_406),
.A2(n_416),
.B(n_407),
.Y(n_473)
);

AO31x2_ASAP7_75t_L g474 ( 
.A1(n_363),
.A2(n_394),
.A3(n_420),
.B(n_415),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_405),
.A2(n_409),
.B(n_422),
.C(n_423),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g476 ( 
.A1(n_418),
.A2(n_421),
.B(n_415),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_SL g477 ( 
.A(n_395),
.B(n_404),
.C(n_363),
.Y(n_477)
);

OAI21x1_ASAP7_75t_SL g478 ( 
.A1(n_399),
.A2(n_385),
.B(n_394),
.Y(n_478)
);

AOI221xp5_ASAP7_75t_L g479 ( 
.A1(n_424),
.A2(n_403),
.B1(n_408),
.B2(n_420),
.C(n_416),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_408),
.Y(n_480)
);

NAND2x1p5_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_455),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_429),
.B(n_470),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_432),
.B(n_441),
.Y(n_484)
);

AO21x2_ASAP7_75t_L g485 ( 
.A1(n_440),
.A2(n_461),
.B(n_453),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_426),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_454),
.A2(n_434),
.B(n_428),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_465),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_472),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_477),
.A2(n_478),
.B(n_430),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_448),
.A2(n_433),
.B(n_450),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_425),
.A2(n_431),
.B(n_462),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_427),
.B(n_469),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_459),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_457),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_465),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_456),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_445),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_480),
.Y(n_502)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_449),
.A2(n_471),
.B(n_438),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_451),
.B(n_479),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_475),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

AO31x2_ASAP7_75t_L g507 ( 
.A1(n_452),
.A2(n_468),
.A3(n_446),
.B(n_474),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

BUFx2_ASAP7_75t_SL g509 ( 
.A(n_447),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_467),
.B(n_437),
.Y(n_510)
);

OAI221xp5_ASAP7_75t_SL g511 ( 
.A1(n_445),
.A2(n_439),
.B1(n_464),
.B2(n_444),
.C(n_436),
.Y(n_511)
);

O2A1O1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_444),
.A2(n_442),
.B(n_474),
.C(n_463),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_442),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_474),
.A2(n_373),
.B1(n_367),
.B2(n_429),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_442),
.A2(n_476),
.B(n_432),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_458),
.B(n_472),
.Y(n_516)
);

BUFx12f_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_459),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_473),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_429),
.B(n_361),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_429),
.B(n_373),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_373),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_426),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_429),
.B(n_373),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_520),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_523),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_523),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_482),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_514),
.A2(n_503),
.B(n_505),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_486),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_486),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_483),
.A2(n_521),
.B1(n_494),
.B2(n_520),
.Y(n_533)
);

BUFx2_ASAP7_75t_R g534 ( 
.A(n_499),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_499),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_495),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_484),
.B(n_493),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_498),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_498),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_489),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_505),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_518),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_522),
.A2(n_524),
.B1(n_494),
.B2(n_516),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_496),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_516),
.B(n_489),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_500),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_491),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_509),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_491),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_510),
.A2(n_487),
.B(n_512),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_501),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_491),
.B(n_485),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_506),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

NAND2x1_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_519),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_506),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_560),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_485),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_562),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_551),
.B(n_517),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_517),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_552),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_540),
.B(n_519),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_563),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_544),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_558),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_544),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_546),
.B(n_511),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_533),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_525),
.B(n_519),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_562),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_541),
.B(n_519),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_527),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_525),
.B(n_547),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_531),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_550),
.A2(n_485),
.B1(n_487),
.B2(n_506),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_531),
.B(n_513),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_538),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_542),
.A2(n_487),
.B1(n_508),
.B2(n_504),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_542),
.A2(n_487),
.B1(n_508),
.B2(n_519),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_549),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_528),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_529),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_L g594 ( 
.A1(n_558),
.A2(n_503),
.B(n_504),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_532),
.B(n_507),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_539),
.B(n_559),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_549),
.B(n_507),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_535),
.Y(n_601)
);

NOR2x1_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_488),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_554),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_559),
.B(n_507),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_558),
.B(n_507),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_603),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_603),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_569),
.Y(n_609)
);

NAND2x1p5_ASAP7_75t_SL g610 ( 
.A(n_602),
.B(n_556),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_599),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_569),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_583),
.B(n_545),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_598),
.B(n_530),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_530),
.Y(n_615)
);

INVx3_ASAP7_75t_SL g616 ( 
.A(n_599),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_572),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_599),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_507),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_595),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_595),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_600),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_549),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_567),
.B(n_548),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_577),
.B(n_515),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_564),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_597),
.B(n_561),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_566),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_571),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_565),
.B(n_537),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_605),
.B(n_543),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_571),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_605),
.B(n_543),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_576),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_579),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_577),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_637),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_637),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_585),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_622),
.B(n_575),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_627),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_634),
.B(n_597),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_635),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_635),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_622),
.B(n_575),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_609),
.B(n_591),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_634),
.B(n_589),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_624),
.Y(n_650)
);

AOI211xp5_ASAP7_75t_L g651 ( 
.A1(n_625),
.A2(n_568),
.B(n_594),
.C(n_578),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_L g652 ( 
.A(n_612),
.B(n_573),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_615),
.B(n_586),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_627),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_624),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_615),
.B(n_586),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_633),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_613),
.B(n_582),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_628),
.B(n_582),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_619),
.B(n_594),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_631),
.B(n_574),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_633),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_630),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_606),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_646),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_642),
.B(n_647),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_659),
.B(n_636),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_646),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_644),
.B(n_631),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_620),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_652),
.B(n_639),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_648),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_660),
.B(n_619),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_661),
.B(n_621),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_660),
.B(n_621),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_661),
.B(n_620),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_639),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_640),
.Y(n_678)
);

NOR2x1_ASAP7_75t_L g679 ( 
.A(n_667),
.B(n_636),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_675),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_672),
.B(n_638),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_666),
.B(n_651),
.C(n_658),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_673),
.B(n_638),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_SL g684 ( 
.A(n_671),
.B(n_534),
.Y(n_684)
);

OAI332xp33_ASAP7_75t_L g685 ( 
.A1(n_675),
.A2(n_662),
.A3(n_657),
.B1(n_645),
.B2(n_650),
.B3(n_655),
.C1(n_664),
.C2(n_663),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_670),
.A2(n_623),
.B1(n_573),
.B2(n_628),
.Y(n_686)
);

NAND2xp67_ASAP7_75t_L g687 ( 
.A(n_677),
.B(n_678),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_677),
.Y(n_688)
);

AOI21xp33_ASAP7_75t_SL g689 ( 
.A1(n_682),
.A2(n_681),
.B(n_680),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_683),
.B(n_669),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_682),
.A2(n_671),
.B(n_665),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_687),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_684),
.A2(n_573),
.B1(n_616),
.B2(n_618),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_691),
.A2(n_685),
.B(n_689),
.Y(n_694)
);

OAI21xp33_ASAP7_75t_SL g695 ( 
.A1(n_692),
.A2(n_679),
.B(n_686),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_693),
.A2(n_671),
.B(n_668),
.Y(n_696)
);

OAI32xp33_ASAP7_75t_L g697 ( 
.A1(n_690),
.A2(n_579),
.A3(n_601),
.B1(n_688),
.B2(n_649),
.Y(n_697)
);

OAI221xp5_ASAP7_75t_L g698 ( 
.A1(n_691),
.A2(n_601),
.B1(n_678),
.B2(n_573),
.C(n_616),
.Y(n_698)
);

OAI211xp5_ASAP7_75t_L g699 ( 
.A1(n_689),
.A2(n_649),
.B(n_641),
.C(n_548),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_694),
.B(n_669),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_699),
.A2(n_616),
.B(n_628),
.C(n_611),
.Y(n_701)
);

NOR3x1_ASAP7_75t_L g702 ( 
.A(n_698),
.B(n_611),
.C(n_664),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_697),
.B(n_670),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_703),
.Y(n_704)
);

NOR2x1_ASAP7_75t_L g705 ( 
.A(n_700),
.B(n_696),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_701),
.B(n_695),
.C(n_618),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_705),
.B(n_602),
.C(n_702),
.Y(n_707)
);

NOR2x1_ASAP7_75t_L g708 ( 
.A(n_704),
.B(n_618),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_SL g709 ( 
.A(n_706),
.B(n_590),
.C(n_641),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_704),
.Y(n_710)
);

NAND4xp75_ASAP7_75t_L g711 ( 
.A(n_708),
.B(n_710),
.C(n_707),
.D(n_709),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_707),
.A2(n_670),
.B1(n_674),
.B2(n_676),
.Y(n_712)
);

NAND4xp75_ASAP7_75t_L g713 ( 
.A(n_708),
.B(n_596),
.C(n_674),
.D(n_676),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_708),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_707),
.B(n_630),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_710),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_710),
.B(n_656),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_714),
.B(n_716),
.C(n_715),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_717),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_711),
.B(n_656),
.Y(n_720)
);

OR4x1_ASAP7_75t_L g721 ( 
.A(n_713),
.B(n_596),
.C(n_588),
.D(n_587),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_712),
.B(n_653),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_716),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_716),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_623),
.C(n_629),
.Y(n_725)
);

XNOR2xp5_ASAP7_75t_L g726 ( 
.A(n_719),
.B(n_623),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_720),
.A2(n_629),
.B1(n_626),
.B2(n_640),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_718),
.A2(n_654),
.B1(n_643),
.B2(n_626),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_723),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_725),
.A2(n_653),
.B1(n_629),
.B2(n_614),
.Y(n_730)
);

OA21x2_ASAP7_75t_L g731 ( 
.A1(n_724),
.A2(n_654),
.B(n_643),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_722),
.Y(n_732)
);

BUFx2_ASAP7_75t_SL g733 ( 
.A(n_721),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_732),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_733),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_726),
.A2(n_581),
.B1(n_570),
.B2(n_614),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_729),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_728),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_730),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_727),
.A2(n_592),
.B(n_593),
.Y(n_740)
);

OAI21x1_ASAP7_75t_SL g741 ( 
.A1(n_735),
.A2(n_731),
.B(n_593),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_734),
.B(n_592),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_738),
.A2(n_580),
.B1(n_566),
.B2(n_617),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_739),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_742),
.A2(n_737),
.B(n_740),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_736),
.B(n_481),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_581),
.B1(n_570),
.B2(n_580),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_745),
.A2(n_741),
.B(n_481),
.Y(n_748)
);

AO21x2_ASAP7_75t_L g749 ( 
.A1(n_746),
.A2(n_610),
.B(n_584),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_748),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_750),
.B(n_749),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_751),
.A2(n_747),
.B1(n_581),
.B2(n_570),
.Y(n_752)
);


endmodule