module fake_jpeg_5652_n_101 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_0),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_51),
.B1(n_43),
.B2(n_55),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_53),
.B(n_54),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_0),
.B(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_46),
.B1(n_45),
.B2(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_80),
.B(n_81),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_52),
.B(n_49),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_12),
.C(n_15),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_58),
.B(n_1),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_10),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_89),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_88),
.C(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_91),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_17),
.C(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_22),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_25),
.B(n_26),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_28),
.B(n_31),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_32),
.Y(n_101)
);


endmodule