module real_jpeg_5422_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_0),
.A2(n_189),
.B1(n_207),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_0),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_0),
.A2(n_101),
.B1(n_274),
.B2(n_355),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_0),
.A2(n_93),
.B1(n_274),
.B2(n_389),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g451 ( 
.A1(n_0),
.A2(n_139),
.B1(n_274),
.B2(n_452),
.Y(n_451)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_1),
.Y(n_240)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_1),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_1),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_2),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_2),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_2),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_2),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_3),
.A2(n_90),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_3),
.A2(n_90),
.B1(n_186),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_3),
.A2(n_90),
.B1(n_399),
.B2(n_402),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_4),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_4),
.A2(n_158),
.B1(n_188),
.B2(n_252),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_4),
.A2(n_188),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_4),
.A2(n_188),
.B1(n_344),
.B2(n_345),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_158),
.B1(n_159),
.B2(n_163),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_5),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_5),
.B(n_173),
.C(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_5),
.B(n_78),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_5),
.B(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_5),
.B(n_123),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_5),
.B(n_258),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_33),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_6),
.A2(n_51),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_6),
.A2(n_51),
.B1(n_375),
.B2(n_379),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_6),
.A2(n_51),
.B1(n_76),
.B2(n_392),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_7),
.A2(n_158),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_7),
.A2(n_184),
.B1(n_204),
.B2(n_212),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_7),
.A2(n_212),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_7),
.A2(n_143),
.B1(n_212),
.B2(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_9),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_10),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_13),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_13),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_14),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_14),
.A2(n_80),
.B1(n_95),
.B2(n_125),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_95),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_14),
.A2(n_95),
.B1(n_185),
.B2(n_370),
.Y(n_369)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_16),
.A2(n_55),
.B1(n_58),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_16),
.A2(n_61),
.B1(n_204),
.B2(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_16),
.A2(n_61),
.B1(n_214),
.B2(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_16),
.A2(n_61),
.B1(n_431),
.B2(n_436),
.Y(n_430)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_18),
.A2(n_126),
.B1(n_166),
.B2(n_169),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_18),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_18),
.A2(n_169),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_18),
.A2(n_169),
.B1(n_264),
.B2(n_267),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_18),
.A2(n_132),
.B1(n_169),
.B2(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_528),
.B(n_531),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_147),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_145),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_137),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_23),
.B(n_137),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_128),
.C(n_134),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_24),
.A2(n_25),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_62),
.C(n_96),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_26),
.B(n_516),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_27),
.A2(n_52),
.B1(n_54),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_27),
.A2(n_52),
.B1(n_129),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_27),
.A2(n_342),
.B(n_394),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_27),
.A2(n_38),
.B1(n_394),
.B2(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_27),
.A2(n_48),
.B1(n_52),
.B2(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_28),
.A2(n_339),
.B(n_341),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_28),
.B(n_343),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g317 ( 
.A1(n_33),
.A2(n_318),
.A3(n_319),
.B1(n_320),
.B2(n_322),
.Y(n_317)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_35),
.Y(n_139)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_36),
.Y(n_319)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_37),
.Y(n_321)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_38),
.B(n_163),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_38)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_40),
.Y(n_351)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_42),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_42),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_42),
.Y(n_435)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_43),
.Y(n_261)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_43),
.Y(n_269)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g277 ( 
.A(n_45),
.Y(n_277)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_49),
.Y(n_419)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_50),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_52),
.A2(n_417),
.B(n_455),
.Y(n_465)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_53),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_53),
.B(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_62),
.A2(n_96),
.B1(n_97),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_62),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_63),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_63),
.A2(n_91),
.B1(n_290),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_63),
.A2(n_91),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_63),
.A2(n_86),
.B1(n_91),
.B2(n_505),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_75),
.B(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g255 ( 
.A1(n_76),
.A2(n_163),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_77),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_78),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_78),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_78),
.A2(n_135),
.B1(n_297),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_78),
.A2(n_135),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_78)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_80),
.Y(n_385)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_81),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_83),
.Y(n_355)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_83),
.Y(n_381)
);

AOI32xp33_ASAP7_75t_L g276 ( 
.A1(n_84),
.A2(n_158),
.A3(n_257),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_85),
.Y(n_279)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_91),
.B(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_91),
.A2(n_290),
.B(n_296),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_96),
.A2(n_97),
.B1(n_503),
.B2(n_504),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_96),
.B(n_500),
.C(n_503),
.Y(n_511)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_122),
.B(n_124),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_98),
.A2(n_157),
.B(n_164),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_98),
.A2(n_122),
.B1(n_211),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_98),
.A2(n_164),
.B(n_251),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_98),
.A2(n_122),
.B1(n_354),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_99),
.B(n_165),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_99),
.A2(n_123),
.B1(n_374),
.B2(n_382),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_99),
.A2(n_123),
.B1(n_382),
.B2(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_99),
.A2(n_123),
.B1(n_398),
.B2(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_110),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_111),
.Y(n_403)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_112),
.A2(n_211),
.B(n_215),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_119),
.B2(n_121),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_120),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_122),
.A2(n_215),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_124),
.Y(n_442)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_128),
.B(n_134),
.Y(n_525)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_135),
.A2(n_255),
.B(n_262),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_135),
.B(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_135),
.A2(n_262),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_522),
.B(n_527),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_494),
.B(n_519),
.Y(n_148)
);

OAI311xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_358),
.A3(n_470),
.B1(n_488),
.C1(n_489),
.Y(n_149)
);

AOI21x1_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_311),
.B(n_357),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_281),
.B(n_310),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_245),
.B(n_280),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_218),
.B(n_244),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_181),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_155),
.B(n_181),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_170),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_156),
.A2(n_170),
.B1(n_171),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_156),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_162),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_163),
.A2(n_193),
.B(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_163),
.B(n_323),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g339 ( 
.A1(n_163),
.A2(n_322),
.B(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_167),
.Y(n_252)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_208),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_182),
.B(n_209),
.C(n_217),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_193),
.B(n_200),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_193),
.A2(n_275),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_193),
.A2(n_364),
.B1(n_367),
.B2(n_369),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_193),
.A2(n_369),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_203),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_194),
.A2(n_273),
.B1(n_301),
.B2(n_306),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_194),
.A2(n_330),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_196),
.Y(n_405)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_202),
.Y(n_368)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_206),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_216),
.B2(n_217),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_213),
.B(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_235),
.B(n_243),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_228),
.B(n_234),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_233),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_241),
.Y(n_243)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_247),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_270),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_253),
.C(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_261),
.Y(n_439)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_266),
.Y(n_390)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_282),
.B(n_283),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_309),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_287),
.C(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_298),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_299),
.C(n_300),
.Y(n_333)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_291),
.Y(n_352)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_312),
.B(n_313),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_336),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_314)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_315),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_326),
.B2(n_327),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_317),
.B(n_326),
.Y(n_466)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_333),
.B(n_334),
.C(n_336),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_347),
.B2(n_356),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_337),
.B(n_348),
.C(n_353),
.Y(n_479)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_349),
.Y(n_468)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_456),
.Y(n_358)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_359),
.A2(n_456),
.B(n_490),
.C(n_493),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_422),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_360),
.B(n_422),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_395),
.C(n_407),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_361),
.B(n_395),
.CI(n_407),
.CON(n_469),
.SN(n_469)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_386),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_387),
.C(n_393),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_373),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_363),
.B(n_373),
.Y(n_462)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_393),
.Y(n_386)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_404),
.B2(n_406),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_404),
.Y(n_446)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_404),
.A2(n_406),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_404),
.A2(n_446),
.B(n_449),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_415),
.C(n_420),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_409),
.B(n_411),
.Y(n_478)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_415),
.A2(n_416),
.B1(n_420),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_426),
.C(n_444),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_444),
.B2(n_445),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_440),
.B(n_443),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_441),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

FAx1_ASAP7_75t_SL g496 ( 
.A(n_443),
.B(n_497),
.CI(n_498),
.CON(n_496),
.SN(n_496)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_497),
.C(n_498),
.Y(n_518)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_455),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx8_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_469),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_469),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_462),
.C(n_463),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_458),
.A2(n_459),
.B1(n_462),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.C(n_467),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_467),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_469),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_483),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_472),
.A2(n_491),
.B(n_492),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_480),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_480),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.C(n_479),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_486),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_478),
.B1(n_479),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_479),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_484),
.B(n_485),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_508),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_507),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_507),
.Y(n_520)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_496),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_500),
.B1(n_502),
.B2(n_506),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_499),
.A2(n_500),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_510),
.C(n_514),
.Y(n_526)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_502),
.Y(n_506)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_508),
.A2(n_520),
.B(n_521),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_518),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_518),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_526),
.Y(n_527)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx13_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_530),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_534),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);


endmodule