module fake_ibex_493_n_1017 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1017);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1017;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_375;
wire n_340;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_262;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_597;
wire n_415;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_885;
wire n_588;
wire n_212;
wire n_513;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_890;
wire n_874;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_988;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_947;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_1),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_92),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_68),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_34),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_71),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_64),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_116),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_108),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_109),
.B(n_198),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_87),
.B(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_18),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_102),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_23),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_34),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_25),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_2),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_104),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_119),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_66),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_80),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_133),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_60),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_126),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_146),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_179),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_149),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_74),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_132),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_75),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_129),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_51),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_137),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_59),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_163),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_117),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_185),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_19),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_107),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_0),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_120),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_125),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_44),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_91),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_147),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_85),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_52),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_12),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_189),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_57),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_69),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_90),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_58),
.B(n_30),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_49),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_139),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_142),
.B(n_177),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_33),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_128),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_22),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_32),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_100),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_159),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_32),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_86),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_39),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_101),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_93),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_167),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_45),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_38),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_25),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_115),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_98),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_118),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_36),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_78),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_6),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_178),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_76),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_195),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_0),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_193),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_175),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_141),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_36),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_144),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_38),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_134),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_215),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_213),
.B(n_255),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_222),
.A2(n_275),
.B1(n_295),
.B2(n_229),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_257),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_202),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_211),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_211),
.B(n_3),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_202),
.B(n_4),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_213),
.B(n_7),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_8),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_9),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_285),
.B(n_9),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_269),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_201),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_211),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_201),
.Y(n_347)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_233),
.A2(n_84),
.B(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_209),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_220),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_247),
.B(n_260),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_216),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_224),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_247),
.B(n_14),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_230),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_260),
.B(n_15),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_300),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_L g364 ( 
.A(n_210),
.B(n_53),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_256),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_243),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_269),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_270),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_280),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_243),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_219),
.B(n_16),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_282),
.B(n_16),
.Y(n_377)
);

BUFx8_ASAP7_75t_L g378 ( 
.A(n_200),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g380 ( 
.A1(n_316),
.A2(n_103),
.B(n_188),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_306),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_219),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_225),
.B(n_17),
.Y(n_383)
);

OAI22x1_ASAP7_75t_SL g384 ( 
.A1(n_222),
.A2(n_229),
.B1(n_295),
.B2(n_275),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_225),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_220),
.Y(n_386)
);

OR2x6_ASAP7_75t_L g387 ( 
.A(n_288),
.B(n_17),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_248),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_287),
.B(n_18),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_287),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_293),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_304),
.B(n_20),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_304),
.B(n_20),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_269),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_299),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_248),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_314),
.B(n_21),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_252),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_305),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_21),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_207),
.C(n_206),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_402),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_280),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_360),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

BUFx4f_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_329),
.B(n_210),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_208),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_214),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_377),
.A2(n_323),
.B1(n_250),
.B2(n_267),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_364),
.B(n_212),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_387),
.B(n_204),
.Y(n_427)
);

NOR2x1p5_ASAP7_75t_L g428 ( 
.A(n_381),
.B(n_214),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_221),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_343),
.B(n_226),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_327),
.B(n_223),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_346),
.B(n_351),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_347),
.B(n_382),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_228),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_359),
.B(n_372),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_377),
.B(n_252),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_400),
.A2(n_249),
.B1(n_308),
.B2(n_232),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_372),
.B(n_223),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_235),
.C(n_234),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_328),
.B(n_292),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_382),
.B(n_236),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_385),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_292),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_331),
.B(n_296),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_391),
.B(n_296),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_380),
.B(n_237),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_334),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_350),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_330),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_348),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g466 ( 
.A1(n_387),
.A2(n_307),
.B1(n_305),
.B2(n_277),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_336),
.B(n_302),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_334),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_374),
.B(n_302),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_340),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_340),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_340),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_340),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_338),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_339),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_342),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_342),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_383),
.B(n_326),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_341),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_349),
.A2(n_244),
.B(n_239),
.Y(n_482)
);

BUFx4f_ASAP7_75t_L g483 ( 
.A(n_352),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_354),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_354),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_353),
.B(n_366),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_339),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_367),
.B(n_205),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_356),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_356),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_356),
.Y(n_491)
);

NOR2x1p5_ASAP7_75t_L g492 ( 
.A(n_378),
.B(n_245),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_384),
.B(n_307),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_356),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_358),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_358),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_358),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_358),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_389),
.B(n_279),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_361),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_361),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_361),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_392),
.B(n_395),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_357),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_361),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_362),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_397),
.B(n_231),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_362),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_362),
.Y(n_509)
);

AOI221xp5_ASAP7_75t_L g510 ( 
.A1(n_433),
.A2(n_399),
.B1(n_332),
.B2(n_393),
.C(n_390),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_394),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_419),
.A2(n_337),
.B1(n_378),
.B2(n_344),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_419),
.A2(n_277),
.B1(n_204),
.B2(n_227),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

NOR2x1p5_ASAP7_75t_L g516 ( 
.A(n_454),
.B(n_457),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_462),
.B(n_435),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_479),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_419),
.B(n_238),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_427),
.A2(n_355),
.B1(n_227),
.B2(n_241),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_453),
.B(n_376),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_483),
.B(n_240),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_241),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_480),
.B(n_251),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_427),
.A2(n_283),
.B1(n_271),
.B2(n_273),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_483),
.B(n_258),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_410),
.B(n_246),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_412),
.A2(n_289),
.B1(n_259),
.B2(n_261),
.Y(n_528)
);

O2A1O1Ixp5_ASAP7_75t_L g529 ( 
.A1(n_450),
.A2(n_290),
.B(n_278),
.C(n_284),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_416),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_416),
.A2(n_301),
.B(n_309),
.C(n_294),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_412),
.A2(n_274),
.B1(n_315),
.B2(n_303),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_22),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_483),
.B(n_426),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_404),
.Y(n_537)
);

O2A1O1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_441),
.A2(n_322),
.B(n_313),
.C(n_311),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_480),
.B(n_203),
.Y(n_539)
);

NOR2x1p5_ASAP7_75t_L g540 ( 
.A(n_432),
.B(n_253),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_458),
.A2(n_217),
.B(n_218),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_411),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_467),
.B(n_475),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_410),
.B(n_467),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_442),
.A2(n_321),
.B1(n_272),
.B2(n_242),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_430),
.B(n_254),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_426),
.B(n_262),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_426),
.B(n_268),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_408),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_492),
.B(n_281),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_406),
.B(n_276),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_406),
.B(n_286),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_428),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_442),
.A2(n_324),
.B1(n_310),
.B2(n_368),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_404),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_470),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_436),
.B(n_363),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_420),
.B(n_363),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_420),
.B(n_499),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_417),
.Y(n_562)
);

AND2x6_ASAP7_75t_SL g563 ( 
.A(n_493),
.B(n_23),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_409),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_488),
.B(n_368),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_458),
.A2(n_373),
.B(n_370),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_423),
.A2(n_373),
.B1(n_370),
.B2(n_27),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_486),
.B(n_370),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_417),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_446),
.B(n_373),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_422),
.B(n_373),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_503),
.B(n_24),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_452),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_442),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_458),
.B(n_54),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_418),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_470),
.B(n_26),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_487),
.B(n_55),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_455),
.Y(n_580)
);

AND2x2_ASAP7_75t_SL g581 ( 
.A(n_464),
.B(n_29),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_507),
.B(n_56),
.Y(n_582)
);

AND2x4_ASAP7_75t_SL g583 ( 
.A(n_476),
.B(n_29),
.Y(n_583)
);

BUFx8_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

AO221x1_ASAP7_75t_L g585 ( 
.A1(n_466),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.C(n_35),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_451),
.B(n_31),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_493),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_442),
.A2(n_405),
.B1(n_447),
.B2(n_482),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_421),
.B(n_61),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_407),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_476),
.B(n_62),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_449),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_444),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_481),
.B(n_41),
.C(n_42),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_429),
.B(n_63),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_481),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_450),
.B(n_479),
.Y(n_600)
);

AOI33xp33_ASAP7_75t_L g601 ( 
.A1(n_543),
.A2(n_459),
.A3(n_438),
.B1(n_434),
.B2(n_425),
.B3(n_463),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_517),
.B(n_476),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_566),
.A2(n_450),
.B(n_479),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_524),
.A2(n_438),
.B(n_434),
.C(n_425),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_523),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_518),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_515),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g608 ( 
.A(n_550),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_593),
.Y(n_609)
);

AO32x1_ASAP7_75t_L g610 ( 
.A1(n_596),
.A2(n_450),
.A3(n_567),
.B1(n_583),
.B2(n_515),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_599),
.Y(n_611)
);

O2A1O1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_561),
.A2(n_456),
.B(n_448),
.C(n_459),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_593),
.B(n_469),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_544),
.B(n_449),
.Y(n_614)
);

OAI22x1_ASAP7_75t_L g615 ( 
.A1(n_525),
.A2(n_492),
.B1(n_445),
.B2(n_46),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_516),
.B(n_540),
.Y(n_616)
);

BUFx2_ASAP7_75t_SL g617 ( 
.A(n_578),
.Y(n_617)
);

OA22x2_ASAP7_75t_L g618 ( 
.A1(n_521),
.A2(n_588),
.B1(n_585),
.B2(n_583),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_531),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_539),
.B(n_445),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_581),
.A2(n_413),
.B1(n_414),
.B2(n_460),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_511),
.B(n_43),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_524),
.B(n_45),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_539),
.B(n_46),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_589),
.A2(n_431),
.B1(n_437),
.B2(n_443),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_532),
.A2(n_439),
.B(n_440),
.C(n_443),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_518),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_R g628 ( 
.A(n_584),
.B(n_47),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_584),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_595),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_584),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_513),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_536),
.A2(n_559),
.B(n_526),
.Y(n_633)
);

INVx6_ASAP7_75t_L g634 ( 
.A(n_551),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_514),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_576),
.A2(n_509),
.B(n_477),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_526),
.A2(n_545),
.B(n_537),
.Y(n_637)
);

AND2x6_ASAP7_75t_SL g638 ( 
.A(n_551),
.B(n_48),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_554),
.B(n_48),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_556),
.A2(n_560),
.B(n_565),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_520),
.A2(n_501),
.B1(n_494),
.B2(n_505),
.C(n_502),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_573),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

O2A1O1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_587),
.A2(n_501),
.B(n_491),
.C(n_505),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_574),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_580),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_512),
.A2(n_485),
.B1(n_502),
.B2(n_500),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_L g648 ( 
.A1(n_572),
.A2(n_50),
.B1(n_484),
.B2(n_474),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_597),
.A2(n_474),
.B1(n_485),
.B2(n_500),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_546),
.B(n_484),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_579),
.B(n_484),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_551),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_580),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_530),
.A2(n_489),
.B(n_506),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_557),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_548),
.A2(n_549),
.B(n_527),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_575),
.A2(n_508),
.B1(n_498),
.B2(n_497),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_547),
.B(n_528),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_SL g659 ( 
.A(n_535),
.B(n_461),
.Y(n_659)
);

AOI21x1_ASAP7_75t_L g660 ( 
.A1(n_594),
.A2(n_496),
.B(n_495),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_547),
.B(n_65),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_591),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_577),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_533),
.B(n_67),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_586),
.B(n_564),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_552),
.A2(n_478),
.B(n_471),
.Y(n_666)
);

O2A1O1Ixp5_ASAP7_75t_L g667 ( 
.A1(n_529),
.A2(n_478),
.B(n_471),
.C(n_468),
.Y(n_667)
);

CKINVDCx11_ASAP7_75t_R g668 ( 
.A(n_563),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_538),
.B(n_519),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_571),
.A2(n_490),
.B(n_473),
.Y(n_670)
);

OAI21xp33_ASAP7_75t_L g671 ( 
.A1(n_541),
.A2(n_490),
.B(n_473),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_522),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_562),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_562),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_568),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_558),
.A2(n_472),
.B(n_415),
.Y(n_676)
);

OAI21xp33_ASAP7_75t_L g677 ( 
.A1(n_555),
.A2(n_415),
.B(n_73),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_534),
.A2(n_569),
.B(n_582),
.C(n_542),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_558),
.A2(n_415),
.B(n_77),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_582),
.B(n_72),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_611),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_653),
.B(n_570),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_624),
.A2(n_590),
.B(n_598),
.C(n_570),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_602),
.A2(n_620),
.B(n_656),
.C(n_601),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_608),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_629),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_643),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_634),
.Y(n_688)
);

O2A1O1Ixp5_ASAP7_75t_L g689 ( 
.A1(n_651),
.A2(n_592),
.B(n_81),
.C(n_82),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_678),
.A2(n_619),
.B(n_607),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_645),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_605),
.B(n_592),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_617),
.A2(n_79),
.B1(n_83),
.B2(n_94),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_605),
.B(n_96),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_614),
.A2(n_99),
.B(n_105),
.C(n_106),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_606),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_652),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_658),
.A2(n_110),
.B(n_111),
.C(n_112),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_636),
.A2(n_113),
.B(n_114),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_616),
.B(n_121),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_668),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_616),
.B(n_122),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_633),
.A2(n_123),
.B(n_124),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_665),
.A2(n_640),
.B(n_637),
.Y(n_704)
);

CKINVDCx8_ASAP7_75t_R g705 ( 
.A(n_638),
.Y(n_705)
);

AO31x2_ASAP7_75t_L g706 ( 
.A1(n_604),
.A2(n_136),
.A3(n_138),
.B(n_140),
.Y(n_706)
);

INVx8_ASAP7_75t_L g707 ( 
.A(n_652),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_625),
.A2(n_145),
.A3(n_148),
.B(n_150),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_623),
.A2(n_151),
.B(n_152),
.C(n_154),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_660),
.A2(n_158),
.B(n_160),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_645),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_627),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_641),
.B(n_649),
.C(n_621),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_631),
.B(n_162),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_628),
.Y(n_715)
);

AO32x2_ASAP7_75t_L g716 ( 
.A1(n_657),
.A2(n_164),
.A3(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_615),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_612),
.A2(n_170),
.B(n_171),
.C(n_172),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_L g719 ( 
.A1(n_618),
.A2(n_669),
.B1(n_639),
.B2(n_672),
.C(n_622),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_676),
.A2(n_182),
.B(n_183),
.Y(n_720)
);

AO31x2_ASAP7_75t_L g721 ( 
.A1(n_679),
.A2(n_184),
.A3(n_187),
.B(n_670),
.Y(n_721)
);

BUFx4f_ASAP7_75t_L g722 ( 
.A(n_638),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_642),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_632),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_646),
.B(n_662),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_626),
.A2(n_675),
.B(n_680),
.C(n_659),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_647),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_680),
.A2(n_644),
.B(n_671),
.C(n_677),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_655),
.B(n_673),
.Y(n_729)
);

CKINVDCx16_ASAP7_75t_R g730 ( 
.A(n_627),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_630),
.A2(n_657),
.B1(n_613),
.B2(n_650),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_648),
.A2(n_630),
.B1(n_664),
.B2(n_609),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_666),
.A2(n_667),
.B(n_609),
.C(n_654),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_674),
.B(n_610),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_663),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_603),
.A2(n_600),
.B(n_602),
.Y(n_736)
);

AND2x6_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_617),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_635),
.B(n_521),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_635),
.B(n_521),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_602),
.B(n_517),
.Y(n_740)
);

AO31x2_ASAP7_75t_L g741 ( 
.A1(n_604),
.A2(n_450),
.A3(n_465),
.B(n_566),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_608),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_602),
.B(n_517),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_629),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_603),
.A2(n_566),
.B(n_636),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_602),
.B(n_517),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_603),
.A2(n_600),
.B(n_602),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_608),
.Y(n_748)
);

NAND2x1p5_ASAP7_75t_L g749 ( 
.A(n_629),
.B(n_419),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_624),
.A2(n_602),
.B(n_620),
.C(n_656),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_643),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_602),
.B(n_517),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_603),
.A2(n_566),
.B(n_636),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_603),
.A2(n_600),
.B(n_602),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_603),
.A2(n_600),
.B(n_602),
.Y(n_755)
);

AO31x2_ASAP7_75t_L g756 ( 
.A1(n_604),
.A2(n_450),
.A3(n_465),
.B(n_566),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_603),
.A2(n_600),
.B(n_602),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_608),
.Y(n_758)
);

AOI221x1_ASAP7_75t_L g759 ( 
.A1(n_671),
.A2(n_541),
.B1(n_677),
.B2(n_657),
.C(n_597),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_602),
.B(n_517),
.Y(n_760)
);

AOI21xp33_ASAP7_75t_L g761 ( 
.A1(n_602),
.A2(n_487),
.B(n_481),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_633),
.A2(n_600),
.B(n_529),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_602),
.B(n_616),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_611),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_602),
.A2(n_523),
.B1(n_427),
.B2(n_521),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_611),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_602),
.B(n_517),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_SL g768 ( 
.A1(n_661),
.A2(n_576),
.B(n_604),
.C(n_651),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_663),
.Y(n_769)
);

AO31x2_ASAP7_75t_L g770 ( 
.A1(n_604),
.A2(n_450),
.A3(n_465),
.B(n_566),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_602),
.A2(n_523),
.B1(n_427),
.B2(n_521),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_611),
.B(n_402),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_602),
.B(n_616),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_603),
.A2(n_566),
.B(n_636),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_602),
.B(n_427),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_603),
.A2(n_600),
.B(n_602),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_602),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_602),
.B(n_517),
.Y(n_778)
);

NAND3xp33_ASAP7_75t_L g779 ( 
.A(n_624),
.B(n_541),
.C(n_510),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_740),
.B(n_743),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_724),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_738),
.A2(n_739),
.B1(n_717),
.B2(n_746),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_711),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_711),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_752),
.B(n_760),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_767),
.B(n_778),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_735),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_772),
.B(n_681),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_684),
.A2(n_754),
.B(n_757),
.Y(n_789)
);

BUFx2_ASAP7_75t_R g790 ( 
.A(n_748),
.Y(n_790)
);

AND2x2_ASAP7_75t_SL g791 ( 
.A(n_722),
.B(n_730),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_734),
.A2(n_759),
.B(n_745),
.Y(n_792)
);

NOR2x1_ASAP7_75t_SL g793 ( 
.A(n_711),
.B(n_712),
.Y(n_793)
);

AO21x2_ASAP7_75t_L g794 ( 
.A1(n_726),
.A2(n_753),
.B(n_774),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_742),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_777),
.B(n_779),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_742),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_736),
.A2(n_776),
.B(n_747),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_765),
.B(n_771),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_768),
.A2(n_704),
.B(n_733),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_719),
.B(n_775),
.C(n_750),
.Y(n_801)
);

INVx8_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_769),
.Y(n_803)
);

OA21x2_ASAP7_75t_L g804 ( 
.A1(n_710),
.A2(n_699),
.B(n_703),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_764),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_755),
.A2(n_690),
.B(n_762),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_715),
.A2(n_744),
.B1(n_705),
.B2(n_701),
.Y(n_807)
);

OA21x2_ASAP7_75t_L g808 ( 
.A1(n_720),
.A2(n_718),
.B(n_689),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_713),
.A2(n_727),
.B(n_683),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_707),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_712),
.B(n_723),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_766),
.B(n_773),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_761),
.A2(n_732),
.B(n_731),
.C(n_694),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_763),
.B(n_714),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_686),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_763),
.B(n_725),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_729),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_692),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_749),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_696),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_737),
.B(n_751),
.Y(n_821)
);

AO31x2_ASAP7_75t_L g822 ( 
.A1(n_698),
.A2(n_709),
.A3(n_695),
.B(n_693),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_687),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_682),
.A2(n_691),
.B(n_700),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_741),
.B(n_770),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_707),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_697),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_702),
.Y(n_828)
);

BUFx8_ASAP7_75t_L g829 ( 
.A(n_688),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_685),
.B(n_758),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_682),
.A2(n_716),
.B1(n_756),
.B2(n_721),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_682),
.B(n_721),
.Y(n_832)
);

AO21x2_ASAP7_75t_L g833 ( 
.A1(n_708),
.A2(n_716),
.B(n_706),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_716),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_721),
.B(n_711),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_711),
.B(n_740),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_738),
.B(n_523),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_711),
.B(n_740),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_740),
.B(n_743),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_724),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_SL g841 ( 
.A1(n_693),
.A2(n_777),
.B(n_728),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_707),
.B(n_617),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_779),
.B(n_624),
.C(n_597),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_684),
.A2(n_747),
.B(n_736),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_724),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_684),
.A2(n_747),
.B(n_736),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_740),
.A2(n_743),
.B(n_752),
.C(n_746),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_738),
.A2(n_618),
.B1(n_581),
.B2(n_739),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_740),
.B(n_743),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_711),
.B(n_427),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_724),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_711),
.B(n_427),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_796),
.Y(n_853)
);

CKINVDCx6p67_ASAP7_75t_R g854 ( 
.A(n_795),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_802),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_817),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_835),
.B(n_824),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_805),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_799),
.B(n_780),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_780),
.B(n_785),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_847),
.A2(n_843),
.B(n_813),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_781),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_840),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_799),
.B(n_785),
.Y(n_864)
);

OAI21x1_ASAP7_75t_L g865 ( 
.A1(n_800),
.A2(n_806),
.B(n_798),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_845),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_783),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_837),
.B(n_788),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_851),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_818),
.Y(n_870)
);

OAI21x1_ASAP7_75t_SL g871 ( 
.A1(n_793),
.A2(n_824),
.B(n_832),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_786),
.B(n_839),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_802),
.B(n_841),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_849),
.B(n_782),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_849),
.B(n_809),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_809),
.B(n_787),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_783),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_816),
.B(n_825),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_848),
.B(n_812),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_798),
.A2(n_831),
.B(n_846),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_835),
.B(n_842),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_842),
.B(n_811),
.Y(n_882)
);

AO21x2_ASAP7_75t_L g883 ( 
.A1(n_789),
.A2(n_844),
.B(n_846),
.Y(n_883)
);

INVx3_ASAP7_75t_SL g884 ( 
.A(n_842),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_803),
.B(n_836),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_834),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_838),
.B(n_816),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_801),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_815),
.B(n_828),
.Y(n_889)
);

OAI332xp33_ASAP7_75t_L g890 ( 
.A1(n_826),
.A2(n_850),
.A3(n_852),
.B1(n_823),
.B2(n_821),
.B3(n_807),
.C1(n_790),
.C2(n_791),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_819),
.B(n_814),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_811),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_784),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_784),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_830),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_833),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_797),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_830),
.B(n_810),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_829),
.B(n_820),
.Y(n_899)
);

BUFx2_ASAP7_75t_SL g900 ( 
.A(n_855),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_878),
.B(n_792),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_860),
.B(n_792),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_881),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_890),
.B(n_861),
.C(n_874),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_878),
.B(n_794),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_872),
.B(n_827),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_875),
.B(n_822),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_882),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_857),
.B(n_887),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_853),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_887),
.B(n_822),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_857),
.B(n_804),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_876),
.B(n_808),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_876),
.B(n_790),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_896),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_857),
.B(n_829),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_856),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_868),
.A2(n_879),
.B1(n_864),
.B2(n_859),
.Y(n_919)
);

NOR2x1_ASAP7_75t_L g920 ( 
.A(n_881),
.B(n_882),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_885),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_883),
.B(n_880),
.Y(n_922)
);

AND2x4_ASAP7_75t_SL g923 ( 
.A(n_881),
.B(n_882),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_883),
.B(n_880),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_873),
.B(n_883),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_892),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_880),
.B(n_870),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_926),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_902),
.B(n_880),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_912),
.B(n_886),
.Y(n_931)
);

NAND2x1_ASAP7_75t_L g932 ( 
.A(n_910),
.B(n_871),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_912),
.B(n_886),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_911),
.B(n_888),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_922),
.B(n_924),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_908),
.B(n_927),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_923),
.B(n_855),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_913),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_927),
.B(n_922),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_901),
.B(n_865),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_936),
.B(n_918),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_935),
.B(n_901),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_935),
.B(n_905),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_905),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_936),
.B(n_907),
.Y(n_945)
);

AND2x4_ASAP7_75t_SL g946 ( 
.A(n_937),
.B(n_917),
.Y(n_946)
);

OAI31xp33_ASAP7_75t_L g947 ( 
.A1(n_928),
.A2(n_904),
.A3(n_917),
.B(n_915),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_929),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_939),
.B(n_919),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_934),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_939),
.B(n_914),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_931),
.B(n_921),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_929),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_928),
.Y(n_954)
);

AND2x4_ASAP7_75t_SL g955 ( 
.A(n_937),
.B(n_917),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_930),
.B(n_914),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_930),
.B(n_925),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_930),
.B(n_925),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_942),
.B(n_940),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_950),
.B(n_931),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_948),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_956),
.B(n_938),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_945),
.B(n_854),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_948),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_956),
.B(n_938),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_949),
.B(n_933),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_953),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_953),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_954),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_942),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_969),
.A2(n_947),
.B(n_904),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_970),
.A2(n_955),
.B1(n_946),
.B2(n_941),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_962),
.B(n_957),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_961),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_963),
.A2(n_906),
.B(n_915),
.Y(n_975)
);

OAI21xp33_ASAP7_75t_L g976 ( 
.A1(n_959),
.A2(n_958),
.B(n_957),
.Y(n_976)
);

AOI322xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_952),
.A3(n_951),
.B1(n_958),
.B2(n_917),
.C1(n_937),
.C2(n_920),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_959),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_961),
.Y(n_979)
);

NOR2xp67_ASAP7_75t_L g980 ( 
.A(n_962),
.B(n_909),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_968),
.Y(n_981)
);

XNOR2xp5_ASAP7_75t_L g982 ( 
.A(n_966),
.B(n_946),
.Y(n_982)
);

OAI221xp5_ASAP7_75t_L g983 ( 
.A1(n_971),
.A2(n_960),
.B1(n_932),
.B2(n_943),
.C(n_944),
.Y(n_983)
);

OAI221xp5_ASAP7_75t_L g984 ( 
.A1(n_977),
.A2(n_932),
.B1(n_943),
.B2(n_944),
.C(n_964),
.Y(n_984)
);

OAI211xp5_ASAP7_75t_SL g985 ( 
.A1(n_975),
.A2(n_899),
.B(n_920),
.C(n_889),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_976),
.A2(n_955),
.B(n_965),
.C(n_923),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_978),
.A2(n_965),
.B1(n_938),
.B2(n_951),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_SL g988 ( 
.A1(n_978),
.A2(n_923),
.B1(n_909),
.B2(n_900),
.Y(n_988)
);

AOI222xp33_ASAP7_75t_L g989 ( 
.A1(n_984),
.A2(n_982),
.B1(n_981),
.B2(n_980),
.C1(n_973),
.C2(n_967),
.Y(n_989)
);

OAI211xp5_ASAP7_75t_L g990 ( 
.A1(n_983),
.A2(n_972),
.B(n_897),
.C(n_898),
.Y(n_990)
);

AOI211xp5_ASAP7_75t_L g991 ( 
.A1(n_985),
.A2(n_890),
.B(n_982),
.C(n_884),
.Y(n_991)
);

NAND4xp25_ASAP7_75t_L g992 ( 
.A(n_989),
.B(n_986),
.C(n_988),
.D(n_897),
.Y(n_992)
);

NAND4xp25_ASAP7_75t_L g993 ( 
.A(n_991),
.B(n_987),
.C(n_855),
.D(n_903),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_992),
.B(n_990),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_L g995 ( 
.A(n_993),
.B(n_895),
.C(n_893),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_994),
.A2(n_854),
.B1(n_973),
.B2(n_873),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_995),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_997),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_996),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_998),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_999),
.B(n_974),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_998),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_1000),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_1002),
.A2(n_884),
.B1(n_909),
.B2(n_900),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_1001),
.A2(n_884),
.B1(n_882),
.B2(n_873),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_1000),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_1006),
.A2(n_882),
.B(n_891),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_974),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_1004),
.B(n_979),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_1005),
.A2(n_894),
.B(n_877),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_1006),
.A2(n_867),
.B(n_873),
.Y(n_1011)
);

AOI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_1006),
.A2(n_869),
.B(n_862),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_862),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_1011),
.A2(n_869),
.B(n_863),
.Y(n_1014)
);

AO21x2_ASAP7_75t_L g1015 ( 
.A1(n_1008),
.A2(n_863),
.B(n_866),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_1013),
.A2(n_1010),
.B(n_1009),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_1016),
.A2(n_1015),
.B1(n_1014),
.B2(n_1012),
.Y(n_1017)
);


endmodule