module fake_jpeg_8557_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_4),
.B(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_2),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_14),
.C(n_12),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_16),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_36),
.B1(n_13),
.B2(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_13),
.B1(n_8),
.B2(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.C(n_34),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_30),
.B1(n_33),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_42),
.B1(n_30),
.B2(n_25),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_26),
.C(n_38),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_51),
.B(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_26),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_47),
.C(n_26),
.Y(n_54)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_10),
.B(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_53),
.B1(n_10),
.B2(n_4),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_6),
.C(n_7),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_2),
.B(n_3),
.Y(n_58)
);


endmodule