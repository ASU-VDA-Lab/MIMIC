module real_aes_4593_n_391 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_1331, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_1330, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_391);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_1331;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_1330;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_391;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_905;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g879 ( .A(n_0), .Y(n_879) );
INVx1_ASAP7_75t_L g949 ( .A(n_1), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_2), .A2(n_377), .B1(n_523), .B2(n_733), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_3), .A2(n_232), .B1(n_598), .B2(n_634), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_4), .A2(n_313), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_5), .A2(n_375), .B1(n_561), .B2(n_681), .Y(n_687) );
AOI21xp33_ASAP7_75t_SL g756 ( .A1(n_6), .A2(n_569), .B(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_7), .A2(n_201), .B1(n_658), .B2(n_659), .Y(n_657) );
AO22x1_ASAP7_75t_L g698 ( .A1(n_8), .A2(n_237), .B1(n_664), .B2(n_665), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_9), .A2(n_284), .B1(n_530), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_10), .A2(n_170), .B1(n_744), .B2(n_745), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_11), .A2(n_319), .B1(n_467), .B2(n_523), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_12), .A2(n_205), .B1(n_561), .B2(n_673), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_13), .A2(n_24), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_14), .A2(n_38), .B1(n_519), .B2(n_545), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_15), .A2(n_357), .B1(n_528), .B2(n_774), .Y(n_773) );
AOI21xp33_ASAP7_75t_SL g1057 ( .A1(n_16), .A2(n_886), .B(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g887 ( .A(n_17), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_18), .A2(n_208), .B1(n_614), .B2(n_616), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_19), .B(n_421), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_20), .A2(n_177), .B1(n_821), .B2(n_822), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_21), .A2(n_191), .B1(n_494), .B2(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_22), .A2(n_346), .B1(n_1099), .B2(n_1105), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_23), .A2(n_354), .B1(n_518), .B2(n_598), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_25), .A2(n_307), .B1(n_467), .B2(n_523), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_26), .A2(n_299), .B1(n_726), .B2(n_742), .C(n_818), .Y(n_817) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_27), .Y(n_421) );
INVx1_ASAP7_75t_L g942 ( .A(n_28), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_29), .A2(n_74), .B1(n_916), .B2(n_1300), .Y(n_1299) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_30), .A2(n_89), .B1(n_658), .B2(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_31), .A2(n_376), .B1(n_460), .B2(n_463), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_32), .A2(n_44), .B1(n_569), .B2(n_571), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_33), .A2(n_901), .B(n_902), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_34), .A2(n_36), .B1(n_445), .B2(n_769), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_35), .A2(n_152), .B1(n_600), .B2(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_37), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_39), .B(n_563), .Y(n_562) );
AO22x2_ASAP7_75t_L g870 ( .A1(n_40), .A2(n_871), .B1(n_876), .B2(n_896), .Y(n_870) );
INVxp33_ASAP7_75t_SL g895 ( .A(n_40), .Y(n_895) );
INVx1_ASAP7_75t_L g504 ( .A(n_41), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_42), .A2(n_215), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_43), .A2(n_125), .B1(n_550), .B2(n_632), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_45), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_46), .A2(n_155), .B1(n_523), .B2(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_47), .A2(n_209), .B1(n_632), .B2(n_828), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_48), .A2(n_371), .B1(n_546), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g807 ( .A(n_49), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_50), .A2(n_102), .B1(n_415), .B2(n_525), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_51), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_52), .B(n_989), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_53), .A2(n_336), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_54), .A2(n_204), .B1(n_632), .B2(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_55), .A2(n_213), .B1(n_519), .B2(n_550), .Y(n_1043) );
INVx1_ASAP7_75t_L g976 ( .A(n_56), .Y(n_976) );
INVx1_ASAP7_75t_L g803 ( .A(n_57), .Y(n_803) );
OA22x2_ASAP7_75t_L g427 ( .A1(n_58), .A2(n_162), .B1(n_421), .B2(n_425), .Y(n_427) );
INVx1_ASAP7_75t_L g455 ( .A(n_58), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_59), .A2(n_223), .B1(n_467), .B2(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_60), .A2(n_145), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_61), .A2(n_273), .B1(n_448), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_62), .A2(n_389), .B1(n_415), .B2(n_545), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_63), .A2(n_206), .B1(n_1089), .B2(n_1091), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_64), .A2(n_75), .B1(n_480), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_65), .A2(n_105), .B1(n_415), .B2(n_440), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_66), .A2(n_247), .B1(n_545), .B2(n_737), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_67), .A2(n_184), .B1(n_1079), .B2(n_1086), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_68), .A2(n_133), .B1(n_445), .B2(n_448), .Y(n_1012) );
INVx1_ASAP7_75t_L g1059 ( .A(n_69), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_70), .A2(n_173), .B1(n_528), .B2(n_569), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_71), .A2(n_100), .B1(n_528), .B2(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_72), .A2(n_370), .B1(n_664), .B2(n_665), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_73), .A2(n_193), .B1(n_445), .B2(n_525), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_76), .A2(n_254), .B1(n_664), .B2(n_665), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_77), .A2(n_172), .B1(n_658), .B2(n_659), .Y(n_794) );
INVx1_ASAP7_75t_L g1306 ( .A(n_78), .Y(n_1306) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_79), .A2(n_387), .B1(n_661), .B2(n_662), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_80), .A2(n_310), .B1(n_415), .B2(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_81), .B(n_175), .Y(n_402) );
INVx1_ASAP7_75t_L g424 ( .A(n_81), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_81), .A2(n_162), .B(n_457), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g1038 ( .A(n_82), .Y(n_1038) );
AO221x2_ASAP7_75t_L g1108 ( .A1(n_83), .A2(n_350), .B1(n_1079), .B2(n_1097), .C(n_1109), .Y(n_1108) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_84), .A2(n_556), .B(n_558), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_85), .A2(n_248), .B1(n_445), .B2(n_448), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_86), .A2(n_373), .B1(n_491), .B2(n_494), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_87), .A2(n_378), .B1(n_856), .B2(n_894), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g1111 ( .A1(n_88), .A2(n_338), .B1(n_1086), .B2(n_1112), .Y(n_1111) );
XNOR2x1_ASAP7_75t_L g972 ( .A(n_90), .B(n_973), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_90), .A2(n_361), .B1(n_1091), .B2(n_1099), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_91), .B(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_92), .A2(n_178), .B1(n_445), .B2(n_828), .Y(n_874) );
INVx1_ASAP7_75t_L g1083 ( .A(n_93), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_93), .B(n_285), .Y(n_1090) );
INVx1_ASAP7_75t_L g580 ( .A(n_94), .Y(n_580) );
AO22x1_ASAP7_75t_L g1109 ( .A1(n_95), .A2(n_183), .B1(n_1089), .B2(n_1105), .Y(n_1109) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_96), .A2(n_120), .B1(n_861), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_97), .A2(n_216), .B1(n_667), .B2(n_668), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_98), .A2(n_343), .B1(n_658), .B2(n_659), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_99), .B(n_537), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_101), .A2(n_276), .B1(n_673), .B2(n_674), .Y(n_688) );
INVx1_ASAP7_75t_L g926 ( .A(n_103), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_103), .A2(n_134), .B1(n_1100), .B2(n_1115), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_104), .A2(n_291), .B1(n_737), .B2(n_1000), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_106), .A2(n_217), .B1(n_634), .B2(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g728 ( .A(n_107), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_108), .A2(n_259), .B1(n_477), .B2(n_480), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_109), .A2(n_227), .B1(n_440), .B2(n_737), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_110), .Y(n_841) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_111), .A2(n_306), .B1(n_502), .B2(n_690), .C(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_112), .A2(n_243), .B1(n_598), .B2(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_113), .A2(n_265), .B1(n_561), .B2(n_681), .Y(n_680) );
XOR2x2_ASAP7_75t_L g897 ( .A(n_114), .B(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_115), .A2(n_221), .B1(n_744), .B2(n_745), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_116), .B(n_502), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_117), .A2(n_164), .B1(n_821), .B2(n_822), .Y(n_1061) );
INVx1_ASAP7_75t_L g1081 ( .A(n_118), .Y(n_1081) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_118), .B(n_398), .Y(n_1087) );
INVx1_ASAP7_75t_SL g1113 ( .A(n_118), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_119), .A2(n_151), .B1(n_521), .B2(n_600), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_121), .A2(n_333), .B1(n_545), .B2(n_600), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_122), .A2(n_257), .B1(n_681), .B2(n_932), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_123), .A2(n_322), .B1(n_445), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_124), .A2(n_356), .B1(n_561), .B2(n_681), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_126), .A2(n_159), .B1(n_1099), .B2(n_1105), .Y(n_1133) );
OAI22x1_ASAP7_75t_L g1296 ( .A1(n_126), .A2(n_1297), .B1(n_1310), .B2(n_1320), .Y(n_1296) );
NAND3xp33_ASAP7_75t_L g1297 ( .A(n_126), .B(n_1298), .C(n_1302), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_126), .A2(n_1322), .B1(n_1325), .B2(n_1327), .Y(n_1321) );
INVx1_ASAP7_75t_L g713 ( .A(n_127), .Y(n_713) );
INVx1_ASAP7_75t_L g981 ( .A(n_128), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_129), .A2(n_194), .B1(n_856), .B2(n_857), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_130), .A2(n_146), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_130), .A2(n_146), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_131), .A2(n_324), .B1(n_460), .B2(n_632), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_132), .B(n_906), .Y(n_905) );
XNOR2x1_ASAP7_75t_L g411 ( .A(n_135), .B(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_136), .A2(n_195), .B1(n_643), .B2(n_839), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_137), .A2(n_280), .B1(n_445), .B2(n_553), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_138), .A2(n_326), .B1(n_849), .B2(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g1020 ( .A(n_139), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_140), .A2(n_314), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_141), .A2(n_142), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_143), .A2(n_185), .B1(n_440), .B2(n_600), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_144), .A2(n_260), .B1(n_445), .B2(n_967), .Y(n_966) );
AO22x1_ASAP7_75t_L g696 ( .A1(n_147), .A2(n_296), .B1(n_667), .B2(n_668), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_148), .A2(n_179), .B1(n_614), .B2(n_616), .Y(n_859) );
INVx1_ASAP7_75t_L g540 ( .A(n_149), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_150), .A2(n_342), .B1(n_553), .B2(n_737), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g915 ( .A1(n_153), .A2(n_374), .B1(n_733), .B2(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_154), .A2(n_327), .B1(n_467), .B2(n_471), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_156), .A2(n_200), .B1(n_471), .B2(n_637), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_157), .A2(n_362), .B1(n_998), .B2(n_999), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_158), .A2(n_272), .B1(n_637), .B2(n_639), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_160), .B(n_671), .Y(n_950) );
INVx1_ASAP7_75t_L g439 ( .A(n_161), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_161), .B(n_212), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_161), .B(n_453), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_162), .B(n_293), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_163), .A2(n_225), .B1(n_1077), .B2(n_1084), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_165), .A2(n_348), .B1(n_497), .B2(n_500), .C(n_503), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_166), .A2(n_317), .B1(n_519), .B2(n_521), .Y(n_596) );
INVx1_ASAP7_75t_L g952 ( .A(n_167), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_168), .A2(n_332), .B1(n_445), .B2(n_553), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_169), .A2(n_351), .B1(n_537), .B2(n_856), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_171), .A2(n_353), .B1(n_667), .B2(n_668), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_174), .A2(n_390), .B1(n_553), .B2(n_839), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_175), .B(n_431), .Y(n_430) );
AO22x1_ASAP7_75t_L g697 ( .A1(n_176), .A2(n_329), .B1(n_661), .B2(n_662), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_180), .A2(n_266), .B1(n_460), .B2(n_632), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_181), .B(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_182), .A2(n_676), .B(n_677), .Y(n_675) );
XOR2x2_ASAP7_75t_SL g1006 ( .A(n_183), .B(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_186), .A2(n_220), .B1(n_991), .B2(n_992), .Y(n_990) );
AOI21xp33_ASAP7_75t_SL g586 ( .A1(n_187), .A2(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g1015 ( .A(n_188), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_189), .A2(n_325), .B1(n_497), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_190), .A2(n_349), .B1(n_661), .B2(n_662), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_192), .A2(n_379), .B1(n_467), .B2(n_640), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_196), .A2(n_690), .B(n_691), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_197), .A2(n_383), .B1(n_909), .B2(n_983), .Y(n_1315) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_198), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g903 ( .A(n_199), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_202), .A2(n_365), .B1(n_494), .B2(n_528), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g929 ( .A(n_203), .B(n_930), .Y(n_929) );
XNOR2x1_ASAP7_75t_L g1032 ( .A(n_206), .B(n_1033), .Y(n_1032) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_207), .A2(n_724), .B(n_727), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g1096 ( .A1(n_210), .A2(n_242), .B1(n_1079), .B2(n_1097), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_211), .A2(n_214), .B1(n_630), .B2(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g422 ( .A(n_212), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_218), .A2(n_321), .B1(n_1079), .B2(n_1086), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_219), .A2(n_360), .B1(n_467), .B2(n_523), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_222), .A2(n_252), .B1(n_661), .B2(n_662), .Y(n_796) );
INVx1_ASAP7_75t_L g589 ( .A(n_224), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_226), .A2(n_298), .B1(n_440), .B2(n_600), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_228), .A2(n_279), .B1(n_1079), .B2(n_1086), .Y(n_1106) );
INVx1_ASAP7_75t_L g884 ( .A(n_229), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_230), .A2(n_235), .B1(n_640), .B2(n_733), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_231), .A2(n_358), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_233), .A2(n_337), .B1(n_637), .B2(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_234), .A2(n_264), .B1(n_415), .B2(n_440), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_236), .A2(n_295), .B1(n_415), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_238), .A2(n_335), .B1(n_909), .B2(n_983), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_239), .A2(n_290), .B1(n_467), .B2(n_640), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_240), .A2(n_328), .B1(n_742), .B2(n_911), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g1312 ( .A1(n_241), .A2(n_261), .B1(n_1313), .B2(n_1314), .Y(n_1312) );
XNOR2x2_ASAP7_75t_L g683 ( .A(n_244), .B(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_245), .A2(n_318), .B1(n_1079), .B2(n_1084), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_246), .B(n_856), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_249), .A2(n_315), .B1(n_1089), .B2(n_1105), .Y(n_1125) );
INVx1_ASAP7_75t_L g1019 ( .A(n_250), .Y(n_1019) );
AOI21xp5_ASAP7_75t_SL g801 ( .A1(n_251), .A2(n_690), .B(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_253), .A2(n_308), .B1(n_673), .B2(n_674), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_255), .A2(n_385), .B1(n_467), .B2(n_523), .Y(n_551) );
XOR2xp5_ASAP7_75t_L g1322 ( .A(n_256), .B(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g881 ( .A(n_258), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_262), .A2(n_288), .B1(n_467), .B2(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g1053 ( .A(n_263), .Y(n_1053) );
AOI22xp5_ASAP7_75t_L g1098 ( .A1(n_263), .A2(n_344), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
INVx1_ASAP7_75t_L g984 ( .A(n_267), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_268), .A2(n_275), .B1(n_545), .B2(n_1319), .Y(n_1318) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_269), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_270), .A2(n_341), .B1(n_548), .B2(n_550), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_271), .A2(n_300), .B1(n_566), .B2(n_744), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_274), .A2(n_384), .B1(n_445), .B2(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_277), .Y(n_863) );
INVx1_ASAP7_75t_L g625 ( .A(n_278), .Y(n_625) );
AOI22xp5_ASAP7_75t_SL g672 ( .A1(n_281), .A2(n_382), .B1(n_673), .B2(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g1016 ( .A(n_282), .Y(n_1016) );
INVx1_ASAP7_75t_L g682 ( .A(n_283), .Y(n_682) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_285), .Y(n_403) );
AND2x4_ASAP7_75t_L g1082 ( .A(n_285), .B(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_SL g789 ( .A(n_286), .Y(n_789) );
INVx1_ASAP7_75t_L g805 ( .A(n_287), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_289), .A2(n_1036), .B(n_1037), .Y(n_1035) );
INVx1_ASAP7_75t_L g1022 ( .A(n_292), .Y(n_1022) );
INVx1_ASAP7_75t_L g437 ( .A(n_293), .Y(n_437) );
INVxp67_ASAP7_75t_L g489 ( .A(n_293), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_294), .A2(n_316), .B1(n_861), .B2(n_862), .Y(n_860) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_297), .A2(n_705), .B(n_720), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_297), .B(n_706), .C(n_710), .D(n_717), .Y(n_720) );
INVxp67_ASAP7_75t_R g750 ( .A(n_301), .Y(n_750) );
INVx1_ASAP7_75t_L g777 ( .A(n_301), .Y(n_777) );
INVx2_ASAP7_75t_L g398 ( .A(n_302), .Y(n_398) );
XNOR2x1_ASAP7_75t_L g541 ( .A(n_303), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g977 ( .A(n_304), .Y(n_977) );
INVx1_ASAP7_75t_L g810 ( .A(n_305), .Y(n_810) );
INVx1_ASAP7_75t_L g957 ( .A(n_309), .Y(n_957) );
INVx1_ASAP7_75t_L g1308 ( .A(n_311), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_312), .B(n_561), .Y(n_812) );
XNOR2x1_ASAP7_75t_L g943 ( .A(n_315), .B(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g692 ( .A(n_320), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_323), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_330), .A2(n_366), .B1(n_667), .B2(n_668), .Y(n_936) );
INVx1_ASAP7_75t_L g890 ( .A(n_331), .Y(n_890) );
INVx1_ASAP7_75t_L g678 ( .A(n_334), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_339), .A2(n_345), .B1(n_658), .B2(n_659), .Y(n_935) );
INVx1_ASAP7_75t_L g987 ( .A(n_340), .Y(n_987) );
AOI21xp33_ASAP7_75t_L g947 ( .A1(n_347), .A2(n_530), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g559 ( .A(n_352), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_355), .B(n_537), .Y(n_1039) );
INVx1_ASAP7_75t_L g954 ( .A(n_359), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_363), .A2(n_372), .B1(n_550), .B2(n_632), .Y(n_1068) );
AOI21xp5_ASAP7_75t_L g1302 ( .A1(n_364), .A2(n_1303), .B(n_1305), .Y(n_1302) );
INVx1_ASAP7_75t_L g800 ( .A(n_367), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_368), .Y(n_814) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_369), .Y(n_626) );
AOI21xp33_ASAP7_75t_SL g940 ( .A1(n_380), .A2(n_690), .B(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_381), .A2(n_388), .B1(n_587), .B2(n_745), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_386), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_404), .B(n_1072), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
BUFx10_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .C(n_403), .Y(n_395) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_396), .B(n_1293), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_396), .B(n_1294), .Y(n_1326) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OA21x2_ASAP7_75t_L g1327 ( .A1(n_397), .A2(n_1113), .B(n_1328), .Y(n_1327) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_398), .B(n_1081), .Y(n_1080) );
AND3x4_ASAP7_75t_L g1112 ( .A(n_398), .B(n_1082), .C(n_1113), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_399), .B(n_1294), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_400), .A2(n_509), .B(n_510), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g1294 ( .A(n_403), .Y(n_1294) );
XNOR2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_782), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_649), .B1(n_650), .B2(n_781), .Y(n_405) );
INVx2_ASAP7_75t_L g781 ( .A(n_406), .Y(n_781) );
AOI22x1_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_573), .B2(n_574), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OA22x2_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_512), .B1(n_513), .B2(n_572), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g572 ( .A(n_410), .Y(n_572) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND4xp75_ASAP7_75t_L g412 ( .A(n_413), .B(n_458), .C(n_475), .D(n_496), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_444), .Y(n_413) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx12f_ASAP7_75t_L g600 ( .A(n_416), .Y(n_600) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_416), .Y(n_737) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_428), .Y(n_416) );
AND2x4_ASAP7_75t_L g441 ( .A(n_417), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g468 ( .A(n_417), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g472 ( .A(n_417), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g661 ( .A(n_417), .B(n_428), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_417), .B(n_462), .Y(n_662) );
AND2x4_ASAP7_75t_L g664 ( .A(n_417), .B(n_469), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_417), .B(n_473), .Y(n_665) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_426), .Y(n_417) );
AND2x2_ASAP7_75t_L g479 ( .A(n_418), .B(n_427), .Y(n_479) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_427), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
NAND2xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_L g425 ( .A(n_421), .Y(n_425) );
INVx3_ASAP7_75t_L g431 ( .A(n_421), .Y(n_431) );
NAND2xp33_ASAP7_75t_L g438 ( .A(n_421), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_421), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_422), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_424), .A2(n_457), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g487 ( .A(n_427), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g446 ( .A(n_428), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g450 ( .A(n_428), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g549 ( .A(n_428), .B(n_447), .Y(n_549) );
AND2x4_ASAP7_75t_L g667 ( .A(n_428), .B(n_447), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_428), .B(n_451), .Y(n_668) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
OR2x2_ASAP7_75t_L g443 ( .A(n_429), .B(n_434), .Y(n_443) );
AND2x4_ASAP7_75t_L g469 ( .A(n_429), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g474 ( .A(n_429), .Y(n_474) );
AND2x2_ASAP7_75t_L g483 ( .A(n_429), .B(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_431), .B(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g453 ( .A(n_431), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_432), .B(n_452), .C(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g470 ( .A(n_435), .Y(n_470) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
BUFx3_ASAP7_75t_L g630 ( .A(n_440), .Y(n_630) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_441), .Y(n_521) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_441), .Y(n_545) );
BUFx6f_ASAP7_75t_L g1000 ( .A(n_441), .Y(n_1000) );
AND2x4_ASAP7_75t_L g465 ( .A(n_442), .B(n_451), .Y(n_465) );
AND2x4_ASAP7_75t_L g658 ( .A(n_442), .B(n_447), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_442), .B(n_451), .Y(n_659) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g462 ( .A(n_443), .Y(n_462) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx8_ASAP7_75t_L g839 ( .A(n_446), .Y(n_839) );
AND2x4_ASAP7_75t_L g461 ( .A(n_447), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g493 ( .A(n_447), .B(n_469), .Y(n_493) );
AND2x2_ASAP7_75t_L g502 ( .A(n_447), .B(n_473), .Y(n_502) );
AND2x2_ASAP7_75t_L g536 ( .A(n_447), .B(n_473), .Y(n_536) );
AND2x4_ASAP7_75t_L g681 ( .A(n_447), .B(n_469), .Y(n_681) );
INVx4_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx4_ASAP7_75t_L g525 ( .A(n_449), .Y(n_525) );
INVx4_ASAP7_75t_L g553 ( .A(n_449), .Y(n_553) );
INVx1_ASAP7_75t_L g601 ( .A(n_449), .Y(n_601) );
INVx2_ASAP7_75t_L g769 ( .A(n_449), .Y(n_769) );
INVx2_ASAP7_75t_SL g967 ( .A(n_449), .Y(n_967) );
INVx8_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g495 ( .A(n_451), .B(n_473), .Y(n_495) );
AND2x4_ASAP7_75t_L g674 ( .A(n_451), .B(n_473), .Y(n_674) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_456), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
BUFx3_ASAP7_75t_L g849 ( .A(n_460), .Y(n_849) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx12f_ASAP7_75t_L g518 ( .A(n_461), .Y(n_518) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_461), .Y(n_550) );
BUFx3_ASAP7_75t_L g739 ( .A(n_461), .Y(n_739) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_461), .Y(n_828) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_463), .Y(n_850) );
INVx1_ASAP7_75t_L g996 ( .A(n_463), .Y(n_996) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx5_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
INVx2_ASAP7_75t_L g546 ( .A(n_464), .Y(n_546) );
INVx3_ASAP7_75t_L g709 ( .A(n_464), .Y(n_709) );
INVx1_ASAP7_75t_L g1319 ( .A(n_464), .Y(n_1319) );
INVx6_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx12f_ASAP7_75t_L g632 ( .A(n_465), .Y(n_632) );
BUFx12f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g638 ( .A(n_468), .Y(n_638) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_468), .Y(n_733) );
AND2x4_ASAP7_75t_L g478 ( .A(n_469), .B(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g673 ( .A(n_469), .B(n_479), .Y(n_673) );
AND2x4_ASAP7_75t_L g473 ( .A(n_470), .B(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g837 ( .A(n_471), .Y(n_837) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
BUFx5_ASAP7_75t_L g640 ( .A(n_472), .Y(n_640) );
INVx1_ASAP7_75t_L g918 ( .A(n_472), .Y(n_918) );
AND2x4_ASAP7_75t_L g499 ( .A(n_473), .B(n_479), .Y(n_499) );
AND2x2_ASAP7_75t_L g690 ( .A(n_473), .B(n_479), .Y(n_690) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
INVx2_ASAP7_75t_L g615 ( .A(n_477), .Y(n_615) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g530 ( .A(n_478), .Y(n_530) );
INVx1_ASAP7_75t_L g570 ( .A(n_478), .Y(n_570) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_478), .Y(n_742) );
INVx2_ASAP7_75t_L g729 ( .A(n_480), .Y(n_729) );
INVx4_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g622 ( .A(n_481), .Y(n_622) );
INVx2_ASAP7_75t_L g774 ( .A(n_481), .Y(n_774) );
INVx2_ASAP7_75t_L g822 ( .A(n_481), .Y(n_822) );
INVx3_ASAP7_75t_L g991 ( .A(n_481), .Y(n_991) );
INVx5_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g585 ( .A(n_482), .Y(n_585) );
BUFx4f_ASAP7_75t_L g856 ( .A(n_482), .Y(n_856) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
AND2x4_ASAP7_75t_L g561 ( .A(n_483), .B(n_487), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g509 ( .A(n_485), .Y(n_509) );
INVx1_ASAP7_75t_L g958 ( .A(n_491), .Y(n_958) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g571 ( .A(n_492), .Y(n_571) );
BUFx6f_ASAP7_75t_L g912 ( .A(n_492), .Y(n_912) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_493), .Y(n_528) );
BUFx3_ASAP7_75t_L g821 ( .A(n_493), .Y(n_821) );
BUFx3_ASAP7_75t_L g619 ( .A(n_494), .Y(n_619) );
INVx3_ASAP7_75t_L g955 ( .A(n_494), .Y(n_955) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g567 ( .A(n_495), .Y(n_567) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_495), .Y(n_909) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_SL g983 ( .A(n_498), .Y(n_983) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g533 ( .A(n_499), .Y(n_533) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_499), .Y(n_587) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_499), .Y(n_676) );
BUFx3_ASAP7_75t_L g744 ( .A(n_499), .Y(n_744) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g799 ( .A1(n_501), .A2(n_800), .B(n_801), .Y(n_799) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_502), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
NOR2xp33_ASAP7_75t_R g624 ( .A(n_505), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_507), .Y(n_564) );
INVx2_ASAP7_75t_L g760 ( .A(n_507), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_507), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g906 ( .A(n_507), .Y(n_906) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g539 ( .A(n_508), .Y(n_539) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
XNOR2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_541), .Y(n_513) );
XOR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_540), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .C(n_522), .D(n_524), .Y(n_516) );
BUFx3_ASAP7_75t_L g634 ( .A(n_518), .Y(n_634) );
BUFx2_ASAP7_75t_L g643 ( .A(n_525), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .C(n_531), .D(n_534), .Y(n_526) );
BUFx3_ASAP7_75t_L g616 ( .A(n_528), .Y(n_616) );
INVx3_ASAP7_75t_L g888 ( .A(n_528), .Y(n_888) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g861 ( .A(n_533), .Y(n_861) );
BUFx3_ASAP7_75t_L g854 ( .A(n_535), .Y(n_854) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g557 ( .A(n_536), .Y(n_557) );
INVx2_ASAP7_75t_L g593 ( .A(n_536), .Y(n_593) );
INVx2_ASAP7_75t_L g1309 ( .A(n_537), .Y(n_1309) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_538), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g857 ( .A(n_538), .Y(n_857) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g679 ( .A(n_539), .Y(n_679) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_554), .Y(n_542) );
NAND4xp25_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .C(n_551), .D(n_552), .Y(n_543) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_545), .Y(n_843) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_549), .Y(n_598) );
NAND3xp33_ASAP7_75t_SL g554 ( .A(n_555), .B(n_565), .C(n_568), .Y(n_554) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_556), .Y(n_623) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g671 ( .A(n_557), .Y(n_671) );
INVx2_ASAP7_75t_L g726 ( .A(n_557), .Y(n_726) );
INVx2_ASAP7_75t_L g1024 ( .A(n_557), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_562), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g1037 ( .A1(n_560), .A2(n_1038), .B(n_1039), .Y(n_1037) );
INVx4_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_564), .B(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_564), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g894 ( .A(n_564), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_564), .B(n_942), .Y(n_941) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g745 ( .A(n_567), .Y(n_745) );
INVx2_ASAP7_75t_L g862 ( .A(n_567), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_567), .A2(n_880), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g886 ( .A(n_570), .Y(n_886) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_609), .B1(n_646), .B2(n_647), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g646 ( .A(n_577), .Y(n_646) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B(n_603), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_579), .B(n_594), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
NOR2xp67_ASAP7_75t_L g581 ( .A(n_582), .B(n_595), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .C(n_594), .Y(n_582) );
INVx1_ASAP7_75t_L g607 ( .A(n_583), .Y(n_607) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVxp67_ASAP7_75t_L g904 ( .A(n_585), .Y(n_904) );
BUFx3_ASAP7_75t_L g618 ( .A(n_587), .Y(n_618) );
INVxp67_ASAP7_75t_L g605 ( .A(n_590), .Y(n_605) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g755 ( .A(n_592), .Y(n_755) );
INVx2_ASAP7_75t_L g989 ( .A(n_592), .Y(n_989) );
INVx2_ASAP7_75t_L g1036 ( .A(n_592), .Y(n_1036) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g892 ( .A(n_593), .Y(n_892) );
INVx1_ASAP7_75t_L g608 ( .A(n_595), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .C(n_599), .D(n_602), .Y(n_595) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_600), .Y(n_642) );
BUFx12f_ASAP7_75t_L g998 ( .A(n_600), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_608), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .C(n_607), .Y(n_604) );
AO22x2_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_626), .B1(n_627), .B2(n_644), .Y(n_609) );
AO22x2_ASAP7_75t_L g648 ( .A1(n_610), .A2(n_626), .B1(n_627), .B2(n_644), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_620), .C(n_626), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND4xp75_ASAP7_75t_SL g644 ( .A(n_612), .B(n_628), .C(n_635), .D(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_617), .Y(n_612) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_615), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_975) );
INVx2_ASAP7_75t_L g1313 ( .A(n_615), .Y(n_1313) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_635), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_633), .Y(n_628) );
BUFx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g1002 ( .A(n_638), .Y(n_1002) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g845 ( .A(n_642), .Y(n_845) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_699), .B2(n_780), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_683), .Y(n_653) );
XOR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_682), .Y(n_654) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_669), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .C(n_663), .D(n_666), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .C(n_675), .D(n_680), .Y(n_669) );
INVx2_ASAP7_75t_L g806 ( .A(n_673), .Y(n_806) );
INVx2_ASAP7_75t_L g808 ( .A(n_674), .Y(n_808) );
INVx2_ASAP7_75t_L g953 ( .A(n_676), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_679), .B(n_713), .Y(n_712) );
INVx4_ASAP7_75t_L g992 ( .A(n_679), .Y(n_992) );
INVx1_ASAP7_75t_L g811 ( .A(n_681), .Y(n_811) );
OA22x2_ASAP7_75t_L g747 ( .A1(n_683), .A2(n_748), .B1(n_749), .B2(n_778), .Y(n_747) );
INVx1_ASAP7_75t_L g778 ( .A(n_683), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_693), .Y(n_684) );
AND4x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .C(n_688), .D(n_689), .Y(n_685) );
NOR4xp25_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .C(n_697), .D(n_698), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g780 ( .A(n_699), .Y(n_780) );
AO22x1_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_747), .B2(n_779), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
XNOR2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_721), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND3x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .C(n_717), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
XNOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_746), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g722 ( .A(n_723), .B(n_731), .C(n_735), .D(n_740), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B(n_730), .Y(n_727) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx2_ASAP7_75t_L g880 ( .A(n_744), .Y(n_880) );
INVx1_ASAP7_75t_L g779 ( .A(n_747), .Y(n_779) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B(n_775), .Y(n_749) );
NOR4xp75_ASAP7_75t_L g751 ( .A(n_752), .B(n_761), .C(n_765), .D(n_770), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND4xp75_ASAP7_75t_L g775 ( .A(n_753), .B(n_762), .C(n_766), .D(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_759), .B(n_949), .Y(n_948) );
NOR2xp33_ASAP7_75t_L g1058 ( .A(n_759), .B(n_1059), .Y(n_1058) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx2_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g776 ( .A(n_771), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B1(n_969), .B2(n_1071), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
XNOR2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_867), .Y(n_784) );
AO22x2_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_832), .B1(n_833), .B2(n_866), .Y(n_785) );
INVx1_ASAP7_75t_L g866 ( .A(n_786), .Y(n_866) );
OA22x2_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_813), .B1(n_830), .B2(n_831), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
XNOR2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
XNOR2xp5_ASAP7_75t_L g831 ( .A(n_789), .B(n_790), .Y(n_831) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_798), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_795), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_804), .C(n_809), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_804) );
INVxp67_ASAP7_75t_L g932 ( .A(n_808), .Y(n_932) );
OAI21xp5_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_811), .B(n_812), .Y(n_809) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_813), .Y(n_830) );
XNOR2x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
OR2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_824), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_820), .C(n_823), .Y(n_816) );
INVx2_ASAP7_75t_L g1017 ( .A(n_821), .Y(n_1017) );
NAND4xp25_ASAP7_75t_SL g824 ( .A(n_825), .B(n_826), .C(n_827), .D(n_829), .Y(n_824) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AO211x2_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_846), .B(n_864), .C(n_865), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_840), .Y(n_834) );
AO22x2_ASAP7_75t_L g865 ( .A1(n_835), .A2(n_847), .B1(n_863), .B2(n_1331), .Y(n_865) );
NAND2xp5_ASAP7_75t_SL g835 ( .A(n_836), .B(n_838), .Y(n_835) );
AO22x1_ASAP7_75t_L g864 ( .A1(n_840), .A2(n_858), .B1(n_863), .B2(n_1330), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_844), .B2(n_845), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NOR3xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_858), .C(n_863), .Y(n_846) );
NAND2x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_851), .Y(n_847) );
OA21x2_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B(n_855), .Y(n_851) );
INVx1_ASAP7_75t_SL g853 ( .A(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g882 ( .A(n_862), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_923), .B2(n_968), .Y(n_867) );
INVxp67_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_897), .B1(n_921), .B2(n_922), .Y(n_869) );
INVx2_ASAP7_75t_L g921 ( .A(n_870), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_871), .B(n_877), .Y(n_896) );
AND4x1_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .C(n_874), .D(n_875), .Y(n_871) );
AND2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_895), .Y(n_876) );
NOR3xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_883), .C(n_889), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_880), .B1(n_881), .B2(n_882), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_887), .B2(n_888), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_885), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OAI21xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_891), .B(n_893), .Y(n_889) );
INVxp67_ASAP7_75t_L g901 ( .A(n_891), .Y(n_901) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g922 ( .A(n_897), .Y(n_922) );
NOR2x1_ASAP7_75t_L g898 ( .A(n_899), .B(n_913), .Y(n_898) );
NAND3xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_907), .C(n_910), .Y(n_899) );
OAI21xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B(n_905), .Y(n_902) );
BUFx3_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx4_ASAP7_75t_L g985 ( .A(n_909), .Y(n_985) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx2_ASAP7_75t_L g979 ( .A(n_912), .Y(n_979) );
INVx2_ASAP7_75t_L g1314 ( .A(n_912), .Y(n_1314) );
NAND4xp25_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .C(n_919), .D(n_920), .Y(n_913) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g1004 ( .A(n_917), .Y(n_1004) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g968 ( .A(n_923), .Y(n_968) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
XNOR2xp5_ASAP7_75t_L g924 ( .A(n_925), .B(n_943), .Y(n_924) );
INVx3_ASAP7_75t_SL g1047 ( .A(n_925), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_925), .Y(n_1048) );
XNOR2x1_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
NOR2x1_ASAP7_75t_L g927 ( .A(n_928), .B(n_934), .Y(n_927) );
NAND3xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_931), .C(n_933), .Y(n_928) );
NAND4xp25_ASAP7_75t_SL g934 ( .A(n_935), .B(n_936), .C(n_937), .D(n_940), .Y(n_934) );
AND2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_960), .Y(n_944) );
NOR3xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_951), .C(n_956), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_950), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B1(n_954), .B2(n_955), .Y(n_951) );
OAI21xp33_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_958), .B(n_959), .Y(n_956) );
NOR2xp33_ASAP7_75t_SL g960 ( .A(n_961), .B(n_964), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
INVx1_ASAP7_75t_L g1071 ( .A(n_969), .Y(n_1071) );
AO22x1_ASAP7_75t_L g969 ( .A1(n_970), .A2(n_971), .B1(n_1028), .B2(n_1029), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_1006), .B1(n_1026), .B2(n_1027), .Y(n_971) );
INVx1_ASAP7_75t_SL g1027 ( .A(n_972), .Y(n_1027) );
AND2x4_ASAP7_75t_L g973 ( .A(n_974), .B(n_993), .Y(n_973) );
NOR3xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_980), .C(n_986), .Y(n_974) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B1(n_984), .B2(n_985), .Y(n_980) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
OAI21xp33_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_988), .B(n_990), .Y(n_986) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1307 ( .A(n_991), .Y(n_1307) );
AND4x1_ASAP7_75t_L g993 ( .A(n_994), .B(n_997), .C(n_1001), .D(n_1005), .Y(n_993) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
BUFx3_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
BUFx4f_ASAP7_75t_L g1300 ( .A(n_1002), .Y(n_1300) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1006), .Y(n_1026) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1013), .Y(n_1007) );
AND4x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .C(n_1011), .D(n_1012), .Y(n_1008) );
NOR3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1018), .C(n_1021), .Y(n_1013) );
OAI21xp33_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1023), .B(n_1025), .Y(n_1021) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1024), .Y(n_1304) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
OAI22x1_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1031), .B1(n_1050), .B2(n_1069), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
OA22x2_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1047), .B1(n_1048), .B2(n_1049), .Y(n_1031) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1032), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1042), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1040), .C(n_1041), .Y(n_1034) );
NAND4xp25_ASAP7_75t_SL g1042 ( .A(n_1043), .B(n_1044), .C(n_1045), .D(n_1046), .Y(n_1042) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1052), .Y(n_1070) );
XNOR2x1_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
NOR4xp75_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1060), .C(n_1063), .D(n_1066), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1062), .Y(n_1060) );
NAND2xp5_ASAP7_75t_SL g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
NAND2xp5_ASAP7_75t_SL g1066 ( .A(n_1067), .B(n_1068), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
OAI221xp5_ASAP7_75t_SL g1072 ( .A1(n_1073), .A2(n_1288), .B1(n_1290), .B2(n_1295), .C(n_1321), .Y(n_1072) );
AND5x1_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1224), .C(n_1253), .D(n_1268), .E(n_1275), .Y(n_1073) );
AOI211xp5_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1092), .B(n_1183), .C(n_1200), .Y(n_1074) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1075), .B(n_1119), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_1075), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1088), .Y(n_1075) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx3_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
AND2x4_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1082), .Y(n_1079) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_1080), .B(n_1090), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1080), .B(n_1090), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1080), .B(n_1090), .Y(n_1115) );
AND2x4_ASAP7_75t_L g1086 ( .A(n_1082), .B(n_1087), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1097 ( .A(n_1082), .B(n_1087), .Y(n_1097) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_1086), .Y(n_1085) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_1087), .B(n_1090), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1087), .B(n_1090), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1087), .B(n_1090), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g1328 ( .A(n_1090), .Y(n_1328) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_1091), .Y(n_1289) );
NAND5xp2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1150), .C(n_1161), .D(n_1165), .E(n_1178), .Y(n_1092) );
AOI21xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1116), .B(n_1127), .Y(n_1093) );
OAI21xp5_ASAP7_75t_L g1198 ( .A1(n_1094), .A2(n_1164), .B(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1101), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1095), .B(n_1137), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1095), .B(n_1144), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1095), .B(n_1110), .Y(n_1149) );
CKINVDCx6p67_ASAP7_75t_R g1153 ( .A(n_1095), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1095), .B(n_1142), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1095), .B(n_1170), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1095), .B(n_1169), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1095), .B(n_1107), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1095), .B(n_1179), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1098), .Y(n_1095) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1101), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1107), .Y(n_1101) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1102), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1102), .B(n_1181), .Y(n_1180) );
INVx3_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1103), .B(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1103), .Y(n_1148) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1103), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1103), .B(n_1153), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1103), .B(n_1182), .Y(n_1205) );
NOR2xp33_ASAP7_75t_L g1240 ( .A(n_1103), .B(n_1132), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1103), .B(n_1139), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1106), .Y(n_1103) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1107), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1107), .B(n_1153), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1107), .B(n_1193), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1110), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1108), .B(n_1137), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1108), .B(n_1110), .Y(n_1155) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1108), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1108), .B(n_1153), .Y(n_1209) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1110), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1110), .B(n_1170), .Y(n_1169) );
AOI31xp33_ASAP7_75t_L g1260 ( .A1(n_1110), .A2(n_1210), .A3(n_1261), .B(n_1263), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1114), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1116), .B(n_1247), .Y(n_1266) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
NOR3xp33_ASAP7_75t_L g1283 ( .A(n_1117), .B(n_1141), .C(n_1190), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1122), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1118), .B(n_1157), .Y(n_1166) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1118), .Y(n_1210) );
NOR2xp33_ASAP7_75t_L g1218 ( .A(n_1118), .B(n_1219), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1118), .B(n_1123), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1118), .B(n_1196), .Y(n_1280) );
INVx4_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1119), .B(n_1130), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1119), .B(n_1163), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1119), .B(n_1124), .Y(n_1177) );
NAND3xp33_ASAP7_75t_L g1267 ( .A(n_1119), .B(n_1169), .C(n_1240), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
INVxp67_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1123), .B(n_1132), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1123), .B(n_1131), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1123), .B(n_1132), .Y(n_1182) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1123), .Y(n_1196) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1124), .B(n_1132), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1126), .Y(n_1124) );
OAI211xp5_ASAP7_75t_SL g1127 ( .A1(n_1128), .A2(n_1135), .B(n_1138), .C(n_1145), .Y(n_1127) );
A2O1A1O1Ixp25_ASAP7_75t_L g1255 ( .A1(n_1128), .A2(n_1235), .B(n_1256), .C(n_1257), .D(n_1260), .Y(n_1255) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
AOI211xp5_ASAP7_75t_L g1246 ( .A1(n_1130), .A2(n_1194), .B(n_1235), .C(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1131), .Y(n_1176) );
INVx4_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1132), .B(n_1148), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1132), .B(n_1148), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1134), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1137), .B(n_1153), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
AOI22xp5_ASAP7_75t_L g1150 ( .A1(n_1139), .A2(n_1151), .B1(n_1156), .B2(n_1158), .Y(n_1150) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1139), .Y(n_1199) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1142), .B(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1142), .B(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1142), .Y(n_1204) );
AOI322xp5_ASAP7_75t_L g1201 ( .A1(n_1143), .A2(n_1156), .A3(n_1160), .B1(n_1180), .B2(n_1202), .C1(n_1205), .C2(n_1206), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1143), .B(n_1179), .Y(n_1278) );
NOR2x1_ASAP7_75t_L g1154 ( .A(n_1144), .B(n_1155), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1144), .B(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1144), .B(n_1250), .Y(n_1249) );
NOR2x1_ASAP7_75t_L g1271 ( .A(n_1144), .B(n_1251), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1149), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1148), .B(n_1209), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1148), .B(n_1259), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1149), .B(n_1159), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1151), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
NOR2xp33_ASAP7_75t_L g1225 ( .A(n_1152), .B(n_1226), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1154), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1153), .B(n_1179), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1153), .B(n_1169), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1153), .B(n_1170), .Y(n_1286) );
OAI21xp5_ASAP7_75t_L g1252 ( .A1(n_1154), .A2(n_1156), .B(n_1250), .Y(n_1252) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1155), .Y(n_1179) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1171 ( .A(n_1159), .B(n_1172), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g1222 ( .A(n_1159), .B(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1160), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g1220 ( .A1(n_1162), .A2(n_1221), .B(n_1222), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1163), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1167), .B1(n_1171), .B2(n_1173), .Y(n_1165) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
OAI21xp33_ASAP7_75t_L g1276 ( .A1(n_1168), .A2(n_1235), .B(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1169), .Y(n_1203) );
OAI211xp5_ASAP7_75t_L g1284 ( .A1(n_1169), .A2(n_1186), .B(n_1285), .C(n_1287), .Y(n_1284) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1171), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1177), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1175), .Y(n_1191) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1176), .Y(n_1214) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1177), .Y(n_1264) );
AOI221xp5_ASAP7_75t_L g1275 ( .A1(n_1177), .A2(n_1271), .B1(n_1276), .B2(n_1279), .C(n_1281), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1179), .B(n_1193), .Y(n_1197) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1182), .A2(n_1188), .B1(n_1194), .B2(n_1197), .Y(n_1187) );
O2A1O1Ixp33_ASAP7_75t_SL g1183 ( .A1(n_1184), .A2(n_1185), .B(n_1187), .C(n_1198), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_1184), .B(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
OAI211xp5_ASAP7_75t_L g1233 ( .A1(n_1189), .A2(n_1195), .B(n_1234), .C(n_1235), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1192), .Y(n_1189) );
HB1xp67_ASAP7_75t_L g1226 ( .A(n_1190), .Y(n_1226) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1191), .Y(n_1243) );
O2A1O1Ixp33_ASAP7_75t_L g1253 ( .A1(n_1192), .A2(n_1225), .B(n_1254), .C(n_1255), .Y(n_1253) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx3_ASAP7_75t_SL g1195 ( .A(n_1196), .Y(n_1195) );
OAI221xp5_ASAP7_75t_L g1227 ( .A1(n_1196), .A2(n_1199), .B1(n_1228), .B2(n_1230), .C(n_1231), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1196), .B(n_1219), .Y(n_1245) );
NOR4xp25_ASAP7_75t_L g1237 ( .A(n_1197), .B(n_1238), .C(n_1241), .D(n_1245), .Y(n_1237) );
OAI221xp5_ASAP7_75t_L g1200 ( .A1(n_1201), .A2(n_1210), .B1(n_1211), .B2(n_1217), .C(n_1220), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1208), .Y(n_1206) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
A2O1A1Ixp33_ASAP7_75t_SL g1268 ( .A1(n_1210), .A2(n_1269), .B(n_1271), .C(n_1272), .Y(n_1268) );
INVxp67_ASAP7_75t_SL g1211 ( .A(n_1212), .Y(n_1211) );
NOR2xp33_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1215), .Y(n_1212) );
OAI221xp5_ASAP7_75t_L g1236 ( .A1(n_1213), .A2(n_1237), .B1(n_1246), .B2(n_1248), .C(n_1252), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1213), .B(n_1278), .Y(n_1277) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1270 ( .A(n_1214), .Y(n_1270) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1216), .B(n_1229), .Y(n_1228) );
OAI311xp33_ASAP7_75t_L g1224 ( .A1(n_1217), .A2(n_1225), .A3(n_1227), .B1(n_1233), .C1(n_1236), .Y(n_1224) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1219), .Y(n_1235) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1221), .Y(n_1230) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1244), .Y(n_1241) );
HB1xp67_ASAP7_75t_L g1274 ( .A(n_1242), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
OAI211xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B(n_1266), .C(n_1267), .Y(n_1263) );
CKINVDCx16_ASAP7_75t_R g1269 ( .A(n_1270), .Y(n_1269) );
INVxp67_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1284), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
HB1xp67_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
AND4x1_ASAP7_75t_L g1320 ( .A(n_1298), .B(n_1302), .C(n_1311), .D(n_1316), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1301), .Y(n_1298) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B1(n_1308), .B2(n_1309), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1316), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1315), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1318), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g1324 ( .A(n_1320), .Y(n_1324) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
BUFx2_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
endmodule