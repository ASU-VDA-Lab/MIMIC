module fake_jpeg_31707_n_36 (n_3, n_2, n_1, n_0, n_4, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_SL g5 ( 
.A(n_1),
.Y(n_5)
);

BUFx3_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_3),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_9),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_8),
.B(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_0),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_20),
.B(n_5),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_17),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_17),
.B(n_13),
.C(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_28),
.C(n_22),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_29),
.B2(n_16),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_29),
.C(n_27),
.Y(n_32)
);

OAI33xp33_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_10),
.A3(n_20),
.B1(n_8),
.B2(n_21),
.B3(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_21),
.Y(n_36)
);


endmodule