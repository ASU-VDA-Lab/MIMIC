module fake_jpeg_28792_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_36),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_66),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_58),
.B1(n_57),
.B2(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_25),
.B1(n_45),
.B2(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_96),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_73),
.B1(n_62),
.B2(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_94),
.B1(n_83),
.B2(n_95),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_70),
.B(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_63),
.C(n_57),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.C(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_29),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_51),
.B1(n_67),
.B2(n_52),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_64),
.B(n_63),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_68),
.B1(n_64),
.B2(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_54),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_103),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_72),
.B(n_60),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_105),
.Y(n_134)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_10),
.C(n_12),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_113),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_70),
.B(n_8),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_13),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_28),
.C(n_41),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_27),
.B1(n_40),
.B2(n_39),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_115),
.B1(n_12),
.B2(n_13),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_20),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_7),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_14),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_34),
.C(n_35),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_38),
.B1(n_48),
.B2(n_122),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_33),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_114),
.B1(n_112),
.B2(n_100),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_15),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_15),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_19),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_30),
.C(n_32),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_138),
.A2(n_147),
.B1(n_134),
.B2(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_148),
.C(n_149),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_144),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_145),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_119),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_124),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_147),
.B1(n_140),
.B2(n_131),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_137),
.C(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_151),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_159),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_157),
.B1(n_139),
.B2(n_158),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_156),
.B(n_150),
.C(n_155),
.D(n_153),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_156),
.B(n_141),
.C(n_144),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_136),
.Y(n_164)
);


endmodule