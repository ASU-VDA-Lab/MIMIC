module real_jpeg_31156_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_679, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_678, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_679;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_678;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_666;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_586;
wire n_572;
wire n_120;
wire n_155;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_659;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_625;
wire n_85;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_0),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_2),
.A2(n_34),
.B1(n_242),
.B2(n_246),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_2),
.A2(n_34),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_2),
.A2(n_34),
.B1(n_625),
.B2(n_631),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_3),
.A2(n_140),
.B1(n_223),
.B2(n_227),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_3),
.A2(n_140),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_3),
.A2(n_140),
.B1(n_534),
.B2(n_538),
.Y(n_533)
);

AO22x1_ASAP7_75t_L g255 ( 
.A1(n_4),
.A2(n_256),
.B1(n_259),
.B2(n_262),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_4),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g316 ( 
.A1(n_4),
.A2(n_262),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_4),
.A2(n_262),
.B1(n_617),
.B2(n_618),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g651 ( 
.A1(n_4),
.A2(n_262),
.B1(n_652),
.B2(n_655),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_85),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_5),
.A2(n_337),
.B(n_339),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_5),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_5),
.A2(n_85),
.B1(n_382),
.B2(n_386),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_168),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_6),
.A2(n_173),
.B1(n_288),
.B2(n_291),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_6),
.A2(n_173),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_6),
.A2(n_173),
.B1(n_212),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_7),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_10),
.Y(n_452)
);

AOI22x1_ASAP7_75t_SL g125 ( 
.A1(n_11),
.A2(n_126),
.B1(n_129),
.B2(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_11),
.A2(n_134),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_11),
.A2(n_91),
.B1(n_134),
.B2(n_463),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_11),
.A2(n_134),
.B1(n_478),
.B2(n_480),
.Y(n_477)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_12),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_13),
.A2(n_187),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_13),
.A2(n_234),
.B1(n_369),
.B2(n_372),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_13),
.A2(n_234),
.B1(n_425),
.B2(n_428),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_13),
.A2(n_234),
.B1(n_472),
.B2(n_476),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_14),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_14),
.A2(n_94),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_14),
.A2(n_94),
.B1(n_296),
.B2(n_299),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_14),
.A2(n_587),
.B(n_592),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_14),
.B(n_593),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_15),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_15),
.A2(n_52),
.B1(n_91),
.B2(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_15),
.A2(n_52),
.B1(n_531),
.B2(n_598),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_15),
.A2(n_52),
.B1(n_235),
.B2(n_643),
.Y(n_642)
);

OAI321xp33_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_21),
.A3(n_666),
.B1(n_672),
.B2(n_674),
.C(n_678),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_16),
.B(n_673),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_17),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_17),
.A2(n_205),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_17),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_17),
.B(n_177),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_17),
.A2(n_39),
.B1(n_471),
.B2(n_489),
.Y(n_488)
);

OAI32xp33_ASAP7_75t_L g508 ( 
.A1(n_17),
.A2(n_147),
.A3(n_509),
.B1(n_513),
.B2(n_517),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_17),
.A2(n_390),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_18),
.Y(n_355)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_19),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_19),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_21),
.B(n_675),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_574),
.B(n_659),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_410),
.B(n_569),
.Y(n_23)
);

NAND4xp25_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_304),
.C(n_343),
.D(n_403),
.Y(n_24)
);

A2O1A1O1Ixp25_ASAP7_75t_L g569 ( 
.A1(n_25),
.A2(n_304),
.B(n_570),
.C(n_572),
.D(n_573),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_263),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_26),
.B(n_263),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_184),
.C(n_239),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_28),
.B(n_239),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_98),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_29),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_57),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_30),
.B(n_57),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_39),
.B1(n_45),
.B2(n_53),
.Y(n_30)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_31),
.Y(n_216)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_33),
.Y(n_212)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_33),
.Y(n_388)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_38),
.Y(n_475)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_39),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_39),
.A2(n_45),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_39),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_39),
.A2(n_471),
.B1(n_477),
.B2(n_484),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_42),
.Y(n_380)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_44),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_50),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_51),
.Y(n_258)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_51),
.Y(n_385)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_51),
.Y(n_483)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_54),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.Y(n_496)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_79),
.B1(n_89),
.B2(n_90),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_58),
.A2(n_89),
.B1(n_90),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_58),
.A2(n_89),
.B1(n_241),
.B2(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_58),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_58),
.A2(n_79),
.B1(n_89),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_58),
.A2(n_89),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_58),
.A2(n_555),
.B(n_556),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_58),
.B(n_89),
.Y(n_603)
);

AO21x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_66),
.B(n_73),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_65),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_65),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_65),
.Y(n_464)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_65),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_66),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_67),
.Y(n_245)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g537 ( 
.A(n_69),
.Y(n_537)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_74),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_74),
.Y(n_457)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_78),
.Y(n_214)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_84),
.Y(n_248)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_89),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_89),
.B(n_390),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_93),
.Y(n_319)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_93),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_97),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_144),
.B1(n_145),
.B2(n_183),
.Y(n_98)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_125),
.B1(n_135),
.B2(n_136),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_101),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_101),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_101),
.A2(n_238),
.B1(n_287),
.B2(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_101),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_101),
.A2(n_286),
.B1(n_336),
.B2(n_586),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_105),
.Y(n_630)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_106),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_106),
.Y(n_657)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_110),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_110),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_118),
.B1(n_121),
.B2(n_124),
.Y(n_114)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_116),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_117),
.Y(n_371)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_123),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_123),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_123),
.Y(n_376)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_132),
.Y(n_291)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_132),
.Y(n_644)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_133),
.Y(n_591)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_135),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_135),
.A2(n_233),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

NOR2x1_ASAP7_75t_R g389 ( 
.A(n_135),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_136),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_139),
.Y(n_338)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

BUFx4f_ASAP7_75t_SL g631 ( 
.A(n_143),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22x1_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_167),
.B1(n_176),
.B2(n_178),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_146),
.A2(n_167),
.B1(n_176),
.B2(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_146),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_146),
.A2(n_176),
.B1(n_222),
.B2(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_146),
.A2(n_176),
.B1(n_360),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_146),
.A2(n_176),
.B1(n_368),
.B2(n_529),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_146),
.A2(n_176),
.B1(n_597),
.B2(n_601),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_146),
.A2(n_176),
.B1(n_597),
.B2(n_616),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_154),
.B(n_159),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_149),
.Y(n_617)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_165),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_161),
.Y(n_428)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_172),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g619 ( 
.A(n_175),
.Y(n_619)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22x1_ASAP7_75t_L g292 ( 
.A1(n_177),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_177),
.A2(n_293),
.B1(n_295),
.B2(n_325),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g639 ( 
.A1(n_177),
.A2(n_293),
.B(n_640),
.Y(n_639)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_182),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_184),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_219),
.C(n_230),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_185),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_209),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_186),
.A2(n_209),
.B1(n_210),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_186),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_189),
.A3(n_190),
.B1(n_195),
.B2(n_204),
.Y(n_186)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_211),
.A2(n_215),
.B1(n_379),
.B2(n_381),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_214),
.Y(n_433)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_215),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_215),
.A2(n_381),
.B1(n_456),
.B2(n_522),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_221),
.B(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_226),
.Y(n_362)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_226),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_231),
.Y(n_396)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_249),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_248),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

INVx3_ASAP7_75t_SL g280 ( 
.A(n_251),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_254),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_254),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_254),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_260),
.Y(n_476)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_306),
.C(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_281),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

XNOR2x2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_277),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_278),
.Y(n_333)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_278),
.A2(n_579),
.B1(n_580),
.B2(n_679),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_282),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_286),
.Y(n_623)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_SL g594 ( 
.A(n_291),
.Y(n_594)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_296),
.Y(n_530)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_299),
.Y(n_531)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_305),
.B(n_308),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_309),
.B(n_332),
.C(n_341),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_332),
.B1(n_341),
.B2(n_342),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_324),
.B(n_331),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_324),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_315)
);

NAND2x1_ASAP7_75t_L g602 ( 
.A(n_316),
.B(n_603),
.Y(n_602)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_321),
.A2(n_323),
.B1(n_418),
.B2(n_424),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_321),
.A2(n_323),
.B1(n_533),
.B2(n_543),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_321),
.B(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_325),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_330),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_331),
.Y(n_582)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_333),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_335),
.Y(n_580)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_393),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_344),
.B(n_393),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_366),
.C(n_391),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_345),
.B(n_566),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_347),
.A2(n_622),
.B1(n_623),
.B2(n_624),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_347),
.A2(n_623),
.B1(n_624),
.B2(n_642),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_347),
.A2(n_623),
.B1(n_642),
.B2(n_651),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_347),
.A2(n_623),
.B(n_651),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_359),
.Y(n_350)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_352),
.Y(n_557)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_355),
.Y(n_520)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_355),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_366),
.B(n_391),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_377),
.C(n_389),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_367),
.B(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_377),
.A2(n_378),
.B1(n_389),
.B2(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_389),
.Y(n_551)
);

OAI21xp33_ASAP7_75t_SL g418 ( 
.A1(n_390),
.A2(n_419),
.B(n_421),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_390),
.B(n_484),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_390),
.B(n_518),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_397),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_405),
.C(n_406),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_399),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.C(n_402),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_404),
.B(n_407),
.C(n_571),
.Y(n_570)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

AOI21x1_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_564),
.B(n_568),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_547),
.B(n_563),
.Y(n_411)
);

AOI21x1_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_504),
.B(n_546),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_467),
.B(n_503),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_443),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_415),
.B(n_443),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_429),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_416),
.A2(n_417),
.B1(n_429),
.B2(n_430),
.Y(n_495)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_438),
.B1(n_439),
.B2(n_442),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_458),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_460),
.C(n_465),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_453),
.B2(n_455),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_445),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_446),
.Y(n_499)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_460),
.B1(n_465),
.B2(n_466),
.Y(n_458)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_459),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_460),
.Y(n_466)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

OAI31xp33_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_494),
.A3(n_500),
.B(n_502),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_487),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_486),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_470),
.B(n_486),
.Y(n_501)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_491),
.Y(n_487)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_496),
.Y(n_502)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_SL g546 ( 
.A(n_505),
.B(n_506),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_527),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_532),
.C(n_545),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_521),
.B1(n_525),
.B2(n_526),
.Y(n_507)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_508),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_508),
.B(n_526),
.Y(n_553)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_532),
.B1(n_544),
.B2(n_545),
.Y(n_527)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_528),
.Y(n_545)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_532),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_533),
.Y(n_555)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_562),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_562),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_549),
.A2(n_552),
.B1(n_560),
.B2(n_561),
.Y(n_548)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_549),
.Y(n_561)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_552),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_553),
.A2(n_554),
.B1(n_558),
.B2(n_559),
.Y(n_552)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_553),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_554),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_558),
.C(n_561),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_565),
.B(n_567),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_567),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_632),
.C(n_649),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_576),
.B(n_605),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_577),
.B(n_604),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_577),
.B(n_604),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_581),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_582),
.C(n_583),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_583),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_595),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_584),
.B(n_610),
.C(n_611),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_621),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_584),
.B(n_609),
.C(n_646),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_586),
.Y(n_622)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_590),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_602),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_596),
.Y(n_611)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_602),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_602),
.B(n_615),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_602),
.B(n_615),
.C(n_621),
.Y(n_636)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_606),
.A2(n_662),
.B(n_663),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_608),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_607),
.B(n_608),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_609),
.B(n_612),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_620),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_613),
.A2(n_614),
.B1(n_647),
.B2(n_648),
.Y(n_646)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_616),
.Y(n_640)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_621),
.Y(n_648)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_633),
.A2(n_661),
.B(n_664),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_634),
.B(n_645),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_634),
.B(n_645),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_635),
.A2(n_636),
.B1(n_637),
.B2(n_638),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_635),
.B(n_639),
.C(n_641),
.Y(n_658)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_639),
.B(n_641),
.Y(n_638)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_644),
.Y(n_654)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_SL g659 ( 
.A1(n_649),
.A2(n_660),
.B(n_665),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_658),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_650),
.B(n_658),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_650),
.B(n_668),
.Y(n_667)
);

CKINVDCx16_ASAP7_75t_R g671 ( 
.A(n_650),
.Y(n_671)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_654),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_656),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_666),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_667),
.B(n_670),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_669),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_669),
.B(n_671),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_672),
.B(n_676),
.Y(n_675)
);


endmodule