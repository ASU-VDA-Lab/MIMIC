module fake_jpeg_31929_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_1),
.Y(n_100)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_25),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_14),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_56),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_35),
.B1(n_36),
.B2(n_30),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_6),
.B(n_7),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_37),
.B1(n_33),
.B2(n_20),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_77),
.B1(n_78),
.B2(n_86),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_35),
.C(n_31),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_61),
.C(n_90),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_68),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_87),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_88),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_32),
.B1(n_36),
.B2(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_19),
.B(n_31),
.C(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_37),
.B1(n_33),
.B2(n_20),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_1),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_99),
.A2(n_60),
.B1(n_4),
.B2(n_6),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_102),
.B(n_120),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_114),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_3),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_127),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_90),
.B(n_75),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_8),
.C(n_9),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_66),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_73),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_80),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_82),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_72),
.B1(n_64),
.B2(n_96),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_145),
.B1(n_155),
.B2(n_125),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_159),
.B(n_11),
.Y(n_185)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_148),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_64),
.B1(n_96),
.B2(n_97),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_143),
.B1(n_153),
.B2(n_154),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_83),
.B1(n_72),
.B2(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_146),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_103),
.B1(n_117),
.B2(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_110),
.B(n_70),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_83),
.B1(n_92),
.B2(n_93),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_79),
.B1(n_71),
.B2(n_92),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_79),
.B1(n_71),
.B2(n_84),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_113),
.B1(n_112),
.B2(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_82),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_8),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_11),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_8),
.B1(n_11),
.B2(n_63),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_162),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_130),
.B(n_105),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_170),
.B(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_166),
.Y(n_204)
);

OR2x2_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_115),
.Y(n_167)
);

AO32x1_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_135),
.A3(n_145),
.B1(n_148),
.B2(n_142),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_174),
.B(n_175),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_142),
.B(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_181),
.B1(n_129),
.B2(n_107),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_179),
.B1(n_146),
.B2(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_182),
.B(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_105),
.B1(n_101),
.B2(n_121),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_155),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_190),
.B(n_192),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_176),
.B1(n_165),
.B2(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_149),
.B(n_140),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_194),
.C(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_138),
.C(n_144),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_140),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_184),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_160),
.C(n_151),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_147),
.A3(n_152),
.B1(n_115),
.B2(n_121),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_129),
.B(n_63),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_164),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_170),
.B(n_173),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_167),
.B1(n_165),
.B2(n_183),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_166),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_218),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_174),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_198),
.C(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_226),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_215),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_197),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_200),
.C(n_192),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_187),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_234),
.Y(n_239)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_236),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_209),
.B(n_206),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_228),
.B(n_210),
.C(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_218),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_213),
.B(n_209),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_206),
.B1(n_205),
.B2(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

NAND4xp25_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_179),
.C(n_202),
.D(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_204),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_228),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_246),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_247),
.B(n_240),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_213),
.A3(n_235),
.B1(n_207),
.B2(n_204),
.C1(n_214),
.C2(n_177),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_238),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_245),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_240),
.B(n_172),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_252),
.C(n_240),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_254),
.B(n_107),
.CI(n_248),
.CON(n_255),
.SN(n_255)
);


endmodule