module fake_netlist_1_3385_n_561 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_561);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_561;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_75), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_67), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_15), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_63), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_8), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_58), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_24), .Y(n_83) );
INVx1_ASAP7_75t_SL g84 ( .A(n_73), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_22), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_46), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_52), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_36), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_72), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_53), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_60), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_61), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_43), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_31), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_64), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_3), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_74), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_28), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_40), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_70), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_21), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_42), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_23), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_44), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_11), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_54), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_25), .B(n_29), .Y(n_107) );
NOR2xp67_ASAP7_75t_L g108 ( .A(n_17), .B(n_9), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_1), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_47), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_41), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_38), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_39), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_49), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
CKINVDCx8_ASAP7_75t_R g118 ( .A(n_78), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_79), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_82), .Y(n_121) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_100), .A2(n_27), .B(n_71), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_109), .Y(n_123) );
INVx6_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_79), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_126) );
NOR2x1_ASAP7_75t_L g127 ( .A(n_108), .B(n_4), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_106), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_105), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_106), .B(n_4), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_105), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_100), .Y(n_135) );
BUFx8_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_97), .B(n_5), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_132), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_132), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_117), .B(n_99), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g144 ( .A1(n_118), .A2(n_116), .B1(n_113), .B2(n_91), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_134), .B(n_110), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_135), .Y(n_147) );
INVx2_ASAP7_75t_SL g148 ( .A(n_132), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
AO22x2_ASAP7_75t_L g150 ( .A1(n_117), .A2(n_92), .B1(n_90), .B2(n_112), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_134), .B(n_80), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_119), .A2(n_116), .B1(n_113), .B2(n_111), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_130), .B(n_101), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_128), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_135), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_130), .B(n_80), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
NAND3xp33_ASAP7_75t_L g162 ( .A(n_131), .B(n_104), .C(n_115), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_131), .B(n_114), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_137), .B(n_114), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_120), .Y(n_165) );
INVx8_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
AND2x6_ASAP7_75t_SL g167 ( .A(n_151), .B(n_138), .Y(n_167) );
INVx8_ASAP7_75t_L g168 ( .A(n_166), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_153), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_158), .B(n_129), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_153), .A2(n_91), .B1(n_111), .B2(n_137), .Y(n_174) );
INVx8_ASAP7_75t_L g175 ( .A(n_166), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_166), .B(n_121), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_149), .B(n_121), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
AND2x6_ASAP7_75t_SL g179 ( .A(n_151), .B(n_126), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_163), .B(n_128), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_150), .A2(n_139), .B1(n_123), .B2(n_128), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_149), .B(n_118), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_166), .B(n_123), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_166), .B(n_139), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_149), .B(n_98), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_152), .B(n_102), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_144), .B(n_81), .C(n_96), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_146), .B(n_136), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_142), .A2(n_122), .B(n_93), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_146), .B(n_127), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_143), .B(n_5), .Y(n_200) );
NOR2x1p5_ASAP7_75t_L g201 ( .A(n_143), .B(n_89), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_199), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_172), .B(n_164), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_197), .A2(n_148), .B(n_142), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_198), .A2(n_148), .B(n_162), .C(n_122), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_200), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_169), .A2(n_155), .B(n_152), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_174), .B(n_150), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_167), .B(n_155), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_167), .B(n_155), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_169), .A2(n_155), .B(n_159), .Y(n_211) );
AO22x1_ASAP7_75t_L g212 ( .A1(n_174), .A2(n_154), .B1(n_159), .B2(n_127), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_168), .Y(n_213) );
BUFx4f_ASAP7_75t_SL g214 ( .A(n_183), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_170), .B(n_162), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_168), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_168), .A2(n_150), .B1(n_154), .B2(n_159), .Y(n_217) );
NOR2xp67_ASAP7_75t_SL g218 ( .A(n_195), .B(n_103), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_180), .A2(n_150), .B(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_200), .B(n_150), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_168), .A2(n_84), .B1(n_94), .B2(n_154), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_175), .B(n_95), .Y(n_223) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_191), .A2(n_165), .B(n_161), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_107), .B(n_154), .C(n_160), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_171), .A2(n_165), .B(n_161), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_194), .B(n_177), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_175), .B(n_95), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_175), .B(n_95), .Y(n_229) );
BUFx8_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_199), .B(n_154), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_171), .A2(n_161), .B(n_160), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_201), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_199), .B(n_154), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_201), .B(n_154), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_204), .A2(n_175), .B(n_185), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_219), .A2(n_178), .B(n_173), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_206), .B(n_196), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_220), .A2(n_176), .B(n_186), .C(n_181), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_205), .A2(n_175), .B(n_178), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_203), .A2(n_193), .B(n_191), .C(n_188), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_230), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_224), .A2(n_193), .B(n_173), .Y(n_244) );
AOI221xp5_ASAP7_75t_SL g245 ( .A1(n_225), .A2(n_187), .B1(n_190), .B2(n_189), .C(n_184), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g246 ( .A(n_234), .B(n_170), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_230), .Y(n_247) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_226), .A2(n_182), .B(n_190), .Y(n_248) );
AO32x2_ASAP7_75t_L g249 ( .A1(n_222), .A2(n_179), .A3(n_124), .B1(n_133), .B2(n_125), .Y(n_249) );
AO31x2_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_189), .A3(n_145), .B(n_160), .Y(n_250) );
OAI22x1_ASAP7_75t_L g251 ( .A1(n_208), .A2(n_179), .B1(n_7), .B2(n_8), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_203), .B(n_182), .Y(n_252) );
CKINVDCx11_ASAP7_75t_R g253 ( .A(n_213), .Y(n_253) );
INVx8_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_233), .A2(n_182), .B(n_145), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_215), .B(n_154), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_231), .A2(n_195), .B(n_145), .Y(n_258) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_217), .A2(n_211), .B(n_207), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_212), .B(n_195), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_235), .A2(n_195), .B(n_156), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_227), .A2(n_195), .B(n_156), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_223), .A2(n_35), .B(n_59), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_202), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
AO31x2_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_210), .A3(n_209), .B(n_236), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_264), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_257), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_265), .B(n_216), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_239), .B(n_210), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_253), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_257), .B(n_209), .Y(n_272) );
AOI21xp33_ASAP7_75t_SL g273 ( .A1(n_251), .A2(n_229), .B(n_228), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_264), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_254), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_256), .B(n_221), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_246), .B(n_214), .Y(n_279) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_238), .A2(n_133), .B(n_125), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_243), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_259), .B(n_37), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_252), .B(n_214), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_242), .A2(n_218), .B(n_133), .C(n_125), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_240), .A2(n_6), .B(n_9), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_245), .A2(n_6), .B(n_10), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_248), .A2(n_133), .B(n_125), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_237), .A2(n_124), .B(n_125), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_247), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_275), .Y(n_290) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_286), .A2(n_260), .B(n_244), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_277), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_270), .B(n_253), .Y(n_293) );
AOI21x1_ASAP7_75t_L g294 ( .A1(n_287), .A2(n_262), .B(n_255), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_276), .A2(n_255), .B(n_263), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_276), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_281), .B(n_254), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_287), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_287), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_282), .B(n_254), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_277), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_282), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_267), .B(n_250), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_287), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_267), .B(n_249), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_285), .A2(n_261), .B(n_258), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_268), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_274), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_271), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_289), .B(n_254), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_302), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_304), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_304), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_309), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_290), .B(n_275), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_309), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_308), .B(n_272), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_299), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_290), .B(n_282), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_312), .B(n_282), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_303), .B(n_266), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_306), .B(n_266), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_293), .B(n_271), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_306), .B(n_266), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_301), .B(n_266), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_301), .B(n_303), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_301), .B(n_266), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_299), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_301), .B(n_266), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_300), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_297), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_332), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_317), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_335), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_332), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_325), .B(n_305), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_332), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_325), .B(n_305), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_297), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_305), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_331), .A2(n_310), .B1(n_259), .B2(n_298), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_327), .B(n_295), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_339), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_335), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_327), .B(n_295), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_331), .B(n_295), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_339), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_315), .B(n_295), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_315), .B(n_273), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_328), .B(n_291), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_328), .B(n_291), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_328), .B(n_291), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_329), .B(n_302), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_320), .B(n_302), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_328), .B(n_249), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_329), .B(n_294), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_322), .B(n_249), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_316), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_324), .B(n_292), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_322), .B(n_249), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_330), .B(n_280), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_324), .B(n_292), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_318), .B(n_273), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_337), .B(n_280), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_326), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_323), .B(n_311), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_334), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_366), .B(n_334), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_347), .B(n_338), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_344), .Y(n_390) );
AND2x2_ASAP7_75t_SL g391 ( .A(n_345), .B(n_330), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_350), .B(n_323), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_350), .B(n_321), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_355), .B(n_358), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_355), .B(n_321), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_376), .B(n_316), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_373), .B(n_341), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_349), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_349), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_354), .B(n_341), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_354), .B(n_340), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_340), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_359), .B(n_337), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_385), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_367), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_359), .B(n_342), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_372), .B(n_313), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_313), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_379), .B(n_280), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_379), .B(n_294), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_365), .B(n_307), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_343), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_343), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_376), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_371), .B(n_10), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_365), .B(n_288), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_386), .B(n_279), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_363), .B(n_11), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_368), .B(n_288), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_357), .B(n_250), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_368), .B(n_133), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_382), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_357), .A2(n_277), .B1(n_269), .B2(n_283), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_382), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_380), .B(n_250), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_380), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_369), .B(n_250), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_351), .B(n_12), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_351), .B(n_12), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_369), .B(n_124), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_361), .B(n_124), .Y(n_439) );
INVx3_ASAP7_75t_SL g440 ( .A(n_391), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_394), .B(n_361), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_416), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_404), .B(n_363), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_395), .B(n_352), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_405), .B(n_381), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_390), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_395), .B(n_352), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_404), .B(n_381), .Y(n_453) );
INVxp33_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_394), .B(n_373), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_387), .B(n_373), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_420), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_418), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_417), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_403), .B(n_353), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_387), .B(n_374), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_436), .A2(n_370), .B1(n_383), .B2(n_375), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_403), .B(n_434), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_391), .A2(n_383), .B1(n_356), .B2(n_343), .Y(n_466) );
NAND2x1p5_ASAP7_75t_L g467 ( .A(n_436), .B(n_277), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_415), .B(n_374), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g471 ( .A1(n_397), .A2(n_378), .B(n_277), .C(n_384), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_415), .B(n_378), .Y(n_472) );
AOI21xp33_ASAP7_75t_L g473 ( .A1(n_425), .A2(n_384), .B(n_364), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_392), .B(n_364), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_389), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_424), .A2(n_346), .B1(n_360), .B2(n_356), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_409), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_389), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_393), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_392), .B(n_360), .Y(n_482) );
OAI32xp33_ASAP7_75t_L g483 ( .A1(n_437), .A2(n_360), .A3(n_356), .B1(n_348), .B2(n_346), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_414), .B(n_348), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_430), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_461), .B(n_439), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_447), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g489 ( .A(n_442), .B(n_437), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_449), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_449), .B(n_393), .Y(n_491) );
NAND2x1_ASAP7_75t_L g492 ( .A(n_479), .B(n_411), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_448), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_463), .A2(n_431), .B(n_438), .Y(n_494) );
O2A1O1Ixp5_ASAP7_75t_L g495 ( .A1(n_454), .A2(n_411), .B(n_422), .C(n_429), .Y(n_495) );
AOI32xp33_ASAP7_75t_L g496 ( .A1(n_454), .A2(n_411), .A3(n_409), .B1(n_429), .B2(n_439), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_450), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_444), .B(n_388), .Y(n_498) );
OAI21xp33_ASAP7_75t_SL g499 ( .A1(n_455), .A2(n_388), .B(n_433), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_441), .B(n_414), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g501 ( .A(n_473), .B(n_427), .C(n_433), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_477), .B(n_480), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_451), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_458), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_440), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_445), .B(n_410), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_481), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_440), .A2(n_410), .B1(n_412), .B2(n_435), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_455), .B(n_412), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_456), .B(n_435), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_445), .A2(n_426), .B1(n_423), .B2(n_413), .Y(n_511) );
OAI322xp33_ASAP7_75t_L g512 ( .A1(n_463), .A2(n_427), .A3(n_396), .B1(n_432), .B2(n_401), .C1(n_402), .C2(n_423), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_467), .A2(n_426), .B(n_413), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_477), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_375), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_483), .A2(n_13), .B(n_14), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_505), .A2(n_466), .B(n_467), .C(n_471), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_505), .A2(n_464), .B1(n_480), .B2(n_478), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_512), .A2(n_443), .B1(n_453), .B2(n_470), .C(n_457), .Y(n_519) );
NOR2x1_ASAP7_75t_L g520 ( .A(n_492), .B(n_441), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_490), .Y(n_521) );
AOI21xp33_ASAP7_75t_L g522 ( .A1(n_504), .A2(n_485), .B(n_459), .Y(n_522) );
OA33x2_ASAP7_75t_L g523 ( .A1(n_487), .A2(n_469), .A3(n_472), .B1(n_482), .B2(n_476), .B3(n_484), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_498), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_499), .A2(n_484), .B1(n_481), .B2(n_475), .Y(n_525) );
NAND5xp2_ASAP7_75t_L g526 ( .A(n_494), .B(n_284), .C(n_269), .D(n_452), .E(n_462), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_495), .B(n_474), .C(n_468), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_501), .A2(n_462), .B1(n_468), .B2(n_465), .C(n_474), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_486), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_504), .B(n_465), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_513), .A2(n_460), .B1(n_278), .B2(n_263), .C1(n_13), .C2(n_14), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_488), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_491), .Y(n_533) );
OAI222xp33_ASAP7_75t_L g534 ( .A1(n_496), .A2(n_15), .B1(n_16), .B2(n_18), .C1(n_19), .C2(n_20), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_506), .A2(n_511), .B(n_508), .C(n_516), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_489), .A2(n_30), .B(n_32), .C(n_33), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_500), .B(n_34), .C(n_45), .D(n_48), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_489), .A2(n_156), .B1(n_51), .B2(n_55), .C(n_56), .Y(n_538) );
AOI21xp33_ASAP7_75t_SL g539 ( .A1(n_507), .A2(n_50), .B(n_57), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_493), .B(n_62), .C(n_65), .D(n_66), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_497), .A2(n_68), .B(n_69), .C(n_76), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_503), .A2(n_156), .B1(n_514), .B2(n_510), .C(n_515), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_502), .A2(n_156), .B1(n_499), .B2(n_505), .C(n_496), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_533), .B(n_520), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_540), .B(n_543), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_532), .B(n_521), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_529), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g548 ( .A(n_531), .B(n_526), .C(n_535), .D(n_536), .Y(n_548) );
NAND4xp75_ASAP7_75t_L g549 ( .A(n_545), .B(n_519), .C(n_542), .D(n_525), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_544), .B(n_517), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_547), .B(n_524), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_551), .Y(n_552) );
NAND4xp25_ASAP7_75t_SL g553 ( .A(n_550), .B(n_517), .C(n_528), .D(n_548), .Y(n_553) );
AO22x2_ASAP7_75t_L g554 ( .A1(n_552), .A2(n_549), .B1(n_527), .B2(n_546), .Y(n_554) );
XOR2xp5_ASAP7_75t_L g555 ( .A(n_553), .B(n_537), .Y(n_555) );
XNOR2x1_ASAP7_75t_L g556 ( .A(n_555), .B(n_518), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_556), .Y(n_557) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_557), .A2(n_554), .B(n_541), .Y(n_558) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_558), .A2(n_522), .B(n_534), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_559), .A2(n_530), .B1(n_538), .B2(n_539), .Y(n_560) );
AOI21xp33_ASAP7_75t_SL g561 ( .A1(n_560), .A2(n_523), .B(n_509), .Y(n_561) );
endmodule