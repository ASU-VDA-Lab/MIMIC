module fake_jpeg_29082_n_428 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_428);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_428;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_34),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_76),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_86),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_87),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_84),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_44),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_61),
.Y(n_102)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx6p67_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_121),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_47),
.B1(n_39),
.B2(n_42),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_49),
.B1(n_51),
.B2(n_77),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_20),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_59),
.A2(n_41),
.B1(n_32),
.B2(n_37),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_67),
.B1(n_80),
.B2(n_79),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_53),
.B(n_37),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_41),
.B1(n_20),
.B2(n_32),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_43),
.B1(n_44),
.B2(n_35),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_84),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_60),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_136),
.Y(n_184)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_139),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_162),
.B1(n_128),
.B2(n_103),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_43),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_164),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_167),
.B1(n_83),
.B2(n_107),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_R g148 ( 
.A(n_127),
.B(n_77),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_157),
.Y(n_175)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_156),
.Y(n_176)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_158),
.B1(n_160),
.B2(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_96),
.A2(n_89),
.B1(n_101),
.B2(n_103),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_145),
.B1(n_141),
.B2(n_126),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_105),
.B(n_39),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_105),
.B(n_42),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_173),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_114),
.C(n_100),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_126),
.B1(n_119),
.B2(n_89),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_177),
.B1(n_183),
.B2(n_102),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_96),
.B1(n_68),
.B2(n_69),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_188),
.B1(n_193),
.B2(n_145),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_116),
.C(n_100),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_190),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_91),
.B1(n_85),
.B2(n_73),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_40),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_91),
.B1(n_115),
.B2(n_55),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_70),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_143),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_202),
.B1(n_193),
.B2(n_180),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_214),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_115),
.B1(n_149),
.B2(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_145),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_216),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_47),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_153),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_10),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_153),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_217),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_157),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_182),
.B(n_9),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_194),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_173),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_224),
.B(n_202),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_180),
.B1(n_165),
.B2(n_177),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_228),
.A2(n_238),
.B1(n_240),
.B2(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_202),
.B1(n_200),
.B2(n_216),
.Y(n_265)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_175),
.A3(n_181),
.B1(n_186),
.B2(n_191),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_175),
.C(n_191),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_221),
.C(n_212),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_236),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_219),
.Y(n_237)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_179),
.B1(n_50),
.B2(n_192),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_181),
.B1(n_140),
.B2(n_186),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_151),
.B(n_170),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_216),
.B(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_192),
.B1(n_108),
.B2(n_117),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_229),
.Y(n_246)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_201),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_247),
.B(n_253),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_234),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_256),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_249),
.A2(n_265),
.B1(n_225),
.B2(n_245),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_216),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_213),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_209),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_254),
.B(n_255),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_222),
.B(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_215),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_264),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_222),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_262),
.C(n_271),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_212),
.C(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_225),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_235),
.Y(n_278)
);

INVx6_ASAP7_75t_SL g269 ( 
.A(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_226),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_218),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_206),
.C(n_203),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_231),
.B1(n_225),
.B2(n_240),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_265),
.B1(n_238),
.B2(n_250),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_300),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_233),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_292),
.C(n_244),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_227),
.C(n_223),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_301),
.Y(n_308)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_263),
.B1(n_267),
.B2(n_252),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_227),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_223),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_298),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_295),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_226),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_242),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_230),
.Y(n_299)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_262),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_246),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_268),
.B1(n_264),
.B2(n_259),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_303),
.A2(n_316),
.B1(n_172),
.B2(n_106),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_315),
.B1(n_317),
.B2(n_322),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_307),
.B(n_293),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_311),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_250),
.C(n_251),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_321),
.C(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_323),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_276),
.A2(n_228),
.B1(n_263),
.B2(n_267),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_267),
.B1(n_273),
.B2(n_200),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_242),
.B(n_241),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_288),
.B(n_295),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_285),
.A2(n_273),
.B1(n_239),
.B2(n_198),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_286),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_198),
.C(n_170),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_337),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_278),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_330),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_300),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_331),
.A2(n_155),
.B(n_104),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_288),
.B(n_280),
.C(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_335),
.C(n_340),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_290),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_303),
.A2(n_280),
.B1(n_289),
.B2(n_283),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_336),
.A2(n_346),
.B1(n_155),
.B2(n_158),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_308),
.B(n_279),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_282),
.C(n_275),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_313),
.B(n_274),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_310),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_282),
.B1(n_274),
.B2(n_205),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_205),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_345),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_324),
.B(n_10),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_312),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_317),
.C(n_322),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_135),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_348),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_315),
.B(n_318),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_351),
.A2(n_356),
.B(n_342),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_355),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_336),
.B(n_338),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_172),
.C(n_152),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_365),
.C(n_135),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_361),
.A2(n_346),
.B1(n_332),
.B2(n_327),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_340),
.B(n_19),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_7),
.Y(n_376)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_335),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_135),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_125),
.C(n_40),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_367),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_372),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_347),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_349),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_334),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_373),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_376),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_333),
.B1(n_330),
.B2(n_328),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_379),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_381),
.Y(n_389)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_364),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_356),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_390),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_371),
.A2(n_353),
.B(n_360),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_391),
.B(n_12),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_368),
.A2(n_366),
.B(n_365),
.Y(n_391)
);

AND2x2_ASAP7_75t_SL g392 ( 
.A(n_369),
.B(n_361),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_392),
.B(n_370),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_367),
.B1(n_354),
.B2(n_378),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_395),
.B1(n_10),
.B2(n_13),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_370),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_402),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_109),
.C(n_94),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_400),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_385),
.A2(n_384),
.B(n_393),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_11),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_392),
.B(n_11),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_403),
.B(n_6),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_109),
.C(n_70),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_94),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_406),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_52),
.C(n_54),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_401),
.A2(n_7),
.B1(n_6),
.B2(n_5),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_5),
.C(n_1),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_411),
.B(n_412),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_407),
.A2(n_399),
.B(n_403),
.Y(n_413)
);

AOI322xp5_ASAP7_75t_L g422 ( 
.A1(n_413),
.A2(n_416),
.A3(n_52),
.B1(n_54),
.B2(n_58),
.C1(n_0),
.C2(n_2),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_SL g416 ( 
.A1(n_408),
.A2(n_5),
.B(n_4),
.C(n_134),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_0),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_411),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_415),
.C(n_58),
.Y(n_423)
);

OAI321xp33_ASAP7_75t_L g424 ( 
.A1(n_420),
.A2(n_421),
.A3(n_422),
.B1(n_2),
.B2(n_3),
.C(n_30),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_414),
.B(n_0),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_423),
.A2(n_424),
.B1(n_2),
.B2(n_3),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_2),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_30),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_427),
.A2(n_30),
.B(n_102),
.Y(n_428)
);


endmodule