module real_aes_6337_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g173 ( .A1(n_0), .A2(n_174), .B(n_175), .C(n_179), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_1), .B(n_169), .Y(n_180) );
INVx1_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_3), .B(n_134), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_4), .A2(n_115), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_5), .A2(n_120), .B(n_125), .C(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_6), .A2(n_115), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_7), .B(n_169), .Y(n_456) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_8), .A2(n_148), .B(n_198), .Y(n_197) );
AND2x6_ASAP7_75t_L g120 ( .A(n_9), .B(n_121), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_10), .A2(n_120), .B(n_125), .C(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g511 ( .A(n_11), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_12), .B(n_40), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_13), .B(n_178), .Y(n_488) );
INVx1_ASAP7_75t_L g144 ( .A(n_14), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_15), .B(n_134), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_135), .B(n_496), .C(n_498), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_17), .B(n_169), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_18), .B(n_162), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_19), .A2(n_125), .B(n_156), .C(n_161), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_20), .A2(n_177), .B(n_192), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_21), .B(n_178), .Y(n_441) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_22), .A2(n_100), .B1(n_704), .B2(n_705), .C1(n_711), .C2(n_716), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_22), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_23), .B(n_178), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_24), .Y(n_437) );
INVx1_ASAP7_75t_L g462 ( .A(n_25), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_26), .A2(n_125), .B(n_161), .C(n_201), .Y(n_200) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_27), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_28), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_29), .Y(n_716) );
INVx1_ASAP7_75t_L g538 ( .A(n_30), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_31), .A2(n_115), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g118 ( .A(n_32), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_33), .A2(n_123), .B(n_128), .C(n_138), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_34), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_35), .A2(n_177), .B(n_453), .C(n_455), .Y(n_452) );
INVxp67_ASAP7_75t_L g539 ( .A(n_36), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_37), .B(n_203), .Y(n_202) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_38), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_39), .A2(n_125), .B(n_161), .C(n_461), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_41), .A2(n_179), .B(n_509), .C(n_510), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_42), .B(n_154), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_43), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_44), .B(n_134), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_45), .B(n_115), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_46), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_47), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_48), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_49), .A2(n_123), .B(n_138), .C(n_212), .Y(n_211) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_50), .A2(n_99), .B1(n_717), .B2(n_726), .C1(n_733), .C2(n_739), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_50), .A2(n_106), .B1(n_107), .B2(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_50), .Y(n_729) );
INVx1_ASAP7_75t_L g176 ( .A(n_51), .Y(n_176) );
INVx1_ASAP7_75t_L g213 ( .A(n_52), .Y(n_213) );
INVx1_ASAP7_75t_L g474 ( .A(n_53), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_54), .B(n_115), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_55), .Y(n_165) );
CKINVDCx14_ASAP7_75t_R g507 ( .A(n_56), .Y(n_507) );
INVx1_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_58), .B(n_115), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_59), .B(n_169), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_60), .A2(n_160), .B(n_223), .C(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g143 ( .A(n_61), .Y(n_143) );
INVx1_ASAP7_75t_SL g454 ( .A(n_62), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_63), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_64), .B(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_65), .B(n_169), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_66), .B(n_135), .Y(n_189) );
INVx1_ASAP7_75t_L g440 ( .A(n_67), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_68), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_69), .B(n_131), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_70), .A2(n_125), .B(n_138), .C(n_249), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g221 ( .A(n_71), .Y(n_221) );
INVx1_ASAP7_75t_L g721 ( .A(n_72), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_73), .A2(n_115), .B(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_74), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_75), .A2(n_115), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_76), .A2(n_154), .B(n_534), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_77), .Y(n_459) );
INVx1_ASAP7_75t_L g494 ( .A(n_78), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_79), .B(n_130), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_80), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_81), .A2(n_115), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g497 ( .A(n_82), .Y(n_497) );
INVx2_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
INVx1_ASAP7_75t_L g487 ( .A(n_84), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_85), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_86), .B(n_178), .Y(n_190) );
OR2x2_ASAP7_75t_L g102 ( .A(n_87), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g427 ( .A(n_87), .Y(n_427) );
OR2x2_ASAP7_75t_L g725 ( .A(n_87), .B(n_715), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_88), .A2(n_125), .B(n_138), .C(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_89), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
INVxp67_ASAP7_75t_L g226 ( .A(n_91), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_92), .B(n_148), .Y(n_512) );
INVx1_ASAP7_75t_L g185 ( .A(n_93), .Y(n_185) );
INVx1_ASAP7_75t_L g250 ( .A(n_94), .Y(n_250) );
INVx2_ASAP7_75t_L g477 ( .A(n_95), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_96), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g215 ( .A(n_97), .B(n_140), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_106), .B1(n_425), .B2(n_428), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g708 ( .A(n_102), .Y(n_708) );
OR2x2_ASAP7_75t_L g426 ( .A(n_103), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g715 ( .A(n_103), .Y(n_715) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_107), .A2(n_706), .B1(n_709), .B2(n_710), .Y(n_705) );
OR3x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_339), .C(n_382), .Y(n_107) );
NAND5xp2_ASAP7_75t_L g108 ( .A(n_109), .B(n_266), .C(n_296), .D(n_313), .E(n_328), .Y(n_108) );
AOI221xp5_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_181), .B1(n_228), .B2(n_234), .C(n_238), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_150), .Y(n_110) );
OR2x2_ASAP7_75t_L g243 ( .A(n_111), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g283 ( .A(n_111), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g301 ( .A(n_111), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_111), .B(n_236), .Y(n_318) );
OR2x2_ASAP7_75t_L g330 ( .A(n_111), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_111), .B(n_289), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_111), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_111), .B(n_267), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_111), .B(n_275), .Y(n_381) );
AND2x2_ASAP7_75t_L g413 ( .A(n_111), .B(n_167), .Y(n_413) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_111), .Y(n_421) );
INVx5_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_112), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g240 ( .A(n_112), .B(n_216), .Y(n_240) );
BUFx2_ASAP7_75t_L g263 ( .A(n_112), .Y(n_263) );
AND2x2_ASAP7_75t_L g292 ( .A(n_112), .B(n_151), .Y(n_292) );
AND2x2_ASAP7_75t_L g347 ( .A(n_112), .B(n_244), .Y(n_347) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_145), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_122), .B(n_140), .Y(n_113) );
BUFx2_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_116), .B(n_120), .Y(n_186) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx1_ASAP7_75t_L g160 ( .A(n_117), .Y(n_160) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g126 ( .A(n_118), .Y(n_126) );
INVx1_ASAP7_75t_L g193 ( .A(n_118), .Y(n_193) );
INVx1_ASAP7_75t_L g127 ( .A(n_119), .Y(n_127) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_119), .Y(n_132) );
INVx3_ASAP7_75t_L g135 ( .A(n_119), .Y(n_135) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_119), .Y(n_178) );
INVx1_ASAP7_75t_L g203 ( .A(n_119), .Y(n_203) );
INVx4_ASAP7_75t_SL g139 ( .A(n_120), .Y(n_139) );
BUFx3_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_124), .A2(n_139), .B(n_172), .C(n_173), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_124), .A2(n_139), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_124), .A2(n_139), .B(n_451), .C(n_452), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_124), .A2(n_139), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_124), .A2(n_139), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_124), .A2(n_139), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_124), .A2(n_139), .B(n_535), .C(n_536), .Y(n_534) );
INVx5_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
BUFx3_ASAP7_75t_L g137 ( .A(n_126), .Y(n_137) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_126), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_133), .C(n_136), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_130), .A2(n_136), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_130), .A2(n_440), .B(n_441), .C(n_442), .Y(n_439) );
O2A1O1Ixp5_ASAP7_75t_L g486 ( .A1(n_130), .A2(n_442), .B(n_487), .C(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g224 ( .A(n_132), .Y(n_224) );
INVx2_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_134), .B(n_226), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_134), .A2(n_159), .B(n_462), .C(n_463), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_134), .A2(n_224), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_135), .B(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
INVx1_ASAP7_75t_L g498 ( .A(n_137), .Y(n_498) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
INVx1_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_140), .A2(n_210), .B(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_140), .A2(n_186), .B(n_459), .C(n_460), .Y(n_458) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_140), .A2(n_505), .B(n_512), .Y(n_504) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g149 ( .A(n_141), .B(n_142), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx3_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_147), .A2(n_184), .B(n_194), .Y(n_183) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_147), .A2(n_247), .B(n_255), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_147), .B(n_256), .Y(n_255) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_147), .A2(n_436), .B(n_443), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_147), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_147), .B(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_148), .A2(n_199), .B(n_200), .Y(n_198) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g196 ( .A(n_149), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_150), .B(n_301), .Y(n_310) );
OAI32xp33_ASAP7_75t_L g324 ( .A1(n_150), .A2(n_260), .A3(n_325), .B1(n_326), .B2(n_327), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_150), .B(n_326), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_150), .B(n_243), .Y(n_367) );
INVx1_ASAP7_75t_SL g396 ( .A(n_150), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g405 ( .A(n_150), .B(n_183), .C(n_347), .D(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_167), .Y(n_150) );
INVx5_ASAP7_75t_L g237 ( .A(n_151), .Y(n_237) );
AND2x2_ASAP7_75t_L g267 ( .A(n_151), .B(n_168), .Y(n_267) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_151), .Y(n_346) );
AND2x2_ASAP7_75t_L g416 ( .A(n_151), .B(n_363), .Y(n_416) );
OR2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_164), .Y(n_151) );
AOI21xp5_ASAP7_75t_SL g152 ( .A1(n_153), .A2(n_155), .B(n_162), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_159), .Y(n_156) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_160), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_163), .B(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_166), .A2(n_483), .B(n_489), .Y(n_482) );
AND2x4_ASAP7_75t_L g289 ( .A(n_167), .B(n_237), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_167), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g323 ( .A(n_167), .B(n_244), .Y(n_323) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g236 ( .A(n_168), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g275 ( .A(n_168), .B(n_246), .Y(n_275) );
AND2x2_ASAP7_75t_L g284 ( .A(n_168), .B(n_245), .Y(n_284) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_180), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_177), .B(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g509 ( .A(n_178), .Y(n_509) );
INVx2_ASAP7_75t_L g442 ( .A(n_179), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_181), .A2(n_353), .B1(n_355), .B2(n_357), .C1(n_360), .C2(n_361), .Y(n_352) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_205), .Y(n_181) );
AND2x2_ASAP7_75t_L g285 ( .A(n_182), .B(n_286), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_182), .B(n_263), .C(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_197), .Y(n_182) );
INVx5_ASAP7_75t_SL g233 ( .A(n_183), .Y(n_233) );
OAI322xp33_ASAP7_75t_L g238 ( .A1(n_183), .A2(n_239), .A3(n_241), .B1(n_242), .B2(n_257), .C1(n_260), .C2(n_262), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_183), .B(n_231), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_183), .B(n_217), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_186), .A2(n_437), .B(n_438), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_186), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_191), .A2(n_202), .B(n_204), .Y(n_201) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx2_ASAP7_75t_L g532 ( .A(n_196), .Y(n_532) );
INVx2_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_197), .B(n_207), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_205), .B(n_270), .Y(n_325) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g304 ( .A(n_206), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
OR2x2_ASAP7_75t_L g232 ( .A(n_207), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_207), .B(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g272 ( .A(n_207), .B(n_217), .Y(n_272) );
AND2x2_ASAP7_75t_L g295 ( .A(n_207), .B(n_231), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_207), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g311 ( .A(n_207), .B(n_270), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_207), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_207), .B(n_279), .Y(n_369) );
INVx5_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g259 ( .A(n_208), .B(n_233), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_208), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g286 ( .A(n_208), .B(n_217), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_208), .B(n_333), .Y(n_374) );
OR2x2_ASAP7_75t_L g390 ( .A(n_208), .B(n_334), .Y(n_390) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_208), .B(n_351), .Y(n_397) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_208), .Y(n_404) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_215), .Y(n_208) );
AND2x2_ASAP7_75t_L g258 ( .A(n_216), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g308 ( .A(n_216), .B(n_231), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_216), .B(n_233), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_216), .B(n_270), .Y(n_392) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_217), .B(n_233), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_217), .B(n_231), .Y(n_280) );
OR2x2_ASAP7_75t_L g334 ( .A(n_217), .B(n_231), .Y(n_334) );
AND2x2_ASAP7_75t_L g351 ( .A(n_217), .B(n_230), .Y(n_351) );
INVxp67_ASAP7_75t_L g373 ( .A(n_217), .Y(n_373) );
AND2x2_ASAP7_75t_L g400 ( .A(n_217), .B(n_270), .Y(n_400) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_217), .Y(n_407) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_217) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_218), .A2(n_449), .B(n_456), .Y(n_448) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_218), .A2(n_472), .B(n_478), .Y(n_471) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_218), .A2(n_492), .B(n_499), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_223), .A2(n_250), .B(n_251), .C(n_252), .Y(n_249) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_224), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_224), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_230), .B(n_281), .Y(n_354) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g270 ( .A(n_231), .B(n_233), .Y(n_270) );
OR2x2_ASAP7_75t_L g337 ( .A(n_231), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g281 ( .A(n_232), .Y(n_281) );
OR2x2_ASAP7_75t_L g342 ( .A(n_232), .B(n_334), .Y(n_342) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g241 ( .A(n_236), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_236), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g242 ( .A(n_237), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_237), .B(n_244), .Y(n_277) );
INVx2_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_237), .B(n_275), .Y(n_335) );
AND2x2_ASAP7_75t_L g360 ( .A(n_237), .B(n_284), .Y(n_360) );
INVx1_ASAP7_75t_L g312 ( .A(n_242), .Y(n_312) );
INVx2_ASAP7_75t_SL g299 ( .A(n_243), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_244), .Y(n_302) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_245), .Y(n_265) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx2_ASAP7_75t_L g363 ( .A(n_246), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_254), .Y(n_247) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g455 ( .A(n_253), .Y(n_455) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g332 ( .A(n_259), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g338 ( .A(n_259), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_259), .A2(n_341), .B1(n_343), .B2(n_348), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_259), .B(n_351), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_260), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g294 ( .A(n_261), .Y(n_294) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OR2x2_ASAP7_75t_L g276 ( .A(n_263), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_263), .B(n_267), .Y(n_327) );
AND2x2_ASAP7_75t_L g350 ( .A(n_263), .B(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g326 ( .A(n_265), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_273), .C(n_287), .Y(n_266) );
INVx1_ASAP7_75t_L g290 ( .A(n_267), .Y(n_290) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_267), .A2(n_399), .B1(n_401), .B2(n_402), .C(n_405), .Y(n_398) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g417 ( .A(n_270), .Y(n_417) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g366 ( .A(n_272), .B(n_305), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_278), .C(n_282), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OAI32xp33_ASAP7_75t_L g391 ( .A1(n_280), .A2(n_281), .A3(n_344), .B1(n_381), .B2(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g423 ( .A(n_283), .B(n_322), .Y(n_423) );
AND2x2_ASAP7_75t_L g370 ( .A(n_284), .B(n_322), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_284), .B(n_292), .Y(n_388) );
AOI31xp33_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_290), .A3(n_291), .B(n_293), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_289), .B(n_301), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_289), .B(n_299), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_289), .A2(n_319), .B1(n_409), .B2(n_412), .C(n_414), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g314 ( .A(n_294), .B(n_315), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_303), .B1(n_306), .B2(n_309), .C1(n_311), .C2(n_312), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g379 ( .A(n_298), .Y(n_379) );
INVx1_ASAP7_75t_L g401 ( .A(n_301), .Y(n_401) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_304), .A2(n_415), .B1(n_417), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g320 ( .A(n_305), .Y(n_320) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B1(n_319), .B2(n_321), .C(n_324), .Y(n_313) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g410 ( .A(n_316), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx1_ASAP7_75t_L g331 ( .A(n_323), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_326), .B(n_413), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_335), .B2(n_336), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g422 ( .A(n_335), .Y(n_422) );
INVxp33_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_337), .B(n_381), .Y(n_380) );
OAI32xp33_ASAP7_75t_L g371 ( .A1(n_338), .A2(n_372), .A3(n_373), .B1(n_374), .B2(n_375), .Y(n_371) );
NAND4xp25_ASAP7_75t_L g339 ( .A(n_340), .B(n_352), .C(n_364), .D(n_376), .Y(n_339) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NAND2xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_347), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_358), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_361), .A2(n_377), .B1(n_394), .B2(n_397), .C(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g412 ( .A(n_363), .B(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_368), .B2(n_370), .C(n_371), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_373), .B(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_380), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_393), .C(n_408), .D(n_419), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_389), .C(n_391), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g424 ( .A(n_411), .Y(n_424) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B(n_424), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx6_ASAP7_75t_L g709 ( .A(n_426), .Y(n_709) );
NOR2x2_ASAP7_75t_L g714 ( .A(n_427), .B(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g710 ( .A(n_428), .Y(n_710) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_429), .B(n_659), .Y(n_428) );
NOR4xp25_ASAP7_75t_L g429 ( .A(n_430), .B(n_596), .C(n_630), .D(n_646), .Y(n_429) );
NAND4xp25_ASAP7_75t_SL g430 ( .A(n_431), .B(n_525), .C(n_560), .D(n_576), .Y(n_430) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_466), .B1(n_500), .B2(n_513), .C1(n_518), .C2(n_524), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI31xp33_ASAP7_75t_L g692 ( .A1(n_433), .A2(n_693), .A3(n_694), .B(n_696), .Y(n_692) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_445), .Y(n_433) );
AND2x2_ASAP7_75t_L g667 ( .A(n_434), .B(n_447), .Y(n_667) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g517 ( .A(n_435), .Y(n_517) );
AND2x2_ASAP7_75t_L g524 ( .A(n_435), .B(n_457), .Y(n_524) );
AND2x2_ASAP7_75t_L g581 ( .A(n_435), .B(n_448), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_445), .B(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_446), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_446), .B(n_528), .Y(n_571) );
AND2x2_ASAP7_75t_L g664 ( .A(n_446), .B(n_604), .Y(n_664) );
OAI321xp33_ASAP7_75t_L g698 ( .A1(n_446), .A2(n_517), .A3(n_671), .B1(n_699), .B2(n_701), .C(n_702), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_446), .B(n_503), .C(n_611), .D(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_457), .Y(n_446) );
AND2x2_ASAP7_75t_L g566 ( .A(n_447), .B(n_515), .Y(n_566) );
AND2x2_ASAP7_75t_L g585 ( .A(n_447), .B(n_517), .Y(n_585) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g516 ( .A(n_448), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g541 ( .A(n_448), .B(n_457), .Y(n_541) );
AND2x2_ASAP7_75t_L g627 ( .A(n_448), .B(n_515), .Y(n_627) );
INVx3_ASAP7_75t_SL g515 ( .A(n_457), .Y(n_515) );
AND2x2_ASAP7_75t_L g559 ( .A(n_457), .B(n_546), .Y(n_559) );
OR2x2_ASAP7_75t_L g592 ( .A(n_457), .B(n_517), .Y(n_592) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_457), .Y(n_599) );
AND2x2_ASAP7_75t_L g628 ( .A(n_457), .B(n_516), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_457), .B(n_601), .Y(n_643) );
AND2x2_ASAP7_75t_L g675 ( .A(n_457), .B(n_667), .Y(n_675) );
AND2x2_ASAP7_75t_L g684 ( .A(n_457), .B(n_529), .Y(n_684) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_464), .Y(n_457) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_479), .Y(n_467) );
INVx1_ASAP7_75t_SL g652 ( .A(n_468), .Y(n_652) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g520 ( .A(n_469), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g502 ( .A(n_470), .B(n_481), .Y(n_502) );
AND2x2_ASAP7_75t_L g588 ( .A(n_470), .B(n_504), .Y(n_588) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g558 ( .A(n_471), .B(n_491), .Y(n_558) );
OR2x2_ASAP7_75t_L g569 ( .A(n_471), .B(n_504), .Y(n_569) );
AND2x2_ASAP7_75t_L g595 ( .A(n_471), .B(n_504), .Y(n_595) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_471), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_479), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_479), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g568 ( .A(n_480), .B(n_569), .Y(n_568) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_480), .A2(n_558), .A3(n_564), .B1(n_595), .B2(n_645), .C1(n_655), .C2(n_657), .Y(n_654) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_481), .B(n_503), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_481), .B(n_504), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_481), .B(n_521), .Y(n_575) );
AND2x2_ASAP7_75t_L g629 ( .A(n_481), .B(n_595), .Y(n_629) );
INVx1_ASAP7_75t_L g633 ( .A(n_481), .Y(n_633) );
AND2x2_ASAP7_75t_L g645 ( .A(n_481), .B(n_491), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_481), .B(n_520), .Y(n_677) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g542 ( .A(n_482), .B(n_491), .Y(n_542) );
BUFx3_ASAP7_75t_L g556 ( .A(n_482), .Y(n_556) );
AND3x2_ASAP7_75t_L g638 ( .A(n_482), .B(n_618), .C(n_639), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_491), .B(n_502), .C(n_503), .Y(n_501) );
INVx1_ASAP7_75t_SL g521 ( .A(n_491), .Y(n_521) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_491), .Y(n_623) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g617 ( .A(n_502), .B(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g624 ( .A(n_502), .Y(n_624) );
AND2x2_ASAP7_75t_L g662 ( .A(n_503), .B(n_640), .Y(n_662) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx3_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
AND2x2_ASAP7_75t_L g618 ( .A(n_504), .B(n_521), .Y(n_618) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
OR2x2_ASAP7_75t_L g562 ( .A(n_515), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g681 ( .A(n_515), .B(n_581), .Y(n_681) );
AND2x2_ASAP7_75t_L g695 ( .A(n_515), .B(n_517), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_516), .B(n_529), .Y(n_636) );
AND2x2_ASAP7_75t_L g683 ( .A(n_516), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g546 ( .A(n_517), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g563 ( .A(n_517), .B(n_529), .Y(n_563) );
INVx1_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g604 ( .A(n_517), .B(n_529), .Y(n_604) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_519), .A2(n_647), .B1(n_651), .B2(n_653), .C(n_654), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_520), .B(n_522), .Y(n_519) );
AND2x2_ASAP7_75t_L g550 ( .A(n_520), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_523), .B(n_557), .Y(n_700) );
AOI322xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_542), .A3(n_543), .B1(n_544), .B2(n_550), .C1(n_552), .C2(n_559), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_541), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_528), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_528), .B(n_591), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_528), .A2(n_541), .B(n_615), .C(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_528), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_528), .B(n_585), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_528), .B(n_667), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_528), .B(n_695), .Y(n_694) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_529), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_529), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g656 ( .A(n_529), .B(n_543), .Y(n_656) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_533), .B(n_540), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_531), .A2(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g548 ( .A(n_533), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_540), .Y(n_549) );
INVx1_ASAP7_75t_L g631 ( .A(n_541), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g641 ( .A1(n_541), .A2(n_566), .A3(n_642), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_541), .B(n_547), .Y(n_693) );
INVx1_ASAP7_75t_SL g554 ( .A(n_542), .Y(n_554) );
AND2x2_ASAP7_75t_L g587 ( .A(n_542), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g668 ( .A(n_542), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g553 ( .A(n_543), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g578 ( .A(n_543), .Y(n_578) );
AND2x2_ASAP7_75t_L g605 ( .A(n_543), .B(n_558), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_543), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g697 ( .A(n_543), .B(n_645), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_545), .B(n_615), .Y(n_688) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g584 ( .A(n_547), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g602 ( .A(n_547), .Y(n_602) );
NAND2xp33_ASAP7_75t_SL g552 ( .A(n_553), .B(n_555), .Y(n_552) );
OAI211xp5_ASAP7_75t_SL g596 ( .A1(n_554), .A2(n_597), .B(n_603), .C(n_619), .Y(n_596) );
OR2x2_ASAP7_75t_L g671 ( .A(n_554), .B(n_652), .Y(n_671) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g608 ( .A(n_556), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_556), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g577 ( .A(n_558), .B(n_578), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B(n_567), .C(n_570), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g611 ( .A(n_563), .Y(n_611) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_566), .B(n_604), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_566), .Y(n_615) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g574 ( .A(n_569), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g607 ( .A(n_569), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g669 ( .A(n_569), .Y(n_669) );
AOI21xp33_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_572), .B(n_574), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_572), .A2(n_583), .B(n_586), .Y(n_582) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_579), .B(n_582), .C(n_589), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_577), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_580), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_SL g593 ( .A(n_581), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_583), .A2(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_588), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_SL g613 ( .A(n_588), .Y(n_613) );
AOI21xp33_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_593), .B(n_594), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g644 ( .A(n_595), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_601), .B(n_627), .Y(n_653) );
AND2x2_ASAP7_75t_L g666 ( .A(n_601), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g680 ( .A(n_601), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g690 ( .A(n_601), .B(n_628), .Y(n_690) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_606), .C(n_614), .Y(n_603) );
INVx1_ASAP7_75t_L g650 ( .A(n_604), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B1(n_610), .B2(n_612), .Y(n_606) );
OR2x2_ASAP7_75t_L g612 ( .A(n_608), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_608), .B(n_669), .Y(n_691) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g685 ( .A(n_618), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_625), .B1(n_628), .B2(n_629), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g703 ( .A(n_623), .Y(n_703) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g649 ( .A(n_627), .Y(n_649) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_632), .B(n_634), .C(n_641), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_649), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR5xp2_ASAP7_75t_L g659 ( .A(n_660), .B(n_678), .C(n_686), .D(n_692), .E(n_698), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B(n_665), .C(n_672), .Y(n_660) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_670), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_675), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B(n_685), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g701 ( .A(n_681), .Y(n_701) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_SL g738 ( .A(n_720), .Y(n_738) );
INVx1_ASAP7_75t_L g737 ( .A(n_722), .Y(n_737) );
OA21x2_ASAP7_75t_L g740 ( .A1(n_722), .A2(n_738), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_725), .Y(n_730) );
BUFx2_ASAP7_75t_L g741 ( .A(n_725), .Y(n_741) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B(n_731), .Y(n_727) );
NOR2xp33_ASAP7_75t_SL g731 ( .A(n_730), .B(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
endmodule