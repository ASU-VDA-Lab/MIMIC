module fake_jpeg_28530_n_518 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_518);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_518;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_65),
.Y(n_124)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_74),
.Y(n_153)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_48),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_95),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_9),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_18),
.C(n_49),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_19),
.B(n_9),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_45),
.Y(n_143)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_35),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_39),
.B1(n_18),
.B2(n_41),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_103),
.A2(n_109),
.B1(n_136),
.B2(n_138),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_39),
.B1(n_35),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_105),
.A2(n_107),
.B1(n_44),
.B2(n_28),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_52),
.A2(n_34),
.B1(n_23),
.B2(n_43),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_19),
.B1(n_37),
.B2(n_31),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_49),
.B1(n_37),
.B2(n_31),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_112),
.A2(n_113),
.B1(n_141),
.B2(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_24),
.B1(n_29),
.B2(n_18),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_56),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_40),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_63),
.A2(n_29),
.B1(n_24),
.B2(n_35),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_138),
.B1(n_91),
.B2(n_80),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_34),
.B1(n_28),
.B2(n_41),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_40),
.C(n_34),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_25),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_40),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_33),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_33),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_83),
.B(n_33),
.Y(n_156)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_163),
.A2(n_165),
.B1(n_171),
.B2(n_187),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_164),
.B(n_203),
.C(n_208),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_68),
.B1(n_69),
.B2(n_76),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_101),
.B(n_83),
.CI(n_28),
.CON(n_167),
.SN(n_167)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_167),
.B(n_178),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_25),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_105),
.A2(n_79),
.B1(n_71),
.B2(n_89),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_100),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_180),
.Y(n_224)
);

INVx5_ASAP7_75t_SL g174 ( 
.A(n_126),
.Y(n_174)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_25),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_44),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_100),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_120),
.A2(n_44),
.B1(n_97),
.B2(n_45),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_182),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_117),
.A2(n_45),
.B1(n_98),
.B2(n_2),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_103),
.B(n_45),
.Y(n_183)
);

NOR2x1_ASAP7_75t_R g245 ( 
.A(n_183),
.B(n_0),
.Y(n_245)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_10),
.B1(n_17),
.B2(n_2),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_108),
.B1(n_129),
.B2(n_122),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_127),
.B(n_11),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_198),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_194),
.Y(n_260)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_115),
.A2(n_45),
.B1(n_11),
.B2(n_3),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_45),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_128),
.B(n_7),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_110),
.B(n_7),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_206),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_140),
.A2(n_6),
.B(n_16),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_207),
.A2(n_14),
.B(n_16),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_126),
.B(n_0),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_6),
.B1(n_16),
.B2(n_3),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_118),
.B1(n_152),
.B2(n_155),
.Y(n_243)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_135),
.Y(n_212)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_6),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_217),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_106),
.A2(n_17),
.B1(n_6),
.B2(n_3),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_129),
.B1(n_122),
.B2(n_118),
.Y(n_240)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_157),
.B(n_106),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_108),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_240),
.B1(n_267),
.B2(n_163),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_162),
.B(n_124),
.C(n_135),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_237),
.B(n_5),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_238),
.B(n_245),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_170),
.A2(n_124),
.B1(n_125),
.B2(n_149),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_149),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_242),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_243),
.A2(n_212),
.B1(n_219),
.B2(n_5),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_184),
.B(n_12),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_266),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_256),
.A2(n_207),
.B(n_208),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_177),
.A2(n_14),
.B1(n_16),
.B2(n_4),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_218),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_210),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_267)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_272),
.A2(n_280),
.B1(n_293),
.B2(n_300),
.Y(n_336)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_183),
.B1(n_174),
.B2(n_209),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_275),
.A2(n_277),
.B1(n_286),
.B2(n_307),
.Y(n_346)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_276),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_183),
.B1(n_161),
.B2(n_213),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_224),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_291),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_162),
.B1(n_175),
.B2(n_178),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_279),
.A2(n_312),
.B1(n_263),
.B2(n_230),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_171),
.B1(n_162),
.B2(n_164),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_167),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_294),
.Y(n_320)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

AO21x2_ASAP7_75t_SL g285 ( 
.A1(n_245),
.A2(n_183),
.B(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_SL g286 ( 
.A(n_237),
.B(n_168),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_287),
.B(n_15),
.Y(n_353)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_226),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_251),
.A2(n_167),
.B1(n_179),
.B2(n_208),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_203),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_295),
.A2(n_303),
.B(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_179),
.C(n_169),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_298),
.C(n_236),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_233),
.C(n_227),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_240),
.A2(n_234),
.B1(n_223),
.B2(n_227),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_234),
.A2(n_227),
.B1(n_241),
.B2(n_258),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_302),
.B1(n_305),
.B2(n_306),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_256),
.A2(n_181),
.B1(n_186),
.B2(n_185),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_235),
.A2(n_220),
.B(n_189),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_304),
.B(n_308),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_225),
.A2(n_172),
.B1(n_215),
.B2(n_216),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_264),
.A2(n_199),
.B1(n_192),
.B2(n_200),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_230),
.A2(n_202),
.B1(n_196),
.B2(n_190),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_263),
.A2(n_182),
.B(n_201),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_265),
.A2(n_166),
.B(n_204),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_310),
.A2(n_270),
.B(n_229),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_195),
.B1(n_176),
.B2(n_217),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_311),
.A2(n_1),
.B1(n_15),
.B2(n_17),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_5),
.Y(n_331)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_274),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_259),
.B(n_265),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_328),
.B(n_347),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_318),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_268),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_323),
.B(n_353),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_268),
.B1(n_259),
.B2(n_248),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_248),
.B1(n_249),
.B2(n_231),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_285),
.A2(n_249),
.B1(n_231),
.B2(n_261),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_261),
.B(n_266),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_335),
.C(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_331),
.B(n_349),
.Y(n_357)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_257),
.C(n_269),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_257),
.C(n_269),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_291),
.B(n_232),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_339),
.B(n_276),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_285),
.A2(n_232),
.B1(n_236),
.B2(n_222),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_343),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_222),
.B1(n_229),
.B2(n_270),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_285),
.A2(n_222),
.B1(n_253),
.B2(n_252),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_352),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_252),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_272),
.A2(n_253),
.B1(n_1),
.B2(n_0),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_354),
.A2(n_312),
.B1(n_290),
.B2(n_289),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_280),
.B(n_1),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_293),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_360),
.C(n_364),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_321),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_358),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_303),
.C(n_289),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_320),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_289),
.C(n_287),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_370),
.C(n_378),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_366),
.A2(n_382),
.B1(n_385),
.B2(n_311),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_320),
.B(n_292),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_367),
.B(n_369),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_316),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_302),
.C(n_301),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_332),
.Y(n_373)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_322),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_376),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_310),
.C(n_296),
.Y(n_378)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_337),
.A2(n_290),
.B1(n_300),
.B2(n_314),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_384),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_337),
.A2(n_313),
.B1(n_304),
.B2(n_315),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_383),
.A2(n_318),
.B1(n_327),
.B2(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_345),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_322),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_386),
.B(n_389),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_340),
.B(n_288),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_388),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_282),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_324),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_391),
.A2(n_384),
.B1(n_375),
.B2(n_371),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_377),
.A2(n_341),
.B1(n_343),
.B2(n_348),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_392),
.A2(n_393),
.B1(n_394),
.B2(n_419),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_341),
.B1(n_346),
.B2(n_328),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_352),
.B1(n_347),
.B2(n_354),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_381),
.A2(n_355),
.B1(n_326),
.B2(n_325),
.Y(n_395)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_353),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_408),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_363),
.A2(n_370),
.B1(n_383),
.B2(n_374),
.Y(n_400)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_350),
.B(n_344),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_405),
.A2(n_406),
.B(n_410),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_368),
.A2(n_350),
.B(n_344),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_333),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_368),
.A2(n_365),
.B(n_378),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_333),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_417),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_324),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_366),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_308),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_374),
.A2(n_317),
.B(n_329),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_418),
.A2(n_357),
.B(n_351),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_371),
.A2(n_351),
.B1(n_329),
.B2(n_299),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_404),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_421),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_399),
.Y(n_421)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_402),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_360),
.C(n_356),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_431),
.C(n_440),
.Y(n_455)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_388),
.C(n_387),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_397),
.B(n_358),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_434),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_435),
.A2(n_394),
.B1(n_405),
.B2(n_415),
.Y(n_463)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_413),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_443),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_438),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_385),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_390),
.B(n_284),
.C(n_271),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_398),
.B(n_380),
.C(n_273),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_444),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_442),
.Y(n_446)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_306),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_426),
.A2(n_400),
.B1(n_391),
.B2(n_416),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_447),
.A2(n_451),
.B1(n_460),
.B2(n_461),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_439),
.A2(n_422),
.B1(n_424),
.B2(n_443),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_398),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_462),
.Y(n_466)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_410),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_463),
.Y(n_472)
);

AOI21xp33_ASAP7_75t_L g458 ( 
.A1(n_427),
.A2(n_406),
.B(n_416),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_429),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_422),
.A2(n_416),
.B1(n_395),
.B2(n_392),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_405),
.B1(n_418),
.B2(n_393),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_412),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_435),
.Y(n_465)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_465),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_411),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_468),
.Y(n_483)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_469),
.B(n_473),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_441),
.C(n_440),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_455),
.C(n_450),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_461),
.A2(n_430),
.B(n_442),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_457),
.B(n_460),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_446),
.A2(n_430),
.B(n_436),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_453),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_456),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_423),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_478),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_463),
.A2(n_444),
.B1(n_409),
.B2(n_417),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_476),
.A2(n_462),
.B1(n_409),
.B2(n_425),
.Y(n_493)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_479),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_431),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_433),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_493),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_450),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_485),
.C(n_478),
.Y(n_497)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_484),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_425),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_471),
.A2(n_459),
.B1(n_454),
.B2(n_415),
.Y(n_487)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_488),
.B(n_490),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_465),
.A2(n_447),
.B(n_428),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_R g496 ( 
.A(n_491),
.B(n_473),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_496),
.B(n_499),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_500),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_470),
.C(n_466),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_475),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_466),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_489),
.A2(n_486),
.B(n_483),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_494),
.B(n_490),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_503),
.A2(n_504),
.B(n_506),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_492),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_492),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_508),
.B(n_480),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_505),
.A2(n_501),
.B(n_502),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_509),
.A2(n_507),
.B(n_480),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_510),
.A2(n_505),
.B(n_488),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_512),
.A2(n_513),
.B(n_511),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_482),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_485),
.B(n_493),
.Y(n_516)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_476),
.C(n_361),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_299),
.B1(n_281),
.B2(n_15),
.Y(n_518)
);


endmodule