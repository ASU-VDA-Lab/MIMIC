module fake_jpeg_28415_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_79),
.B1(n_61),
.B2(n_71),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_88),
.B1(n_54),
.B2(n_52),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_69),
.B1(n_58),
.B2(n_59),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_55),
.B1(n_64),
.B2(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_69),
.B1(n_59),
.B2(n_51),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_72),
.B1(n_64),
.B2(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_71),
.B1(n_72),
.B2(n_62),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_102),
.B(n_107),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_62),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_2),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_93),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_79),
.C(n_70),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_49),
.C(n_53),
.Y(n_117)
);

NAND2x1_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_86),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_67),
.B1(n_66),
.B2(n_60),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_110),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_95),
.B1(n_100),
.B2(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_103),
.B1(n_108),
.B2(n_5),
.Y(n_132)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_118),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_107),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_111),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_21),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_3),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_102),
.C(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_132),
.B1(n_119),
.B2(n_122),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_8),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_118),
.B1(n_23),
.B2(n_24),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_130),
.A2(n_117),
.B1(n_18),
.B2(n_22),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_9),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_156),
.C(n_139),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_27),
.B(n_42),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_30),
.B(n_38),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_26),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_137),
.B1(n_138),
.B2(n_134),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_159),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_150),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_151),
.C(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_151),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_161),
.A3(n_147),
.B1(n_25),
.B2(n_33),
.C(n_14),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_17),
.B1(n_41),
.B2(n_35),
.Y(n_169)
);

OAI321xp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_15),
.A3(n_34),
.B1(n_28),
.B2(n_16),
.C(n_46),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_10),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_12),
.Y(n_172)
);


endmodule