module fake_jpeg_31895_n_401 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_401);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_30),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_40),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_40),
.B1(n_31),
.B2(n_33),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_45),
.B1(n_47),
.B2(n_44),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_49),
.B(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_36),
.B1(n_26),
.B2(n_20),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_25),
.B1(n_19),
.B2(n_18),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_25),
.B1(n_19),
.B2(n_39),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_27),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_52),
.B(n_27),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_39),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_160),
.B1(n_161),
.B2(n_94),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_65),
.C(n_54),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_163),
.C(n_164),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_149),
.B1(n_157),
.B2(n_114),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_93),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_93),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_140),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_90),
.B(n_11),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_152),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_96),
.A2(n_79),
.B1(n_76),
.B2(n_62),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_66),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_107),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_91),
.B(n_68),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_159),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_60),
.B1(n_58),
.B2(n_48),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_46),
.B1(n_69),
.B2(n_114),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_91),
.B(n_69),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_115),
.A2(n_89),
.B1(n_124),
.B2(n_86),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_0),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_106),
.B(n_8),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_120),
.B1(n_86),
.B2(n_119),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_94),
.B1(n_119),
.B2(n_100),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_103),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_138),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_185),
.B1(n_148),
.B2(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_204),
.B1(n_167),
.B2(n_175),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_141),
.B1(n_150),
.B2(n_138),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_200),
.B1(n_201),
.B2(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_141),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_195),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_199),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_183),
.B1(n_181),
.B2(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_134),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_159),
.B1(n_133),
.B2(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_100),
.B1(n_134),
.B2(n_116),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_169),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_146),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_167),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_163),
.B1(n_156),
.B2(n_121),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_116),
.B1(n_161),
.B2(n_144),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_171),
.B(n_174),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_217),
.B1(n_207),
.B2(n_223),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_205),
.A2(n_177),
.B1(n_179),
.B2(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_204),
.B1(n_187),
.B2(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_194),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_175),
.B1(n_181),
.B2(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_178),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_195),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_198),
.B1(n_178),
.B2(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_199),
.B(n_143),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_227),
.B1(n_242),
.B2(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_243),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_200),
.B1(n_201),
.B2(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_234),
.B1(n_237),
.B2(n_223),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_219),
.B(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_203),
.B1(n_196),
.B2(n_190),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_202),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_189),
.B1(n_192),
.B2(n_137),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_239),
.B1(n_235),
.B2(n_210),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_236),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_250),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_251),
.B1(n_225),
.B2(n_241),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_216),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_215),
.B1(n_211),
.B2(n_209),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_214),
.C(n_206),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_261),
.C(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_213),
.B(n_206),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_211),
.B(n_212),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_212),
.B(n_242),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_214),
.C(n_226),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_278),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_229),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_255),
.B(n_256),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_281),
.B1(n_244),
.B2(n_252),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_145),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_186),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_249),
.B1(n_182),
.B2(n_155),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_210),
.B1(n_220),
.B2(n_139),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_183),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_152),
.C(n_182),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_250),
.C(n_253),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_281),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_285),
.B(n_290),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_261),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_258),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_269),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_292),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_271),
.C(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_302),
.C(n_303),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_299),
.B1(n_285),
.B2(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_251),
.B1(n_260),
.B2(n_249),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_266),
.B1(n_264),
.B2(n_186),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_142),
.C(n_151),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_147),
.C(n_153),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.C(n_266),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_153),
.C(n_140),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_276),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_310),
.C(n_324),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_270),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_328),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_274),
.B(n_268),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_306),
.B(n_299),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_319),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_SL g316 ( 
.A(n_300),
.B(n_267),
.C(n_264),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_316),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_318),
.A2(n_294),
.B1(n_297),
.B2(n_298),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_288),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_322),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_186),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_118),
.C(n_125),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_186),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_327),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_169),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_122),
.B1(n_129),
.B2(n_97),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_333),
.A2(n_338),
.B1(n_337),
.B2(n_342),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_294),
.B1(n_298),
.B2(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_296),
.B1(n_129),
.B2(n_127),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_309),
.B(n_13),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_341),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_316),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_320),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_343),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_319),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_313),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_315),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_350),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_312),
.C(n_321),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_348),
.B(n_357),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_333),
.B(n_321),
.CI(n_310),
.CON(n_349),
.SN(n_349)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_349),
.B(n_162),
.Y(n_370)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_355),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_312),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_356),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_324),
.B(n_169),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_337),
.B(n_162),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_344),
.C(n_330),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_363),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_358),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_362),
.A2(n_98),
.B(n_8),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_344),
.C(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_348),
.B(n_345),
.Y(n_364)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_364),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_352),
.B(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_334),
.Y(n_368)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_347),
.B(n_127),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_370),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_349),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_373),
.B(n_375),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_162),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_98),
.C(n_56),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_162),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_377),
.A2(n_9),
.B(n_17),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_8),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_378),
.B(n_17),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_380),
.A2(n_360),
.B(n_362),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_382),
.A2(n_383),
.B(n_372),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_385),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_17),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_376),
.Y(n_391)
);

NOR3xp33_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_15),
.C(n_13),
.Y(n_387)
);

O2A1O1Ixp33_ASAP7_75t_SL g389 ( 
.A1(n_387),
.A2(n_6),
.B(n_15),
.C(n_3),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_388),
.A2(n_390),
.B(n_374),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_391),
.B(n_375),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_393),
.A2(n_394),
.B(n_395),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_392),
.A2(n_6),
.B(n_2),
.Y(n_395)
);

A2O1A1O1Ixp25_ASAP7_75t_L g396 ( 
.A1(n_394),
.A2(n_1),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_396)
);

A2O1A1O1Ixp25_ASAP7_75t_L g398 ( 
.A1(n_396),
.A2(n_5),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_397),
.C(n_4),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_399),
.A2(n_1),
.B(n_5),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g401 ( 
.A1(n_400),
.A2(n_1),
.B(n_5),
.Y(n_401)
);


endmodule