module fake_jpeg_20864_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_1),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_22),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_46),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_19),
.B1(n_12),
.B2(n_16),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_34),
.B1(n_12),
.B2(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_17),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_33),
.B(n_17),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_57),
.C(n_49),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_56),
.B1(n_37),
.B2(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_63),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_13),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_50),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_19),
.B1(n_11),
.B2(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_46),
.B1(n_37),
.B2(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_55),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_72),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_74),
.B(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

A2O1A1O1Ixp25_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_57),
.B(n_58),
.C(n_52),
.D(n_59),
.Y(n_76)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_82),
.B1(n_54),
.B2(n_60),
.C(n_73),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_56),
.B(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_65),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_53),
.C(n_62),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_54),
.C(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_63),
.B1(n_62),
.B2(n_49),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_89),
.A3(n_75),
.B1(n_18),
.B2(n_63),
.C1(n_69),
.C2(n_70),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_87),
.CI(n_88),
.CON(n_91),
.SN(n_91)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_18),
.Y(n_89)
);

OAI321xp33_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_76),
.A3(n_83),
.B1(n_75),
.B2(n_81),
.C(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_93),
.B1(n_84),
.B2(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_69),
.B1(n_71),
.B2(n_10),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_5),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_91),
.B(n_5),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_91),
.C(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_100),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_93),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_101),
.B(n_95),
.Y(n_104)
);


endmodule