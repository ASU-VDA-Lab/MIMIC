module fake_jpeg_5701_n_135 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_4),
.B(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_38),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_17),
.B1(n_22),
.B2(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_23),
.A2(n_14),
.B1(n_17),
.B2(n_11),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_15),
.B(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_49),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_45),
.B1(n_51),
.B2(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_37),
.B(n_40),
.C(n_35),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_17),
.C(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

XNOR2x1_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_36),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_64),
.C(n_48),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_43),
.B1(n_28),
.B2(n_29),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_63),
.B1(n_33),
.B2(n_54),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_41),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_52),
.B1(n_54),
.B2(n_33),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_65),
.B(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_49),
.Y(n_69)
);

OAI322xp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_30),
.A3(n_16),
.B1(n_19),
.B2(n_21),
.C1(n_35),
.C2(n_24),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_60),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_74),
.B(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_65),
.B(n_60),
.C(n_67),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_69),
.C(n_74),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_62),
.C(n_55),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_26),
.B1(n_62),
.B2(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_89),
.C(n_21),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_70),
.C(n_73),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_68),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_15),
.B(n_12),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_26),
.B1(n_16),
.B2(n_38),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_35),
.B(n_42),
.C(n_46),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_55),
.C(n_46),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_6),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_46),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_88),
.C(n_81),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_111),
.C(n_12),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_80),
.B1(n_82),
.B2(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_80),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_109),
.B(n_110),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_102),
.C(n_93),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_38),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_12),
.B1(n_11),
.B2(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_110),
.B1(n_42),
.B2(n_0),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_123),
.C(n_2),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_116),
.B(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_129),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_0),
.B(n_1),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_130),
.B(n_131),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_7),
.A3(n_9),
.B1(n_2),
.B2(n_4),
.C1(n_10),
.C2(n_8),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_10),
.C(n_8),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_121),
.C(n_122),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);


endmodule