module fake_jpeg_14298_n_175 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g68 ( 
.A(n_0),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_1),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_88),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_46),
.B(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_71),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_43),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_61),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_58),
.B1(n_44),
.B2(n_60),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_68),
.B1(n_44),
.B2(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_52),
.B1(n_67),
.B2(n_64),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_69),
.B1(n_51),
.B2(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_114),
.Y(n_130)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_109),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_102),
.B1(n_114),
.B2(n_116),
.Y(n_129)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_108),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_49),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_54),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_48),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_134),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_65),
.B1(n_51),
.B2(n_66),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_132),
.B1(n_133),
.B2(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_129),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_19),
.B(n_36),
.C(n_32),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_24),
.B(n_30),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_104),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_20),
.C(n_31),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_5),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_124),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_21),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_6),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_149),
.C(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_155),
.B1(n_148),
.B2(n_143),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_148),
.B1(n_137),
.B2(n_132),
.C(n_10),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_13),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_152),
.B(n_154),
.Y(n_163)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_131),
.B1(n_125),
.B2(n_130),
.C(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_164),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_167),
.A3(n_159),
.B1(n_156),
.B2(n_146),
.C(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_157),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_161),
.B(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_169),
.B(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_123),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_140),
.Y(n_175)
);


endmodule