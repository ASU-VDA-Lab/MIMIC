module real_aes_2133_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_0), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_1), .B(n_146), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_2), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_3), .B(n_130), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_4), .B(n_148), .Y(n_471) );
INVx1_ASAP7_75t_L g137 ( .A(n_5), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_6), .B(n_130), .Y(n_129) );
NAND2xp33_ASAP7_75t_SL g216 ( .A(n_7), .B(n_136), .Y(n_216) );
INVx1_ASAP7_75t_L g197 ( .A(n_8), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g794 ( .A(n_9), .Y(n_794) );
AND2x2_ASAP7_75t_L g124 ( .A(n_10), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g473 ( .A(n_11), .B(n_187), .Y(n_473) );
AND2x2_ASAP7_75t_L g481 ( .A(n_12), .B(n_213), .Y(n_481) );
INVx2_ASAP7_75t_L g126 ( .A(n_13), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_14), .B(n_148), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_15), .Y(n_113) );
AOI221x1_ASAP7_75t_L g210 ( .A1(n_16), .A2(n_139), .B1(n_211), .B2(n_213), .C(n_215), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_17), .B(n_130), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_18), .B(n_130), .Y(n_504) );
INVx1_ASAP7_75t_L g116 ( .A(n_19), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_20), .A2(n_88), .B1(n_130), .B2(n_198), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_21), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_22), .A2(n_139), .B(n_144), .Y(n_138) );
AOI221xp5_ASAP7_75t_SL g174 ( .A1(n_23), .A2(n_36), .B1(n_130), .B2(n_139), .C(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_24), .B(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g127 ( .A(n_25), .B(n_87), .Y(n_127) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_25), .A2(n_87), .B(n_126), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_26), .B(n_148), .Y(n_186) );
INVxp67_ASAP7_75t_L g209 ( .A(n_27), .Y(n_209) );
AND2x2_ASAP7_75t_L g170 ( .A(n_28), .B(n_160), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_29), .A2(n_139), .B(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_30), .A2(n_213), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_31), .B(n_148), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_32), .A2(n_139), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_33), .B(n_148), .Y(n_499) );
AND2x2_ASAP7_75t_L g136 ( .A(n_34), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g140 ( .A(n_34), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g205 ( .A(n_34), .Y(n_205) );
OR2x6_ASAP7_75t_L g114 ( .A(n_35), .B(n_115), .Y(n_114) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_35), .B(n_793), .C(n_795), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_37), .B(n_130), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_38), .A2(n_80), .B1(n_139), .B2(n_203), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_39), .B(n_148), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_40), .A2(n_104), .B1(n_755), .B2(n_758), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_41), .B(n_130), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_42), .A2(n_72), .B1(n_779), .B2(n_780), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_42), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_43), .B(n_146), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_44), .A2(n_139), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g228 ( .A(n_45), .B(n_160), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_46), .B(n_146), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_47), .B(n_160), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_48), .B(n_130), .Y(n_487) );
INVx1_ASAP7_75t_L g133 ( .A(n_49), .Y(n_133) );
INVx1_ASAP7_75t_L g143 ( .A(n_49), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_50), .B(n_148), .Y(n_479) );
AND2x2_ASAP7_75t_L g515 ( .A(n_51), .B(n_160), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_52), .B(n_130), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_53), .B(n_146), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_54), .B(n_146), .Y(n_498) );
AND2x2_ASAP7_75t_L g161 ( .A(n_55), .B(n_160), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_56), .B(n_130), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_57), .B(n_148), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_58), .B(n_130), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_59), .A2(n_139), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_60), .B(n_146), .Y(n_157) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_61), .B(n_125), .Y(n_189) );
AND2x2_ASAP7_75t_L g510 ( .A(n_62), .B(n_125), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_63), .A2(n_139), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_64), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_65), .B(n_187), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_66), .B(n_146), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_67), .B(n_146), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_68), .A2(n_91), .B1(n_139), .B2(n_203), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_69), .B(n_148), .Y(n_507) );
INVx1_ASAP7_75t_L g135 ( .A(n_70), .Y(n_135) );
INVx1_ASAP7_75t_L g141 ( .A(n_70), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_71), .B(n_146), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_72), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_73), .A2(n_139), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_74), .A2(n_139), .B(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_75), .A2(n_139), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g501 ( .A(n_76), .B(n_125), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_77), .B(n_160), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_78), .B(n_130), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_79), .A2(n_82), .B1(n_130), .B2(n_198), .Y(n_239) );
INVx1_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_83), .B(n_146), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_84), .B(n_146), .Y(n_177) );
AND2x2_ASAP7_75t_L g464 ( .A(n_85), .B(n_187), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_86), .A2(n_139), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_89), .B(n_148), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_90), .A2(n_139), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_92), .B(n_148), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_93), .A2(n_100), .B1(n_105), .B2(n_106), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_93), .Y(n_105) );
INVxp67_ASAP7_75t_L g212 ( .A(n_94), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_95), .B(n_130), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_96), .B(n_148), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_97), .A2(n_139), .B(n_184), .Y(n_183) );
BUFx2_ASAP7_75t_L g509 ( .A(n_98), .Y(n_509) );
BUFx2_ASAP7_75t_L g766 ( .A(n_99), .Y(n_766) );
BUFx2_ASAP7_75t_SL g775 ( .A(n_99), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_100), .Y(n_106) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_786), .B(n_796), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_762), .B(n_773), .Y(n_102) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_107), .B(n_754), .Y(n_103) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_118), .B1(n_451), .B2(n_750), .Y(n_108) );
OAI22x1_ASAP7_75t_L g755 ( .A1(n_109), .A2(n_752), .B1(n_756), .B2(n_757), .Y(n_755) );
CKINVDCx11_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
INVx3_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
AND2x6_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x6_ASAP7_75t_SL g752 ( .A(n_113), .B(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g761 ( .A(n_113), .B(n_114), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_113), .B(n_753), .Y(n_771) );
CKINVDCx16_ASAP7_75t_R g795 ( .A(n_113), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_114), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_116), .B(n_117), .Y(n_791) );
INVx4_ASAP7_75t_L g756 ( .A(n_118), .Y(n_756) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_118), .Y(n_781) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_362), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_284), .C(n_334), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_251), .Y(n_120) );
AOI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_171), .B1(n_190), .B2(n_233), .C(n_243), .Y(n_121) );
INVx1_ASAP7_75t_SL g333 ( .A(n_122), .Y(n_333) );
AND2x4_ASAP7_75t_SL g122 ( .A(n_123), .B(n_151), .Y(n_122) );
INVx2_ASAP7_75t_L g255 ( .A(n_123), .Y(n_255) );
OR2x2_ASAP7_75t_L g277 ( .A(n_123), .B(n_268), .Y(n_277) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_123), .Y(n_292) );
INVx5_ASAP7_75t_L g299 ( .A(n_123), .Y(n_299) );
AND2x4_ASAP7_75t_L g305 ( .A(n_123), .B(n_163), .Y(n_305) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_123), .B(n_235), .Y(n_308) );
OR2x2_ASAP7_75t_L g317 ( .A(n_123), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g324 ( .A(n_123), .B(n_152), .Y(n_324) );
AND2x2_ASAP7_75t_L g425 ( .A(n_123), .B(n_162), .Y(n_425) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_128), .Y(n_123) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_125), .Y(n_160) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x4_ASAP7_75t_L g150 ( .A(n_126), .B(n_127), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_138), .B(n_150), .Y(n_128) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
INVx1_ASAP7_75t_L g217 ( .A(n_131), .Y(n_217) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
AND2x6_ASAP7_75t_L g146 ( .A(n_132), .B(n_141), .Y(n_146) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g148 ( .A(n_134), .B(n_143), .Y(n_148) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx5_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
AND2x2_ASAP7_75t_L g142 ( .A(n_137), .B(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
BUFx3_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
INVx2_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
AND2x4_ASAP7_75t_L g203 ( .A(n_142), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g200 ( .A(n_143), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B(n_149), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_146), .B(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_149), .A2(n_156), .B(n_157), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_149), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_149), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_149), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_149), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_149), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_149), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_149), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_149), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_149), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_149), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_149), .A2(n_520), .B(n_521), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_150), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_150), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_150), .B(n_212), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g215 ( .A(n_150), .B(n_216), .C(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_150), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_150), .A2(n_517), .B(n_518), .Y(n_516) );
INVx3_ASAP7_75t_SL g276 ( .A(n_151), .Y(n_276) );
AND2x2_ASAP7_75t_L g320 ( .A(n_151), .B(n_235), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_151), .A2(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g361 ( .A(n_151), .B(n_299), .Y(n_361) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_162), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_152), .B(n_163), .Y(n_242) );
OR2x2_ASAP7_75t_L g246 ( .A(n_152), .B(n_163), .Y(n_246) );
INVx1_ASAP7_75t_L g254 ( .A(n_152), .Y(n_254) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_152), .Y(n_266) );
INVx2_ASAP7_75t_L g274 ( .A(n_152), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_152), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g383 ( .A(n_152), .B(n_268), .Y(n_383) );
AND2x2_ASAP7_75t_L g398 ( .A(n_152), .B(n_235), .Y(n_398) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_159), .B(n_161), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_158), .Y(n_153) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_159), .A2(n_164), .B(n_170), .Y(n_163) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_159), .A2(n_164), .B(n_170), .Y(n_318) );
AOI21x1_ASAP7_75t_L g466 ( .A1(n_159), .A2(n_467), .B(n_473), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_160), .Y(n_159) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_160), .A2(n_174), .B(n_178), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_160), .A2(n_459), .B(n_460), .Y(n_458) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_160), .A2(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g267 ( .A(n_163), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_163), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_169), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_171), .B(n_391), .Y(n_390) );
NOR2x1p5_ASAP7_75t_L g171 ( .A(n_172), .B(n_179), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g219 ( .A(n_173), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_173), .B(n_180), .Y(n_249) );
INVx1_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
INVx2_ASAP7_75t_L g282 ( .A(n_173), .Y(n_282) );
INVx2_ASAP7_75t_L g288 ( .A(n_173), .Y(n_288) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_173), .Y(n_358) );
OR2x2_ASAP7_75t_L g389 ( .A(n_173), .B(n_180), .Y(n_389) );
OR2x2_ASAP7_75t_L g405 ( .A(n_179), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x4_ASAP7_75t_SL g193 ( .A(n_180), .B(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_L g231 ( .A(n_180), .B(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g269 ( .A(n_180), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g281 ( .A(n_180), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g294 ( .A(n_180), .B(n_260), .Y(n_294) );
OR2x2_ASAP7_75t_L g302 ( .A(n_180), .B(n_194), .Y(n_302) );
INVx2_ASAP7_75t_L g329 ( .A(n_180), .Y(n_329) );
INVx1_ASAP7_75t_L g347 ( .A(n_180), .Y(n_347) );
NOR2xp33_ASAP7_75t_R g380 ( .A(n_180), .B(n_220), .Y(n_380) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_189), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_187), .Y(n_181) );
INVx2_ASAP7_75t_SL g237 ( .A(n_187), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_187), .A2(n_504), .B(n_505), .Y(n_503) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g214 ( .A(n_188), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_191), .B(n_229), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_191), .A2(n_272), .B1(n_275), .B2(n_278), .Y(n_271) );
OR2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_218), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g286 ( .A(n_193), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g321 ( .A(n_193), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g400 ( .A(n_193), .B(n_378), .Y(n_400) );
INVx3_ASAP7_75t_L g232 ( .A(n_194), .Y(n_232) );
AND2x4_ASAP7_75t_L g260 ( .A(n_194), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_194), .B(n_220), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_194), .B(n_282), .Y(n_327) );
AND2x2_ASAP7_75t_L g332 ( .A(n_194), .B(n_329), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_194), .B(n_219), .Y(n_369) );
INVx1_ASAP7_75t_L g439 ( .A(n_194), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_194), .B(n_357), .Y(n_450) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_210), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_198), .B1(n_203), .B2(n_208), .Y(n_195) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_202), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2x1p5_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g494 ( .A(n_213), .Y(n_494) );
INVx4_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI21x1_ASAP7_75t_L g221 ( .A1(n_214), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_214), .A2(n_475), .B(n_481), .Y(n_474) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_220), .B(n_232), .Y(n_250) );
INVx2_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
AND2x2_ASAP7_75t_L g287 ( .A(n_220), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g303 ( .A(n_220), .B(n_282), .Y(n_303) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_220), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_220), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g392 ( .A(n_220), .Y(n_392) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_227), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_230), .B(n_259), .Y(n_270) );
AOI221x1_ASAP7_75t_SL g364 ( .A1(n_231), .A2(n_365), .B1(n_368), .B2(n_370), .C(n_374), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_231), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_231), .B(n_287), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_231), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g353 ( .A(n_232), .B(n_281), .Y(n_353) );
AND2x2_ASAP7_75t_L g391 ( .A(n_232), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_242), .Y(n_234) );
AND2x2_ASAP7_75t_L g244 ( .A(n_235), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g339 ( .A(n_235), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_235), .B(n_255), .Y(n_344) );
AND2x4_ASAP7_75t_L g373 ( .A(n_235), .B(n_274), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_235), .B(n_305), .Y(n_409) );
OR2x2_ASAP7_75t_L g427 ( .A(n_235), .B(n_358), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_235), .B(n_318), .Y(n_437) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g268 ( .A(n_236), .Y(n_268) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_241), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g293 ( .A(n_242), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_242), .A2(n_301), .B1(n_304), .B2(n_306), .Y(n_300) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
INVx2_ASAP7_75t_L g256 ( .A(n_244), .Y(n_256) );
AND2x2_ASAP7_75t_L g395 ( .A(n_245), .B(n_255), .Y(n_395) );
AND2x2_ASAP7_75t_L g441 ( .A(n_245), .B(n_308), .Y(n_441) );
AND2x2_ASAP7_75t_L g446 ( .A(n_245), .B(n_297), .Y(n_446) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_247), .A2(n_317), .A3(n_397), .B1(n_416), .B2(n_418), .Y(n_415) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g283 ( .A(n_250), .Y(n_283) );
AOI211xp5_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_257), .B(n_262), .C(n_271), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .B(n_256), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_254), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_255), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g435 ( .A(n_255), .Y(n_435) );
AND2x2_ASAP7_75t_L g345 ( .A(n_257), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_SL g257 ( .A(n_258), .B(n_260), .Y(n_257) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_258), .Y(n_445) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_259), .Y(n_314) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_259), .Y(n_414) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
AND2x2_ASAP7_75t_L g377 ( .A(n_260), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_260), .B(n_388), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_269), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI21xp33_ASAP7_75t_L g343 ( .A1(n_264), .A2(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_SL g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_268), .B(n_274), .Y(n_273) );
BUFx2_ASAP7_75t_L g297 ( .A(n_268), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_273), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g404 ( .A(n_273), .Y(n_404) );
AND2x2_ASAP7_75t_L g434 ( .A(n_273), .B(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_274), .Y(n_411) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_276), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g351 ( .A(n_277), .Y(n_351) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g310 ( .A(n_281), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_282), .Y(n_378) );
AND2x2_ASAP7_75t_L g387 ( .A(n_283), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_307), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .B1(n_294), .B2(n_295), .C(n_300), .Y(n_285) );
INVx1_ASAP7_75t_L g406 ( .A(n_287), .Y(n_406) );
INVxp33_ASAP7_75t_SL g438 ( .A(n_287), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_289), .A2(n_385), .B(n_393), .Y(n_384) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_293), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g306 ( .A(n_294), .Y(n_306) );
AND2x2_ASAP7_75t_L g341 ( .A(n_294), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g360 ( .A(n_294), .B(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_294), .A2(n_422), .B1(n_423), .B2(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OR2x2_ASAP7_75t_L g316 ( .A(n_297), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_297), .B(n_305), .Y(n_355) );
AND2x4_ASAP7_75t_L g372 ( .A(n_299), .B(n_318), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_299), .B(n_373), .Y(n_419) );
AND2x2_ASAP7_75t_L g431 ( .A(n_299), .B(n_383), .Y(n_431) );
NAND2xp33_ASAP7_75t_L g416 ( .A(n_301), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_SL g359 ( .A(n_302), .Y(n_359) );
INVx1_ASAP7_75t_L g430 ( .A(n_303), .Y(n_430) );
INVx2_ASAP7_75t_SL g382 ( .A(n_305), .Y(n_382) );
AOI211xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_309), .B(n_312), .C(n_330), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI211xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B(n_319), .C(n_323), .Y(n_312) );
OR2x6_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
INVx1_ASAP7_75t_SL g367 ( .A(n_317), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_317), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_326), .A2(n_409), .B1(n_410), .B2(n_412), .Y(n_408) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
OAI211xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_340), .B(n_343), .C(n_348), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B1(n_354), .B2(n_356), .C(n_360), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_359), .A2(n_441), .B1(n_442), .B2(n_446), .C1(n_447), .C2(n_449), .Y(n_440) );
INVx2_ASAP7_75t_L g375 ( .A(n_361), .Y(n_375) );
NOR3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_401), .C(n_420), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_384), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_372), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_373), .B(n_435), .Y(n_448) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_379), .B2(n_381), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVxp33_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_382), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_390), .A2(n_394), .B1(n_396), .B2(n_399), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_405), .B(n_407), .C(n_415), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_428), .C(n_440), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_439), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx5_ASAP7_75t_L g757 ( .A(n_451), .Y(n_757) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_654), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_579), .C(n_615), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_553), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_482), .B(n_511), .C(n_536), .Y(n_454) );
AND2x2_ASAP7_75t_L g644 ( .A(n_455), .B(n_513), .Y(n_644) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_456), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g677 ( .A(n_456), .B(n_559), .Y(n_677) );
AND2x2_ASAP7_75t_L g693 ( .A(n_456), .B(n_528), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_456), .B(n_703), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_456), .B(n_727), .Y(n_726) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_SL g523 ( .A(n_457), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g548 ( .A(n_457), .Y(n_548) );
AND2x2_ASAP7_75t_L g595 ( .A(n_457), .B(n_538), .Y(n_595) );
AND2x2_ASAP7_75t_L g614 ( .A(n_457), .B(n_465), .Y(n_614) );
BUFx2_ASAP7_75t_L g619 ( .A(n_457), .Y(n_619) );
AND2x2_ASAP7_75t_L g663 ( .A(n_457), .B(n_474), .Y(n_663) );
AND2x4_ASAP7_75t_L g735 ( .A(n_457), .B(n_736), .Y(n_735) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_457), .B(n_527), .Y(n_747) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_464), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_465), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g666 ( .A(n_465), .Y(n_666) );
BUFx2_ASAP7_75t_L g715 ( .A(n_465), .Y(n_715) );
INVx1_ASAP7_75t_L g737 ( .A(n_465), .Y(n_737) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_474), .Y(n_465) );
INVx3_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_466), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
INVx2_ASAP7_75t_L g527 ( .A(n_474), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_474), .B(n_524), .Y(n_528) );
INVx2_ASAP7_75t_L g603 ( .A(n_474), .Y(n_603) );
OR2x2_ASAP7_75t_L g610 ( .A(n_474), .B(n_559), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
AND2x2_ASAP7_75t_L g565 ( .A(n_482), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g599 ( .A(n_482), .B(n_562), .Y(n_599) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
AND2x2_ASAP7_75t_L g635 ( .A(n_483), .B(n_534), .Y(n_635) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g592 ( .A(n_484), .B(n_493), .Y(n_592) );
AND2x2_ASAP7_75t_L g711 ( .A(n_484), .B(n_502), .Y(n_711) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g533 ( .A(n_485), .Y(n_533) );
INVx1_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
AND2x2_ASAP7_75t_L g607 ( .A(n_485), .B(n_493), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_485), .B(n_514), .Y(n_612) );
OR2x2_ASAP7_75t_L g675 ( .A(n_485), .B(n_502), .Y(n_675) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_485), .Y(n_684) );
AND2x2_ASAP7_75t_L g513 ( .A(n_492), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
NOR2x1_ASAP7_75t_SL g492 ( .A(n_493), .B(n_502), .Y(n_492) );
AO21x1_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_493) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
AND2x2_ASAP7_75t_L g530 ( .A(n_502), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g578 ( .A(n_502), .Y(n_578) );
NAND2x1_ASAP7_75t_L g588 ( .A(n_502), .B(n_514), .Y(n_588) );
OR2x2_ASAP7_75t_L g593 ( .A(n_502), .B(n_531), .Y(n_593) );
BUFx2_ASAP7_75t_L g649 ( .A(n_502), .Y(n_649) );
AND2x2_ASAP7_75t_L g685 ( .A(n_502), .B(n_564), .Y(n_685) );
AND2x2_ASAP7_75t_L g696 ( .A(n_502), .B(n_534), .Y(n_696) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_522), .B1(n_528), .B2(n_529), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_513), .A2(n_693), .B1(n_743), .B2(n_748), .Y(n_742) );
INVx4_ASAP7_75t_L g531 ( .A(n_514), .Y(n_531) );
INVx2_ASAP7_75t_L g562 ( .A(n_514), .Y(n_562) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_514), .Y(n_633) );
OR2x2_ASAP7_75t_L g648 ( .A(n_514), .B(n_534), .Y(n_648) );
OR2x2_ASAP7_75t_SL g674 ( .A(n_514), .B(n_675), .Y(n_674) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_SL g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx2_ASAP7_75t_SL g555 ( .A(n_523), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_523), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g623 ( .A(n_523), .B(n_571), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_523), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g545 ( .A(n_524), .Y(n_545) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
AND2x2_ASAP7_75t_L g626 ( .A(n_524), .B(n_603), .Y(n_626) );
INVx1_ASAP7_75t_L g736 ( .A(n_524), .Y(n_736) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_526), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_526), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g544 ( .A(n_527), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_528), .B(n_677), .Y(n_676) );
AOI321xp33_ASAP7_75t_L g698 ( .A1(n_529), .A2(n_600), .A3(n_668), .B1(n_699), .B2(n_700), .C(n_704), .Y(n_698) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_530), .Y(n_597) );
AND2x2_ASAP7_75t_L g622 ( .A(n_530), .B(n_551), .Y(n_622) );
AND2x2_ASAP7_75t_L g697 ( .A(n_530), .B(n_607), .Y(n_697) );
INVx1_ASAP7_75t_L g566 ( .A(n_531), .Y(n_566) );
BUFx2_ASAP7_75t_L g576 ( .A(n_531), .Y(n_576) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_531), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g621 ( .A(n_532), .Y(n_621) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
BUFx2_ASAP7_75t_L g628 ( .A(n_533), .Y(n_628) );
INVx2_ASAP7_75t_L g564 ( .A(n_534), .Y(n_564) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_534), .Y(n_587) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI21xp33_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_546), .B(n_549), .Y(n_536) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_537), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .Y(n_538) );
INVx3_ASAP7_75t_L g571 ( .A(n_539), .Y(n_571) );
AND2x2_ASAP7_75t_L g602 ( .A(n_539), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AND2x4_ASAP7_75t_L g559 ( .A(n_540), .B(n_541), .Y(n_559) );
INVx1_ASAP7_75t_L g642 ( .A(n_544), .Y(n_642) );
INVx1_ASAP7_75t_SL g727 ( .A(n_545), .Y(n_727) );
INVxp33_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_548), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g653 ( .A(n_548), .B(n_610), .Y(n_653) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g657 ( .A(n_550), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_550), .B(n_672), .Y(n_671) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_551), .B(n_588), .Y(n_643) );
NOR4xp25_ASAP7_75t_L g738 ( .A(n_551), .B(n_582), .C(n_739), .D(n_740), .Y(n_738) );
OR2x2_ASAP7_75t_L g706 ( .A(n_552), .B(n_707), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_560), .B1(n_565), .B2(n_567), .C(n_572), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g618 ( .A(n_557), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g638 ( .A(n_558), .Y(n_638) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g661 ( .A(n_559), .Y(n_661) );
AND2x2_ASAP7_75t_L g668 ( .A(n_559), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OR2x2_ASAP7_75t_L g605 ( .A(n_562), .B(n_606), .Y(n_605) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_564), .B(n_578), .Y(n_577) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g582 ( .A(n_569), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_569), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g574 ( .A(n_571), .Y(n_574) );
OAI321xp33_ASAP7_75t_L g686 ( .A1(n_571), .A2(n_679), .A3(n_687), .B1(n_692), .B2(n_694), .C(n_698), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
OR2x2_ASAP7_75t_L g641 ( .A(n_574), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g741 ( .A(n_577), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_578), .B(n_621), .Y(n_620) );
NAND2xp33_ASAP7_75t_SL g721 ( .A(n_578), .B(n_592), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_583), .B(n_594), .C(n_598), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g690 ( .A(n_587), .Y(n_690) );
INVx3_ASAP7_75t_L g629 ( .A(n_588), .Y(n_629) );
OR2x2_ASAP7_75t_L g732 ( .A(n_588), .B(n_606), .Y(n_732) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_590), .A2(n_674), .B1(n_676), .B2(n_678), .Y(n_673) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g672 ( .A(n_593), .Y(n_672) );
OR2x2_ASAP7_75t_L g749 ( .A(n_593), .B(n_606), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI21xp5_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_600), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_602), .B(n_619), .Y(n_718) );
AND2x2_ASAP7_75t_L g724 ( .A(n_602), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g669 ( .A(n_603), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B1(n_611), .B2(n_613), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_606), .A2(n_649), .B(n_651), .C(n_653), .Y(n_650) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_609), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_609), .B(n_701), .Y(n_723) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g695 ( .A(n_612), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_614), .A2(n_646), .B(n_649), .C(n_650), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_630), .C(n_645), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B1(n_622), .B2(n_623), .C1(n_624), .C2(n_627), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g679 ( .A(n_619), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_619), .B(n_652), .Y(n_705) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g639 ( .A(n_626), .Y(n_639) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g744 ( .A(n_628), .B(n_661), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_629), .A2(n_720), .B1(n_722), .B2(n_724), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_636), .B1(n_640), .B2(n_643), .C(n_644), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI21xp5_ASAP7_75t_SL g704 ( .A1(n_637), .A2(n_705), .B(n_706), .Y(n_704) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx2_ASAP7_75t_L g652 ( .A(n_638), .Y(n_652) );
AND2x2_ASAP7_75t_L g746 ( .A(n_638), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g730 ( .A(n_642), .Y(n_730) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g659 ( .A(n_648), .B(n_649), .Y(n_659) );
INVx1_ASAP7_75t_L g712 ( .A(n_648), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_686), .C(n_708), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_660), .B(n_662), .C(n_667), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_657), .A2(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_673), .C(n_680), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g691 ( .A(n_674), .Y(n_691) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_675), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_677), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g739 ( .A(n_677), .Y(n_739) );
AND2x2_ASAP7_75t_L g729 ( .A(n_679), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g699 ( .A(n_681), .Y(n_699) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g707 ( .A(n_683), .Y(n_707) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_695), .A2(n_729), .B1(n_731), .B2(n_733), .C(n_738), .Y(n_728) );
OAI21xp33_ASAP7_75t_SL g743 ( .A1(n_700), .A2(n_744), .B(n_745), .Y(n_743) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_719), .C(n_728), .D(n_742), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B1(n_716), .B2(n_717), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx11_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_SL g777 ( .A1(n_756), .A2(n_778), .B1(n_781), .B2(n_782), .Y(n_777) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_768), .A2(n_777), .B(n_783), .Y(n_776) );
NOR2xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_772), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
BUFx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx2_ASAP7_75t_R g785 ( .A(n_771), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_778), .Y(n_782) );
INVx1_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_790), .Y(n_799) );
AND2x4_ASAP7_75t_SL g790 ( .A(n_791), .B(n_792), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
endmodule