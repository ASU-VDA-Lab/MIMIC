module real_aes_17914_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_851, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_851;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
AND2x4_ASAP7_75t_L g112 ( .A(n_0), .B(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_1), .A2(n_4), .B1(n_269), .B2(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_2), .A2(n_43), .B1(n_150), .B2(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_3), .A2(n_23), .B1(n_210), .B2(n_242), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_5), .A2(n_16), .B1(n_182), .B2(n_184), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_6), .A2(n_62), .B1(n_146), .B2(n_212), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_7), .A2(n_17), .B1(n_150), .B2(n_155), .Y(n_508) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_9), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_10), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_11), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_12), .A2(n_18), .B1(n_145), .B2(n_149), .Y(n_144) );
BUFx2_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
OR2x2_ASAP7_75t_L g131 ( .A(n_13), .B(n_38), .Y(n_131) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_14), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_15), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_19), .A2(n_101), .B1(n_182), .B2(n_269), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_20), .A2(n_39), .B1(n_174), .B2(n_176), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_21), .B(n_183), .Y(n_231) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_22), .A2(n_59), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_24), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_25), .A2(n_55), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_25), .Y(n_134) );
INVx4_ASAP7_75t_R g533 ( .A(n_26), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_27), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_28), .B(n_153), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_29), .A2(n_47), .B1(n_195), .B2(n_198), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_30), .A2(n_54), .B1(n_182), .B2(n_198), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_31), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_32), .B(n_174), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_33), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_34), .B(n_242), .Y(n_576) );
INVx1_ASAP7_75t_L g615 ( .A(n_35), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_SL g551 ( .A1(n_36), .A2(n_150), .B(n_152), .C(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_37), .A2(n_56), .B1(n_150), .B2(n_198), .Y(n_560) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_38), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_40), .A2(n_88), .B1(n_150), .B2(n_209), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_41), .A2(n_81), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_41), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_42), .A2(n_46), .B1(n_150), .B2(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_44), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_45), .A2(n_60), .B1(n_182), .B2(n_196), .Y(n_271) );
INVx1_ASAP7_75t_L g573 ( .A(n_48), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_49), .B(n_150), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_50), .Y(n_592) );
INVx2_ASAP7_75t_L g121 ( .A(n_51), .Y(n_121) );
BUFx3_ASAP7_75t_L g116 ( .A(n_52), .Y(n_116) );
INVx1_ASAP7_75t_L g129 ( .A(n_52), .Y(n_129) );
INVx1_ASAP7_75t_L g848 ( .A(n_53), .Y(n_848) );
INVx1_ASAP7_75t_L g135 ( .A(n_55), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_57), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_58), .A2(n_89), .B1(n_150), .B2(n_198), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g830 ( .A1(n_61), .A2(n_831), .B1(n_832), .B2(n_835), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_61), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_63), .A2(n_76), .B1(n_195), .B2(n_196), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_64), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_65), .A2(n_78), .B1(n_150), .B2(n_155), .Y(n_219) );
AOI21xp33_ASAP7_75t_R g839 ( .A1(n_66), .A2(n_485), .B(n_840), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_67), .A2(n_99), .B1(n_149), .B2(n_182), .Y(n_218) );
INVx1_ASAP7_75t_L g162 ( .A(n_68), .Y(n_162) );
AND2x4_ASAP7_75t_L g164 ( .A(n_69), .B(n_165), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_70), .A2(n_91), .B1(n_195), .B2(n_198), .Y(n_611) );
AO22x1_ASAP7_75t_L g520 ( .A1(n_71), .A2(n_77), .B1(n_176), .B2(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g165 ( .A(n_72), .Y(n_165) );
AND2x2_ASAP7_75t_L g554 ( .A(n_73), .B(n_237), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_74), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_75), .B(n_212), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_79), .B(n_242), .Y(n_593) );
INVx2_ASAP7_75t_L g153 ( .A(n_80), .Y(n_153) );
INVx1_ASAP7_75t_L g834 ( .A(n_81), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_82), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_83), .B(n_237), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_84), .A2(n_98), .B1(n_198), .B2(n_212), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_85), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_86), .B(n_160), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_87), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_90), .B(n_237), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_92), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_93), .B(n_237), .Y(n_589) );
INVx1_ASAP7_75t_L g115 ( .A(n_94), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_94), .B(n_491), .Y(n_490) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_95), .B(n_183), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_96), .A2(n_157), .B(n_212), .C(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g535 ( .A(n_97), .B(n_536), .Y(n_535) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_100), .A2(n_123), .B(n_481), .Y(n_122) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_100), .Y(n_483) );
NAND2xp33_ASAP7_75t_L g597 ( .A(n_102), .B(n_175), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_117), .B(n_847), .Y(n_103) );
BUFx12f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx4f_ASAP7_75t_L g849 ( .A(n_105), .Y(n_849) );
AND2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_110), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_114), .C(n_116), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AND3x2_ASAP7_75t_L g127 ( .A(n_114), .B(n_128), .C(n_130), .Y(n_127) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g821 ( .A(n_115), .Y(n_821) );
INVx1_ASAP7_75t_L g828 ( .A(n_116), .Y(n_828) );
NOR2x1_ASAP7_75t_L g846 ( .A(n_116), .B(n_131), .Y(n_846) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_493), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx8_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g826 ( .A(n_121), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_121), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_132), .Y(n_124) );
BUFx2_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_127), .B(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g491 ( .A(n_129), .Y(n_491) );
AND2x6_ASAP7_75t_SL g489 ( .A(n_130), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_130), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_132), .Y(n_484) );
XNOR2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_136), .Y(n_132) );
NAND4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_356), .C(n_410), .D(n_449), .Y(n_136) );
NAND4xp75_ASAP7_75t_L g822 ( .A(n_137), .B(n_356), .C(n_410), .D(n_449), .Y(n_822) );
NOR2x1_ASAP7_75t_L g137 ( .A(n_138), .B(n_314), .Y(n_137) );
NAND3xp33_ASAP7_75t_SL g138 ( .A(n_139), .B(n_257), .C(n_296), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_204), .B1(n_247), .B2(n_252), .Y(n_139) );
INVx1_ASAP7_75t_L g420 ( .A(n_140), .Y(n_420) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_169), .Y(n_140) );
INVx1_ASAP7_75t_L g283 ( .A(n_141), .Y(n_283) );
BUFx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_SL g249 ( .A(n_142), .Y(n_249) );
AND2x2_ASAP7_75t_L g301 ( .A(n_142), .B(n_190), .Y(n_301) );
AND2x2_ASAP7_75t_L g340 ( .A(n_142), .B(n_171), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_142), .B(n_277), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_142), .B(n_476), .Y(n_475) );
AO31x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_158), .A3(n_163), .B(n_166), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_151), .B1(n_154), .B2(n_156), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_147), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g150 ( .A(n_148), .Y(n_150) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
INVx2_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_148), .Y(n_212) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_148), .Y(n_242) );
INVx1_ASAP7_75t_L g270 ( .A(n_148), .Y(n_270) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g155 ( .A(n_150), .Y(n_155) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_151), .A2(n_173), .B1(n_178), .B2(n_181), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_151), .A2(n_178), .B1(n_194), .B2(n_197), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_151), .A2(n_208), .B1(n_211), .B2(n_213), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_151), .A2(n_156), .B1(n_218), .B2(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_151), .A2(n_233), .B(n_234), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_151), .A2(n_178), .B1(n_241), .B2(n_243), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_151), .A2(n_178), .B1(n_268), .B2(n_271), .Y(n_267) );
OAI22x1_ASAP7_75t_L g507 ( .A1(n_151), .A2(n_213), .B1(n_508), .B2(n_509), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_151), .A2(n_516), .B1(n_559), .B2(n_560), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_151), .A2(n_213), .B1(n_611), .B2(n_612), .Y(n_610) );
INVx6_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp5_ASAP7_75t_L g229 ( .A1(n_152), .A2(n_155), .B(n_230), .C(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_152), .B(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_152), .A2(n_597), .B(n_598), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_152), .A2(n_515), .B(n_520), .C(n_523), .Y(n_636) );
BUFx8_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g157 ( .A(n_153), .Y(n_157) );
INVx2_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
INVx1_ASAP7_75t_L g550 ( .A(n_153), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_155), .A2(n_592), .B(n_593), .C(n_594), .Y(n_591) );
INVx1_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
AO31x2_ASAP7_75t_L g216 ( .A1(n_158), .A2(n_217), .A3(n_220), .B(n_222), .Y(n_216) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_158), .A2(n_543), .B(n_554), .Y(n_542) );
AO31x2_ASAP7_75t_L g609 ( .A1(n_158), .A2(n_199), .A3(n_610), .B(n_614), .Y(n_609) );
BUFx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_159), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g536 ( .A(n_159), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_159), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_159), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
INVx2_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
OAI21xp33_ASAP7_75t_L g523 ( .A1(n_160), .A2(n_518), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_163), .A2(n_172), .A3(n_186), .B(n_188), .Y(n_171) );
INVx2_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_163), .A2(n_240), .A3(n_244), .B(n_245), .Y(n_239) );
AO31x2_ASAP7_75t_L g506 ( .A1(n_163), .A2(n_203), .A3(n_507), .B(n_510), .Y(n_506) );
BUFx10_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
INVx1_ASAP7_75t_L g524 ( .A(n_164), .Y(n_524) );
BUFx10_ASAP7_75t_L g561 ( .A(n_164), .Y(n_561) );
NOR2xp33_ASAP7_75t_SL g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx2_ASAP7_75t_L g192 ( .A(n_167), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_167), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g324 ( .A(n_170), .B(n_299), .Y(n_324) );
OR2x2_ASAP7_75t_L g366 ( .A(n_170), .B(n_346), .Y(n_366) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_190), .Y(n_170) );
INVx2_ASAP7_75t_L g251 ( .A(n_171), .Y(n_251) );
INVx1_ASAP7_75t_L g277 ( .A(n_171), .Y(n_277) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_171), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_171), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g431 ( .A(n_171), .Y(n_431) );
AND2x2_ASAP7_75t_L g436 ( .A(n_171), .B(n_265), .Y(n_436) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g195 ( .A(n_175), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g532 ( .A1(n_175), .A2(n_185), .B1(n_533), .B2(n_534), .Y(n_532) );
OAI21xp33_ASAP7_75t_SL g569 ( .A1(n_176), .A2(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g516 ( .A(n_179), .Y(n_516) );
BUFx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g595 ( .A(n_180), .Y(n_595) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_183), .Y(n_521) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AO31x2_ASAP7_75t_L g206 ( .A1(n_186), .A2(n_199), .A3(n_207), .B(n_214), .Y(n_206) );
BUFx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_187), .B(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_187), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_SL g227 ( .A(n_187), .Y(n_227) );
INVx4_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_187), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g577 ( .A(n_187), .B(n_561), .Y(n_577) );
AND2x4_ASAP7_75t_L g250 ( .A(n_190), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g274 ( .A(n_190), .Y(n_274) );
INVx2_ASAP7_75t_L g323 ( .A(n_190), .Y(n_323) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_190), .Y(n_339) );
INVx1_ASAP7_75t_L g476 ( .A(n_190), .Y(n_476) );
AO31x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .A3(n_199), .B(n_201), .Y(n_190) );
AO31x2_ASAP7_75t_L g266 ( .A1(n_191), .A2(n_220), .A3(n_267), .B(n_272), .Y(n_266) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_191), .A2(n_527), .B(n_535), .Y(n_526) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_198), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g613 ( .A(n_198), .Y(n_613) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_SL g235 ( .A(n_200), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_203), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_224), .Y(n_204) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_205), .Y(n_304) );
AND2x2_ASAP7_75t_L g311 ( .A(n_205), .B(n_307), .Y(n_311) );
AND2x2_ASAP7_75t_L g368 ( .A(n_205), .B(n_355), .Y(n_368) );
AND2x4_ASAP7_75t_SL g477 ( .A(n_205), .B(n_279), .Y(n_477) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
BUFx2_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
OR2x2_ASAP7_75t_L g295 ( .A(n_206), .B(n_281), .Y(n_295) );
AND2x4_ASAP7_75t_L g308 ( .A(n_206), .B(n_256), .Y(n_308) );
INVx2_ASAP7_75t_L g336 ( .A(n_206), .Y(n_336) );
OR2x2_ASAP7_75t_L g362 ( .A(n_206), .B(n_239), .Y(n_362) );
INVx1_ASAP7_75t_L g415 ( .A(n_206), .Y(n_415) );
INVx2_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_210), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_213), .B(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g256 ( .A(n_216), .Y(n_256) );
BUFx2_ASAP7_75t_L g334 ( .A(n_216), .Y(n_334) );
AND2x2_ASAP7_75t_L g422 ( .A(n_216), .B(n_336), .Y(n_422) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_221), .A2(n_528), .B(n_531), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_224), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_238), .Y(n_224) );
AND2x4_ASAP7_75t_L g335 ( .A(n_225), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g409 ( .A(n_225), .B(n_256), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_225), .B(n_258), .Y(n_427) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx2_ASAP7_75t_L g360 ( .A(n_226), .Y(n_360) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_236), .Y(n_226) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_227), .A2(n_228), .B(n_236), .Y(n_262) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_232), .B(n_235), .Y(n_228) );
INVx2_ASAP7_75t_L g244 ( .A(n_237), .Y(n_244) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_237), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_238), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g280 ( .A(n_238), .Y(n_280) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_239), .Y(n_294) );
INVx1_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
AND2x2_ASAP7_75t_L g355 ( .A(n_239), .B(n_262), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_242), .B(n_546), .Y(n_545) );
AO31x2_ASAP7_75t_L g557 ( .A1(n_244), .A2(n_558), .A3(n_561), .B(n_562), .Y(n_557) );
AND2x2_ASAP7_75t_L g447 ( .A(n_247), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g480 ( .A(n_247), .B(n_345), .Y(n_480) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
INVx1_ASAP7_75t_L g443 ( .A(n_248), .Y(n_443) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g275 ( .A(n_249), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g310 ( .A(n_249), .B(n_265), .Y(n_310) );
INVx1_ASAP7_75t_L g320 ( .A(n_249), .Y(n_320) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
INVx2_ASAP7_75t_L g352 ( .A(n_249), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_249), .B(n_274), .Y(n_365) );
OR2x2_ASAP7_75t_L g374 ( .A(n_249), .B(n_328), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_249), .B(n_322), .Y(n_384) );
AND2x2_ASAP7_75t_L g453 ( .A(n_249), .B(n_431), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_250), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_250), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_250), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_250), .B(n_286), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_250), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g465 ( .A(n_250), .B(n_351), .Y(n_465) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_253), .A2(n_319), .B1(n_403), .B2(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_254), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g459 ( .A(n_255), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g479 ( .A(n_255), .B(n_355), .Y(n_479) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g291 ( .A(n_256), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_256), .B(n_280), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_256), .B(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_256), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B1(n_285), .B2(n_289), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_258), .B(n_260), .Y(n_347) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_258), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g462 ( .A(n_258), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .B1(n_278), .B2(n_282), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_261), .Y(n_418) );
INVx1_ASAP7_75t_L g460 ( .A(n_261), .Y(n_460) );
INVx1_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_275), .Y(n_263) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_264), .A2(n_349), .B(n_353), .C(n_354), .Y(n_348) );
INVx1_ASAP7_75t_L g386 ( .A(n_264), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_264), .B(n_340), .Y(n_424) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_274), .Y(n_264) );
INVx3_ASAP7_75t_L g346 ( .A(n_265), .Y(n_346) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g284 ( .A(n_266), .B(n_274), .Y(n_284) );
INVx2_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_270), .B(n_548), .Y(n_547) );
NAND2x1_ASAP7_75t_L g367 ( .A(n_275), .B(n_345), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_275), .B(n_338), .Y(n_377) );
INVx1_ASAP7_75t_L g406 ( .A(n_275), .Y(n_406) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_278), .A2(n_464), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_279), .A2(n_298), .B(n_302), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_279), .B(n_433), .Y(n_469) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx3_ASAP7_75t_L g328 ( .A(n_284), .Y(n_328) );
AND2x4_ASAP7_75t_L g446 ( .A(n_284), .B(n_313), .Y(n_446) );
AND2x2_ASAP7_75t_L g452 ( .A(n_284), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g383 ( .A(n_286), .Y(n_383) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g303 ( .A(n_287), .B(n_294), .Y(n_303) );
AND2x2_ASAP7_75t_L g429 ( .A(n_287), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
OR2x2_ASAP7_75t_L g350 ( .A(n_288), .B(n_323), .Y(n_350) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2x1p5_ASAP7_75t_L g361 ( .A(n_291), .B(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_291), .B(n_295), .Y(n_448) );
INVx1_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
NOR2x1_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp67_ASAP7_75t_SL g378 ( .A(n_295), .B(n_379), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_304), .B1(n_305), .B2(n_309), .C1(n_311), .C2(n_312), .Y(n_296) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_298), .A2(n_342), .B(n_347), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_299), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g466 ( .A(n_299), .Y(n_466) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_300), .Y(n_472) );
AND2x4_ASAP7_75t_L g312 ( .A(n_301), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_301), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g456 ( .A(n_301), .Y(n_456) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
AND2x2_ASAP7_75t_L g397 ( .A(n_306), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g390 ( .A(n_307), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g329 ( .A(n_308), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_331), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B1(n_325), .B2(n_329), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_324), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g343 ( .A(n_321), .Y(n_343) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g379 ( .A(n_330), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_330), .B(n_335), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_330), .B(n_433), .Y(n_432) );
AOI211x1_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_337), .B(n_341), .C(n_348), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_332), .A2(n_446), .B(n_447), .Y(n_445) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g398 ( .A(n_334), .B(n_335), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_335), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_335), .Y(n_391) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g455 ( .A(n_338), .B(n_436), .Y(n_455) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g353 ( .A(n_340), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_340), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g373 ( .A(n_346), .B(n_365), .Y(n_373) );
OR2x2_ASAP7_75t_L g474 ( .A(n_346), .B(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
INVx2_ASAP7_75t_L g444 ( .A(n_350), .Y(n_444) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND5xp2_ASAP7_75t_L g450 ( .A(n_353), .B(n_403), .C(n_451), .D(n_454), .E(n_456), .Y(n_450) );
AND2x2_ASAP7_75t_L g421 ( .A(n_355), .B(n_422), .Y(n_421) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_394), .Y(n_356) );
NAND2xp67_ASAP7_75t_SL g357 ( .A(n_358), .B(n_375), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_363), .B1(n_368), .B2(n_369), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND3xp33_ASAP7_75t_SL g363 ( .A(n_364), .B(n_366), .C(n_367), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
NAND3xp33_ASAP7_75t_SL g369 ( .A(n_370), .B(n_373), .C(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_SL g405 ( .A1(n_373), .A2(n_406), .B(n_407), .C(n_408), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_380), .B2(n_381), .C(n_385), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_382), .B(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_390), .B2(n_392), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_386), .A2(n_412), .B(n_438), .C(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g401 ( .A(n_387), .Y(n_401) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g426 ( .A(n_389), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_399), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g404 ( .A(n_398), .Y(n_404) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_402), .C(n_405), .Y(n_399) );
AND3x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_437), .C(n_445), .Y(n_410) );
AOI221x1_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_419), .B1(n_421), .B2(n_423), .C(n_425), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_432), .B2(n_435), .Y(n_425) );
INVx1_ASAP7_75t_L g439 ( .A(n_430), .Y(n_439) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AOI211x1_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_457), .B(n_463), .C(n_478), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B1(n_473), .B2(n_477), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_485), .Y(n_481) );
NOR2xp67_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
CKINVDCx8_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
OAI331xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_823), .A3(n_829), .B1(n_836), .B2(n_837), .B3(n_839), .C1(n_851), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g838 ( .A(n_495), .Y(n_838) );
AO22x2_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_818), .B1(n_819), .B2(n_822), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
NOR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_732), .Y(n_497) );
NAND4xp75_ASAP7_75t_L g498 ( .A(n_499), .B(n_637), .C(n_679), .D(n_703), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_537), .B(n_578), .C(n_616), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g723 ( .A(n_503), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g817 ( .A(n_503), .B(n_754), .Y(n_817) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_512), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g632 ( .A(n_505), .B(n_588), .Y(n_632) );
AND2x2_ASAP7_75t_L g673 ( .A(n_505), .B(n_634), .Y(n_673) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g584 ( .A(n_506), .B(n_526), .Y(n_584) );
OR2x2_ASAP7_75t_L g602 ( .A(n_506), .B(n_526), .Y(n_602) );
INVx2_ASAP7_75t_L g624 ( .A(n_506), .Y(n_624) );
AND2x2_ASAP7_75t_L g654 ( .A(n_506), .B(n_588), .Y(n_654) );
AND2x2_ASAP7_75t_L g683 ( .A(n_506), .B(n_525), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_506), .B(n_635), .Y(n_719) );
AND2x2_ASAP7_75t_L g696 ( .A(n_512), .B(n_625), .Y(n_696) );
INVx2_ASAP7_75t_L g791 ( .A(n_512), .Y(n_791) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .Y(n_512) );
INVx2_ASAP7_75t_L g583 ( .A(n_513), .Y(n_583) );
AND2x4_ASAP7_75t_L g622 ( .A(n_513), .B(n_526), .Y(n_622) );
AOI21x1_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_519), .B(n_522), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_516), .A2(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_524), .A2(n_544), .B(n_551), .Y(n_543) );
AND2x2_ASAP7_75t_L g781 ( .A(n_525), .B(n_583), .Y(n_781) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g645 ( .A(n_526), .Y(n_645) );
AND2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_588), .Y(n_702) );
AND2x2_ASAP7_75t_L g717 ( .A(n_526), .B(n_625), .Y(n_717) );
AND2x2_ASAP7_75t_L g739 ( .A(n_526), .B(n_583), .Y(n_739) );
OAI211xp5_ASAP7_75t_SL g786 ( .A1(n_537), .A2(n_787), .B(n_789), .C(n_796), .Y(n_786) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_564), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g773 ( .A(n_540), .B(n_709), .Y(n_773) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_555), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_541), .B(n_566), .Y(n_672) );
INVxp67_ASAP7_75t_L g686 ( .A(n_541), .Y(n_686) );
AND2x2_ASAP7_75t_L g706 ( .A(n_541), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_541), .B(n_619), .Y(n_713) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B(n_549), .Y(n_544) );
BUFx4f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_550), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g647 ( .A(n_555), .B(n_629), .Y(n_647) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g695 ( .A(n_556), .B(n_606), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_556), .B(n_609), .Y(n_701) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g605 ( .A(n_557), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g670 ( .A(n_557), .B(n_609), .Y(n_670) );
BUFx2_ASAP7_75t_L g677 ( .A(n_557), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_557), .B(n_609), .Y(n_757) );
INVx1_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g687 ( .A(n_565), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g816 ( .A(n_565), .B(n_605), .Y(n_816) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
AND2x2_ASAP7_75t_L g630 ( .A(n_566), .B(n_609), .Y(n_630) );
AND2x2_ASAP7_75t_L g676 ( .A(n_566), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g709 ( .A(n_566), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_566), .B(n_620), .Y(n_726) );
AND2x2_ASAP7_75t_L g765 ( .A(n_566), .B(n_766), .Y(n_765) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_574), .B(n_577), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_585), .B(n_603), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_580), .A2(n_744), .B1(n_745), .B2(n_747), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
AND2x2_ASAP7_75t_L g741 ( .A(n_581), .B(n_632), .Y(n_741) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g656 ( .A(n_582), .Y(n_656) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g805 ( .A(n_583), .B(n_625), .Y(n_805) );
AND2x2_ASAP7_75t_L g769 ( .A(n_584), .B(n_664), .Y(n_769) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_601), .Y(n_585) );
OR2x2_ASAP7_75t_L g666 ( .A(n_586), .B(n_643), .Y(n_666) );
OR2x2_ASAP7_75t_L g778 ( .A(n_586), .B(n_602), .Y(n_778) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g641 ( .A(n_587), .Y(n_641) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g625 ( .A(n_588), .Y(n_625) );
BUFx3_ASAP7_75t_L g707 ( .A(n_588), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_596), .B(n_599), .Y(n_590) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g775 ( .A(n_602), .B(n_634), .Y(n_775) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
AND2x2_ASAP7_75t_L g617 ( .A(n_605), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g658 ( .A(n_605), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g795 ( .A(n_605), .Y(n_795) );
INVx1_ASAP7_75t_L g814 ( .A(n_605), .Y(n_814) );
INVx2_ASAP7_75t_L g629 ( .A(n_606), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_606), .B(n_609), .Y(n_678) );
INVx1_ASAP7_75t_L g742 ( .A(n_607), .Y(n_742) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g803 ( .A(n_608), .Y(n_803) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g620 ( .A(n_609), .Y(n_620) );
INVx1_ASAP7_75t_L g710 ( .A(n_609), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_621), .B1(n_626), .B2(n_631), .Y(n_616) );
AND2x4_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g659 ( .A(n_619), .Y(n_659) );
AND2x2_ASAP7_75t_L g661 ( .A(n_619), .B(n_646), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_619), .B(n_629), .Y(n_721) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx3_ASAP7_75t_L g652 ( .A(n_622), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_622), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g746 ( .A(n_622), .B(n_730), .Y(n_746) );
INVx1_ASAP7_75t_L g650 ( .A(n_623), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_623), .A2(n_661), .B1(n_662), .B2(n_667), .C1(n_673), .C2(n_674), .Y(n_660) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_623), .A2(n_691), .B(n_692), .Y(n_690) );
AND2x2_ASAP7_75t_L g714 ( .A(n_623), .B(n_633), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_623), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
OR2x2_ASAP7_75t_L g643 ( .A(n_624), .B(n_635), .Y(n_643) );
INVx1_ASAP7_75t_L g731 ( .A(n_624), .Y(n_731) );
BUFx2_ASAP7_75t_L g665 ( .A(n_625), .Y(n_665) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_628), .B(n_669), .Y(n_698) );
OR2x2_ASAP7_75t_L g810 ( .A(n_628), .B(n_670), .Y(n_810) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g693 ( .A(n_630), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g808 ( .A(n_630), .Y(n_808) );
OAI31xp33_ASAP7_75t_L g789 ( .A1(n_631), .A2(n_790), .A3(n_792), .B(n_793), .Y(n_789) );
AND2x4_ASAP7_75t_SL g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_632), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_660), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_646), .B(n_648), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x6_ASAP7_75t_L g759 ( .A(n_641), .B(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g691 ( .A(n_644), .Y(n_691) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g782 ( .A(n_645), .B(n_719), .Y(n_782) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_647), .A2(n_736), .B1(n_738), .B2(n_740), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g796 ( .A1(n_647), .A2(n_708), .B(n_770), .C(n_797), .Y(n_796) );
AOI21xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B(n_657), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_652), .B(n_750), .C(n_751), .D(n_753), .Y(n_749) );
NAND2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_654), .B(n_656), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_654), .B(n_739), .Y(n_762) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g728 ( .A(n_659), .B(n_688), .Y(n_728) );
NAND2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_666), .A2(n_810), .B1(n_811), .B2(n_813), .Y(n_809) );
AOI221x1_ASAP7_75t_L g748 ( .A1(n_667), .A2(n_749), .B1(n_755), .B2(n_758), .C(n_761), .Y(n_748) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g688 ( .A(n_670), .Y(n_688) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g700 ( .A(n_672), .B(n_701), .Y(n_700) );
NAND2x1p5_ASAP7_75t_L g763 ( .A(n_673), .B(n_754), .Y(n_763) );
O2A1O1Ixp5_ASAP7_75t_L g776 ( .A1(n_674), .A2(n_758), .B(n_777), .C(n_779), .Y(n_776) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx2_ASAP7_75t_L g725 ( .A(n_677), .Y(n_725) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_689), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_681), .A2(n_699), .B1(n_769), .B2(n_770), .C(n_772), .Y(n_768) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g705 ( .A(n_683), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_683), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g804 ( .A(n_683), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
NAND2x1_ASAP7_75t_L g783 ( .A(n_686), .B(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g807 ( .A(n_686), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g747 ( .A(n_687), .Y(n_747) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B1(n_696), .B2(n_697), .C1(n_699), .C2(n_702), .Y(n_689) );
INVx1_ASAP7_75t_L g774 ( .A(n_693), .Y(n_774) );
INVx1_ASAP7_75t_L g737 ( .A(n_694), .Y(n_737) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g771 ( .A(n_695), .Y(n_771) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g712 ( .A(n_701), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g766 ( .A(n_701), .Y(n_766) );
AND2x2_ASAP7_75t_L g729 ( .A(n_702), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_722), .Y(n_703) );
AOI222xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B1(n_711), .B2(n_714), .C1(n_715), .C2(n_720), .Y(n_704) );
INVx3_ASAP7_75t_L g754 ( .A(n_707), .Y(n_754) );
BUFx2_ASAP7_75t_L g812 ( .A(n_707), .Y(n_812) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g784 ( .A(n_709), .Y(n_784) );
OR2x2_ASAP7_75t_L g794 ( .A(n_709), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_SL g752 ( .A(n_717), .Y(n_752) );
AND2x2_ASAP7_75t_L g797 ( .A(n_718), .B(n_754), .Y(n_797) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_719), .Y(n_750) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g756 ( .A(n_721), .B(n_757), .Y(n_756) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
OR2x2_ASAP7_75t_L g813 ( .A(n_726), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g744 ( .A(n_728), .Y(n_744) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g751 ( .A(n_731), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g801 ( .A(n_731), .Y(n_801) );
NAND4xp75_ASAP7_75t_L g732 ( .A(n_733), .B(n_767), .C(n_785), .D(n_798), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_748), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_742), .B(n_743), .Y(n_734) );
INVxp33_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_737), .B(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g760 ( .A(n_739), .Y(n_760) );
AND2x2_ASAP7_75t_L g800 ( .A(n_739), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g770 ( .A(n_742), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g788 ( .A(n_753), .Y(n_788) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp33_ASAP7_75t_SL g779 ( .A1(n_756), .A2(n_780), .B1(n_782), .B2(n_783), .Y(n_779) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI21xp33_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_763), .B(n_764), .Y(n_761) );
INVx1_ASAP7_75t_L g792 ( .A(n_763), .Y(n_792) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_776), .Y(n_767) );
AOI21xp5_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_774), .B(n_775), .Y(n_772) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_815), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_802), .B1(n_804), .B2(n_806), .C(n_809), .Y(n_799) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
BUFx12f_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
AND2x2_ASAP7_75t_L g845 ( .A(n_821), .B(n_846), .Y(n_845) );
CKINVDCx16_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
BUFx12f_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AND2x6_ASAP7_75t_SL g825 ( .A(n_826), .B(n_827), .Y(n_825) );
CKINVDCx6p67_ASAP7_75t_R g836 ( .A(n_829), .Y(n_836) );
BUFx3_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx10_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR2xp33_ASAP7_75t_R g847 ( .A(n_848), .B(n_849), .Y(n_847) );
endmodule