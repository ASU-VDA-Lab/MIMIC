module fake_netlist_6_3561_n_1712 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1712);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1712;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_44),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_15),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_20),
.Y(n_160)
);

BUFx8_ASAP7_75t_SL g161 ( 
.A(n_111),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_95),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_5),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_46),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_36),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_31),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_43),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_55),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_42),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_58),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_63),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_53),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_103),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_18),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_109),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_128),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_29),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_80),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_33),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_51),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_68),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_133),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_135),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_59),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_122),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_67),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_15),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_14),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_75),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_104),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_89),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_17),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_22),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_71),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_33),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_39),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_37),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_97),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_78),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_57),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_90),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_92),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_0),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_46),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_14),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_137),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_101),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_38),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_39),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_20),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_9),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_21),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_36),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_56),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_32),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_12),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_62),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_115),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_43),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_42),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_116),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_93),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_50),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_112),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_47),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_28),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_31),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_70),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_16),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_49),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_141),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_74),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_121),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_18),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_127),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_21),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_35),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_41),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_123),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_19),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_99),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_41),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_34),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_28),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_144),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_22),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_23),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_91),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_19),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_13),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_27),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_25),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_38),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_94),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_49),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_107),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_190),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_248),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_198),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_161),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_157),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_169),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_179),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_164),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_167),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_175),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_265),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_213),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_265),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_201),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_213),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_236),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_240),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_236),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_235),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_301),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_177),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_178),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_245),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_180),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_159),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_245),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_203),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_181),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_203),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_275),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_211),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_203),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_219),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_169),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_219),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_219),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_247),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_179),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_186),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_168),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_267),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_275),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_168),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_169),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_171),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_171),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_183),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_172),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_172),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_173),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_169),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_173),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_275),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_174),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_159),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_174),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_187),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_188),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_367),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_356),
.A2(n_279),
.B1(n_191),
.B2(n_223),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_303),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_284),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_156),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_317),
.A2(n_323),
.B1(n_321),
.B2(n_327),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_284),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_317),
.A2(n_249),
.B1(n_176),
.B2(n_299),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_284),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_325),
.A2(n_200),
.B(n_183),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_308),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_362),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_200),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_313),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_342),
.B(n_197),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_314),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_314),
.A2(n_195),
.B(n_184),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_232),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_334),
.B(n_193),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_345),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_345),
.B(n_154),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_322),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_315),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_347),
.A2(n_210),
.B(n_209),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_154),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_304),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_368),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_326),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_318),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_350),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_306),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_319),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_L g448 ( 
.A(n_394),
.B(n_320),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_386),
.A2(n_355),
.B1(n_324),
.B2(n_349),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_405),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_397),
.B(n_337),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_423),
.B(n_378),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_339),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_412),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_415),
.B(n_341),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_412),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_423),
.B(n_333),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_407),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_429),
.A2(n_305),
.B1(n_257),
.B2(n_184),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_346),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_417),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_357),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_429),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_396),
.B(n_209),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_394),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

NOR2x1p5_ASAP7_75t_L g482 ( 
.A(n_400),
.B(n_307),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

CKINVDCx6p67_ASAP7_75t_R g484 ( 
.A(n_439),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_415),
.B(n_377),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_SL g486 ( 
.A(n_386),
.B(n_257),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_418),
.B(n_194),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_359),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_409),
.B(n_350),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_409),
.B(n_351),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_409),
.B(n_351),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_427),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_384),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_446),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_446),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_439),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_435),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

INVx11_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

AND3x2_ASAP7_75t_L g507 ( 
.A(n_435),
.B(n_215),
.C(n_210),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_418),
.B(n_400),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_399),
.B(n_199),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_387),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_387),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_393),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_379),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_400),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_399),
.B(n_401),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_393),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_401),
.B(n_202),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_403),
.B(n_212),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_403),
.B(n_195),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_406),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_354),
.C(n_353),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_396),
.B(n_215),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_379),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_406),
.Y(n_531)
);

INVx11_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_380),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_407),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_403),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_406),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_380),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_408),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_419),
.B(n_216),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_392),
.B(n_358),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_383),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_408),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_408),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_438),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_438),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_438),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_413),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_258),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_383),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_420),
.B(n_358),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_413),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_392),
.B(n_360),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_413),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_388),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_421),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_413),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_388),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_426),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_422),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_404),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_422),
.B(n_360),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_389),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_392),
.B(n_361),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_426),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_425),
.B(n_361),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_425),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_389),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_424),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_430),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_424),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_430),
.B(n_166),
.C(n_165),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_432),
.B(n_224),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_424),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_432),
.B(n_226),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_437),
.B(n_227),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_392),
.B(n_228),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_391),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_426),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_391),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_436),
.B(n_165),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_395),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_532),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_450),
.Y(n_592)
);

O2A1O1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_463),
.A2(n_437),
.B(n_442),
.C(n_441),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_456),
.Y(n_594)
);

AOI221xp5_ASAP7_75t_SL g595 ( 
.A1(n_492),
.A2(n_440),
.B1(n_442),
.B2(n_441),
.C(n_302),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_488),
.B(n_424),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_518),
.A2(n_278),
.B1(n_258),
.B2(n_162),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_463),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_450),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_480),
.B(n_424),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_536),
.B(n_233),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_484),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_453),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_508),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_472),
.B(n_230),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_447),
.B(n_155),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_468),
.B(n_411),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_536),
.B(n_160),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_471),
.B(n_411),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_459),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_457),
.B(n_163),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_470),
.A2(n_260),
.B1(n_214),
.B2(n_283),
.Y(n_614)
);

O2A1O1Ixp5_ASAP7_75t_L g615 ( 
.A1(n_470),
.A2(n_402),
.B(n_414),
.C(n_416),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_454),
.B(n_411),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_456),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_477),
.B(n_169),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_548),
.B(n_234),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_464),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_473),
.B(n_395),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_472),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_540),
.B(n_170),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_532),
.Y(n_624)
);

O2A1O1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_476),
.A2(n_440),
.B(n_268),
.C(n_218),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_548),
.B(n_237),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_477),
.B(n_169),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_555),
.B(n_370),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_458),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_489),
.B(n_402),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_490),
.B(n_410),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_230),
.Y(n_632)
);

OA22x2_ASAP7_75t_L g633 ( 
.A1(n_519),
.A2(n_298),
.B1(n_223),
.B2(n_302),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_490),
.B(n_410),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_549),
.B(n_414),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_525),
.A2(n_264),
.B1(n_251),
.B2(n_252),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_461),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_549),
.A2(n_278),
.B1(n_254),
.B2(n_243),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_550),
.B(n_416),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_525),
.A2(n_269),
.B1(n_253),
.B2(n_255),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_462),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_458),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

AND2x6_ASAP7_75t_L g645 ( 
.A(n_561),
.B(n_166),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_464),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_485),
.B(n_189),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_496),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_469),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_560),
.B(n_270),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_451),
.B(n_204),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_476),
.B(n_443),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_483),
.B(n_443),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_483),
.B(n_443),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_505),
.A2(n_214),
.B1(n_244),
.B2(n_298),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_505),
.A2(n_217),
.B1(n_295),
.B2(n_218),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_511),
.B(n_443),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_511),
.A2(n_287),
.B(n_217),
.C(n_244),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_486),
.B(n_225),
.C(n_222),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_560),
.B(n_564),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_475),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_516),
.B(n_381),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_475),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_516),
.B(n_381),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_584),
.A2(n_390),
.B(n_382),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_504),
.B(n_282),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_555),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_574),
.B(n_206),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_529),
.B(n_381),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_529),
.B(n_381),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_533),
.B(n_381),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_533),
.B(n_539),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_561),
.B(n_553),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_539),
.B(n_381),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_560),
.B(n_288),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_477),
.B(n_169),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_448),
.A2(n_574),
.B1(n_522),
.B2(n_521),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_481),
.B(n_370),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_544),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_560),
.B(n_289),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_542),
.A2(n_291),
.B1(n_292),
.B2(n_300),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_557),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_571),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_564),
.B(n_182),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_481),
.A2(n_207),
.B1(n_276),
.B2(n_272),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_564),
.B(n_182),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_460),
.B(n_230),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_494),
.B(n_230),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_527),
.A2(n_436),
.B(n_294),
.C(n_185),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_495),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_479),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_577),
.B(n_208),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_545),
.B(n_382),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_577),
.A2(n_225),
.B1(n_222),
.B2(n_207),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_449),
.B(n_283),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_472),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_564),
.B(n_185),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_506),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_534),
.A2(n_196),
.B1(n_294),
.B2(n_276),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_469),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_487),
.A2(n_272),
.B1(n_196),
.B2(n_205),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_499),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_545),
.B(n_382),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_510),
.A2(n_192),
.B1(n_205),
.B2(n_243),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_382),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_554),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_467),
.B(n_192),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_580),
.B(n_220),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_502),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_499),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_527),
.B(n_254),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_559),
.B(n_382),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_559),
.B(n_382),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_563),
.B(n_382),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_563),
.B(n_382),
.Y(n_717)
);

INVxp33_ASAP7_75t_L g718 ( 
.A(n_449),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_568),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_570),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_221),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_583),
.B(n_229),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_497),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_570),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_561),
.A2(n_271),
.B1(n_231),
.B2(n_281),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_500),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_553),
.A2(n_567),
.B1(n_482),
.B2(n_588),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_573),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_575),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_452),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_500),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_575),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_585),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_385),
.Y(n_734)
);

AND2x6_ASAP7_75t_SL g735 ( 
.A(n_506),
.B(n_295),
.Y(n_735)
);

BUFx6f_ASAP7_75t_SL g736 ( 
.A(n_477),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_477),
.B(n_238),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_588),
.B(n_239),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_590),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_497),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_590),
.B(n_385),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_567),
.A2(n_436),
.B(n_434),
.C(n_433),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_579),
.B(n_241),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_589),
.A2(n_477),
.B1(n_528),
.B2(n_579),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_474),
.B(n_385),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_482),
.B(n_372),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_474),
.B(n_385),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_474),
.B(n_242),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_507),
.B(n_372),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_498),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_603),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_711),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_607),
.A2(n_474),
.B(n_491),
.C(n_501),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_606),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_742),
.A2(n_589),
.B(n_501),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_600),
.A2(n_466),
.B(n_535),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_604),
.B(n_491),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_604),
.A2(n_589),
.B1(n_290),
.B2(n_293),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_620),
.B(n_491),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_610),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_598),
.A2(n_589),
.B1(n_581),
.B2(n_501),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_649),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_612),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_607),
.B(n_478),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_647),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_719),
.B(n_728),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_719),
.B(n_491),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_728),
.B(n_501),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_727),
.A2(n_528),
.B1(n_477),
.B2(n_524),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_637),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_735),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_668),
.B(n_374),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_679),
.B(n_478),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_625),
.A2(n_589),
.B(n_587),
.C(n_586),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_646),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_646),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_675),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_642),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_613),
.A2(n_528),
.B1(n_569),
.B2(n_524),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_647),
.B(n_524),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_598),
.B(n_569),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_647),
.B(n_569),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_647),
.B(n_569),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_592),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_628),
.B(n_374),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_680),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_628),
.B(n_376),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_712),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_680),
.B(n_376),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_708),
.B(n_720),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_739),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_594),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_711),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_648),
.A2(n_528),
.B1(n_576),
.B2(n_581),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_617),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_596),
.A2(n_517),
.B(n_466),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_724),
.B(n_576),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_605),
.B(n_478),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_729),
.B(n_528),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_732),
.Y(n_801)
);

BUFx4f_ASAP7_75t_L g802 ( 
.A(n_700),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_731),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_733),
.B(n_528),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_674),
.B(n_465),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_630),
.B(n_465),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_629),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_663),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_631),
.B(n_465),
.Y(n_809)
);

NOR2x2_ASAP7_75t_L g810 ( 
.A(n_697),
.B(n_433),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_652),
.A2(n_581),
.B1(n_466),
.B2(n_465),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_643),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_634),
.B(n_466),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_675),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_662),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_665),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_614),
.A2(n_578),
.B1(n_517),
.B2(n_535),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_599),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_650),
.B(n_326),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_650),
.B(n_328),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_702),
.B(n_478),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_726),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_614),
.A2(n_552),
.B1(n_586),
.B2(n_572),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_659),
.A2(n_587),
.B(n_572),
.C(n_565),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_671),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_608),
.A2(n_578),
.B(n_535),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_692),
.B(n_543),
.Y(n_827)
);

AND2x4_ASAP7_75t_SL g828 ( 
.A(n_726),
.B(n_543),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_656),
.A2(n_552),
.B1(n_565),
.B2(n_562),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_702),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_692),
.B(n_543),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_609),
.B(n_669),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_672),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_681),
.B(n_578),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_702),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_675),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_591),
.B(n_328),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_632),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_704),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_633),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_664),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_673),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_676),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_669),
.B(n_330),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_330),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_622),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_656),
.A2(n_552),
.B1(n_558),
.B2(n_556),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_702),
.Y(n_848)
);

OAI21xp33_ASAP7_75t_SL g849 ( 
.A1(n_657),
.A2(n_744),
.B(n_640),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_623),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_609),
.B(n_246),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_695),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_694),
.B(n_250),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_635),
.B(n_661),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_744),
.B(n_478),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_730),
.B(n_256),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_705),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_698),
.B(n_331),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_707),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_746),
.B(n_493),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_657),
.A2(n_493),
.B1(n_558),
.B2(n_556),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_684),
.B(n_498),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_714),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_670),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_675),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_602),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_715),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_645),
.Y(n_868)
);

INVxp33_ASAP7_75t_L g869 ( 
.A(n_689),
.Y(n_869)
);

AND3x1_ASAP7_75t_L g870 ( 
.A(n_660),
.B(n_344),
.C(n_338),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_716),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_730),
.B(n_259),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_717),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_749),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_734),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_638),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_693),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_633),
.A2(n_552),
.B1(n_562),
.B2(n_551),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_750),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_685),
.B(n_503),
.Y(n_880)
);

BUFx8_ASAP7_75t_L g881 ( 
.A(n_624),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_SL g882 ( 
.A(n_706),
.B(n_263),
.C(n_286),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_645),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_653),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_623),
.B(n_710),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_690),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_593),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_723),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_SL g889 ( 
.A(n_639),
.B(n_261),
.C(n_262),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_697),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_601),
.B(n_266),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_667),
.Y(n_892)
);

AND3x1_ASAP7_75t_L g893 ( 
.A(n_660),
.B(n_331),
.C(n_344),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_738),
.B(n_509),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_738),
.B(n_509),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_737),
.B(n_493),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_748),
.B(n_512),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_748),
.B(n_611),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_743),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_740),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_645),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_741),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_721),
.B(n_493),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_645),
.A2(n_552),
.B1(n_547),
.B2(n_546),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_722),
.B(n_493),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_621),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_615),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_645),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_619),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_697),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_686),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_616),
.A2(n_390),
.B(n_398),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_654),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_688),
.A2(n_552),
.B1(n_546),
.B2(n_541),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_699),
.A2(n_552),
.B1(n_541),
.B2(n_538),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_626),
.B(n_725),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_655),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_615),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_658),
.B(n_513),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_703),
.B(n_513),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_713),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_745),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_597),
.B(n_514),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_747),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_595),
.B(n_514),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_789),
.B(n_709),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_752),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_832),
.B(n_636),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_832),
.A2(n_736),
.B1(n_718),
.B2(n_651),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_677),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_853),
.A2(n_641),
.B(n_682),
.C(n_691),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_898),
.A2(n_896),
.B(n_805),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_850),
.B(n_683),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_850),
.B(n_696),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_754),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_896),
.A2(n_678),
.B(n_627),
.Y(n_936)
);

NAND2x1_ASAP7_75t_L g937 ( 
.A(n_865),
.B(n_515),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_845),
.B(n_844),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_897),
.A2(n_618),
.B(n_666),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_853),
.A2(n_687),
.B(n_701),
.C(n_526),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_806),
.A2(n_390),
.B(n_398),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_766),
.B(n_273),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_794),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_809),
.A2(n_390),
.B(n_398),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_906),
.B(n_515),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_885),
.A2(n_433),
.B(n_538),
.C(n_537),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_794),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_848),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_838),
.B(n_332),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_751),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_838),
.B(n_332),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_891),
.A2(n_736),
.B1(n_537),
.B2(n_531),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_884),
.B(n_531),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_849),
.A2(n_887),
.B(n_854),
.C(n_758),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_882),
.A2(n_916),
.B1(n_758),
.B2(n_840),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_884),
.B(n_530),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_822),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_851),
.B(n_338),
.Y(n_958)
);

NAND2x1_ASAP7_75t_L g959 ( 
.A(n_865),
.B(n_530),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_813),
.A2(n_755),
.B(n_764),
.Y(n_960)
);

NOR2x1_ASAP7_75t_SL g961 ( 
.A(n_777),
.B(n_526),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_912),
.A2(n_523),
.B(n_520),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_776),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_778),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_891),
.A2(n_856),
.B(n_872),
.C(n_911),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_773),
.A2(n_385),
.B(n_390),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_869),
.B(n_285),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_784),
.B(n_274),
.Y(n_968)
);

AND2x2_ASAP7_75t_SL g969 ( 
.A(n_890),
.B(n_434),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_818),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_886),
.B(n_277),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_787),
.B(n_523),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_775),
.B(n_434),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_L g974 ( 
.A1(n_856),
.A2(n_872),
.B(n_790),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_762),
.B(n_520),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_797),
.A2(n_398),
.B(n_390),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_776),
.B(n_0),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_R g978 ( 
.A(n_892),
.B(n_66),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_803),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_911),
.B(n_1),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_777),
.B(n_398),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_760),
.Y(n_982)
);

INVx6_ASAP7_75t_L g983 ( 
.A(n_881),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_SL g984 ( 
.A(n_889),
.B(n_434),
.C(n_3),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_839),
.B(n_1),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_777),
.B(n_814),
.Y(n_986)
);

BUFx8_ASAP7_75t_L g987 ( 
.A(n_876),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_903),
.A2(n_905),
.B(n_761),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_786),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_848),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_848),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_SL g992 ( 
.A(n_846),
.B(n_398),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_882),
.A2(n_398),
.B1(n_390),
.B2(n_385),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_900),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_900),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_925),
.A2(n_398),
.B(n_390),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_777),
.A2(n_385),
.B1(n_64),
.B2(n_72),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_763),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_790),
.B(n_4),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_817),
.A2(n_385),
.B(n_61),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_756),
.A2(n_73),
.B(n_146),
.Y(n_1001)
);

OA21x2_ASAP7_75t_L g1002 ( 
.A1(n_753),
.A2(n_60),
.B(n_145),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_814),
.B(n_153),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_899),
.B(n_8),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_864),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_770),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_840),
.A2(n_8),
.B(n_10),
.C(n_12),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_866),
.B(n_143),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_801),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_917),
.B(n_10),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_879),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_877),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_923),
.A2(n_17),
.B(n_24),
.C(n_25),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_810),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_848),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_827),
.B(n_24),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_791),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_SL g1018 ( 
.A1(n_890),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_814),
.B(n_87),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_855),
.A2(n_86),
.B(n_129),
.C(n_126),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_827),
.B(n_30),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_831),
.B(n_32),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_781),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_909),
.A2(n_921),
.B1(n_788),
.B2(n_831),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_888),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_819),
.A2(n_98),
.B1(n_110),
.B2(n_108),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_792),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_759),
.B(n_37),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_855),
.A2(n_83),
.B(n_106),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_SL g1030 ( 
.A(n_889),
.B(n_40),
.C(n_45),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_881),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_894),
.A2(n_105),
.B(n_102),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_895),
.A2(n_100),
.B(n_142),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_759),
.B(n_40),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_837),
.B(n_45),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_SL g1036 ( 
.A(n_799),
.B(n_47),
.C(n_48),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_808),
.B(n_50),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_858),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_816),
.B(n_825),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_814),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_793),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_834),
.A2(n_826),
.B(n_774),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_836),
.B(n_802),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_796),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_819),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_865),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_772),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_836),
.A2(n_865),
.B1(n_913),
.B2(n_779),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_807),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_812),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_772),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_802),
.B(n_765),
.Y(n_1052)
);

BUFx4f_ASAP7_75t_L g1053 ( 
.A(n_837),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_836),
.B(n_874),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_858),
.B(n_820),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_774),
.A2(n_804),
.B(n_800),
.C(n_769),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_757),
.B(n_767),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_910),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_833),
.B(n_859),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_842),
.B(n_871),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_820),
.B(n_828),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_836),
.B(n_913),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_771),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_913),
.B(n_765),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_768),
.B(n_913),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_795),
.A2(n_811),
.B1(n_901),
.B2(n_880),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_860),
.A2(n_907),
.B1(n_918),
.B2(n_873),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_870),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_976),
.A2(n_824),
.B(n_798),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_991),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_976),
.A2(n_824),
.B(n_919),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_938),
.B(n_867),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_974),
.B(n_841),
.Y(n_1073)
);

AO32x2_ASAP7_75t_L g1074 ( 
.A1(n_929),
.A2(n_861),
.A3(n_893),
.B1(n_878),
.B2(n_857),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_962),
.A2(n_966),
.B(n_996),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_928),
.A2(n_815),
.B1(n_830),
.B2(n_835),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_955),
.A2(n_823),
.B1(n_829),
.B2(n_847),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1055),
.B(n_830),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_983),
.B(n_868),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1017),
.B(n_875),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_966),
.A2(n_924),
.B(n_922),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_950),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_965),
.A2(n_901),
.B(n_863),
.C(n_852),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1039),
.B(n_843),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_960),
.A2(n_902),
.B(n_862),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_1000),
.A2(n_821),
.B(n_780),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_927),
.B(n_868),
.Y(n_1087)
);

AO31x2_ASAP7_75t_L g1088 ( 
.A1(n_1067),
.A2(n_920),
.A3(n_878),
.B(n_904),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_SL g1089 ( 
.A1(n_1048),
.A2(n_908),
.B(n_883),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_941),
.A2(n_780),
.B(n_783),
.Y(n_1090)
);

NAND2x1_ASAP7_75t_L g1091 ( 
.A(n_1040),
.B(n_868),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_949),
.B(n_1014),
.Y(n_1092)
);

AOI31xp67_ASAP7_75t_L g1093 ( 
.A1(n_952),
.A2(n_783),
.A3(n_915),
.B(n_914),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_983),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_987),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1068),
.B(n_782),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_941),
.A2(n_782),
.B(n_904),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_991),
.Y(n_1098)
);

BUFx2_ASAP7_75t_SL g1099 ( 
.A(n_979),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_982),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_998),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_987),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_931),
.A2(n_954),
.B(n_1000),
.C(n_933),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_958),
.B(n_868),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_970),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_960),
.A2(n_954),
.B(n_1056),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1024),
.B(n_883),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1006),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1066),
.A2(n_829),
.B(n_847),
.Y(n_1109)
);

AO32x2_ASAP7_75t_L g1110 ( 
.A1(n_997),
.A2(n_883),
.A3(n_908),
.B1(n_948),
.B2(n_1013),
.Y(n_1110)
);

INVx3_ASAP7_75t_SL g1111 ( 
.A(n_983),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_SL g1112 ( 
.A1(n_1029),
.A2(n_1033),
.B(n_1032),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_957),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1058),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1042),
.A2(n_988),
.A3(n_1057),
.B(n_1065),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_988),
.A2(n_936),
.A3(n_940),
.B(n_944),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_1016),
.A2(n_1022),
.B(n_1021),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_978),
.Y(n_1118)
);

NAND4xp25_ASAP7_75t_L g1119 ( 
.A(n_1018),
.B(n_985),
.C(n_947),
.D(n_1035),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_1028),
.A2(n_1034),
.B(n_1013),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1029),
.A2(n_1001),
.A3(n_961),
.B(n_1033),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_991),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_968),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_992),
.B(n_1053),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_1001),
.A2(n_1032),
.A3(n_1037),
.B(n_956),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1015),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_946),
.A2(n_959),
.B(n_937),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1009),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_1015),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1031),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1053),
.B(n_969),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_946),
.A2(n_1062),
.B(n_953),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1064),
.A2(n_986),
.B(n_1020),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1010),
.A2(n_1059),
.A3(n_1060),
.B(n_980),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_SL g1136 ( 
.A1(n_1007),
.A2(n_1026),
.B(n_1002),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_951),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_1004),
.A2(n_977),
.B1(n_934),
.B2(n_930),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_L g1139 ( 
.A(n_1008),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_943),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1020),
.A2(n_945),
.B(n_1002),
.Y(n_1141)
);

AO32x2_ASAP7_75t_L g1142 ( 
.A1(n_948),
.A2(n_1007),
.A3(n_1038),
.B1(n_1036),
.B2(n_1040),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1023),
.A2(n_1051),
.B(n_1047),
.C(n_930),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_SL g1144 ( 
.A1(n_942),
.A2(n_972),
.B(n_971),
.C(n_1019),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1023),
.A2(n_981),
.B(n_1054),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_973),
.B(n_1011),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1015),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_SL g1148 ( 
.A1(n_1027),
.A2(n_935),
.B(n_989),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1045),
.B(n_967),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_984),
.A2(n_1003),
.B(n_1030),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_993),
.A2(n_984),
.B(n_1030),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_964),
.B(n_1012),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1005),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1025),
.B(n_1049),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1043),
.A2(n_1061),
.B(n_1046),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1046),
.A2(n_975),
.B(n_990),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_990),
.A2(n_1041),
.B(n_1044),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1050),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_SL g1159 ( 
.A1(n_994),
.A2(n_995),
.B(n_999),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1052),
.A2(n_926),
.B(n_963),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_926),
.A2(n_963),
.B(n_1008),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_943),
.B(n_926),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1063),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1018),
.B(n_938),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_960),
.A2(n_932),
.B(n_954),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_938),
.B(n_604),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_965),
.A2(n_832),
.B(n_853),
.C(n_607),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1040),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_932),
.A2(n_898),
.B(n_939),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_950),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_996),
.A2(n_896),
.B(n_1067),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_976),
.A2(n_962),
.B(n_966),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_938),
.A2(n_832),
.B1(n_853),
.B2(n_607),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_932),
.A2(n_898),
.B(n_939),
.Y(n_1174)
);

OA22x2_ASAP7_75t_L g1175 ( 
.A1(n_1024),
.A2(n_519),
.B1(n_697),
.B2(n_449),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1055),
.B(n_838),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_938),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_938),
.A2(n_832),
.B1(n_656),
.B2(n_657),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_938),
.A2(n_832),
.B1(n_853),
.B2(n_607),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_976),
.A2(n_962),
.B(n_966),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_991),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_947),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_991),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_991),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_SL g1185 ( 
.A1(n_1029),
.A2(n_954),
.B(n_1032),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1067),
.A2(n_1000),
.A3(n_1042),
.B(n_960),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1040),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_938),
.B(n_832),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_938),
.B(n_604),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_991),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_SL g1191 ( 
.A1(n_1029),
.A2(n_954),
.B(n_1032),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_938),
.B(n_832),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_987),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_938),
.B(n_832),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_938),
.B(n_832),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1016),
.A2(n_1022),
.B(n_1021),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_938),
.A2(n_832),
.B1(n_656),
.B2(n_657),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_950),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_976),
.A2(n_962),
.B(n_966),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_938),
.B(n_832),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1055),
.B(n_838),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_938),
.B(n_604),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_970),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_938),
.B(n_832),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_932),
.A2(n_898),
.B(n_939),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_932),
.A2(n_898),
.B(n_939),
.Y(n_1206)
);

AO21x1_ASAP7_75t_L g1207 ( 
.A1(n_1151),
.A2(n_1179),
.B(n_1173),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1169),
.A2(n_1205),
.B(n_1174),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_SL g1209 ( 
.A(n_1099),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1082),
.Y(n_1210)
);

INVx6_ASAP7_75t_L g1211 ( 
.A(n_1094),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1173),
.A2(n_1179),
.B1(n_1188),
.B2(n_1195),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1114),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1194),
.B(n_1204),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1078),
.B(n_1161),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1192),
.A2(n_1200),
.B(n_1197),
.C(n_1178),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1168),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1140),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1177),
.A2(n_1119),
.B1(n_1149),
.B2(n_1132),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1166),
.B(n_1189),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1075),
.A2(n_1199),
.B(n_1172),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1139),
.A2(n_1202),
.B1(n_1166),
.B2(n_1189),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1202),
.B(n_1072),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1077),
.A2(n_1197),
.B(n_1178),
.C(n_1106),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1176),
.B(n_1201),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1102),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1072),
.B(n_1084),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1120),
.A2(n_1144),
.B(n_1143),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1090),
.A2(n_1069),
.B(n_1081),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1083),
.A2(n_1077),
.A3(n_1073),
.B(n_1145),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1071),
.A2(n_1128),
.B(n_1097),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1185),
.A2(n_1191),
.B(n_1112),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1141),
.A2(n_1157),
.B(n_1085),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1120),
.A2(n_1165),
.B(n_1136),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1085),
.A2(n_1133),
.B(n_1134),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1196),
.A2(n_1109),
.B(n_1160),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1119),
.B(n_1164),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1084),
.B(n_1080),
.Y(n_1238)
);

AO21x2_ASAP7_75t_L g1239 ( 
.A1(n_1151),
.A2(n_1117),
.B(n_1086),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1156),
.A2(n_1089),
.B(n_1155),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1091),
.A2(n_1159),
.B(n_1076),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1139),
.A2(n_1164),
.B1(n_1137),
.B2(n_1104),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1146),
.A2(n_1107),
.B(n_1175),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1137),
.B(n_1092),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1113),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1100),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1152),
.A2(n_1154),
.B(n_1129),
.C(n_1198),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1162),
.A2(n_1182),
.B1(n_1170),
.B2(n_1101),
.C(n_1108),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1148),
.A2(n_1187),
.B(n_1087),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1152),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1182),
.B(n_1078),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1094),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1079),
.B(n_1096),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1150),
.A2(n_1122),
.B1(n_1158),
.B2(n_1153),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1105),
.A2(n_1111),
.B1(n_1079),
.B2(n_1154),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1187),
.A2(n_1093),
.B(n_1121),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1135),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1121),
.A2(n_1116),
.B(n_1186),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1135),
.B(n_1079),
.Y(n_1259)
);

AOI222xp33_ASAP7_75t_L g1260 ( 
.A1(n_1193),
.A2(n_1095),
.B1(n_1131),
.B2(n_1203),
.C1(n_1163),
.C2(n_1124),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1125),
.B(n_1130),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1118),
.A2(n_1150),
.B1(n_1181),
.B2(n_1127),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1121),
.A2(n_1116),
.B(n_1186),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1115),
.A2(n_1126),
.B(n_1088),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1126),
.A2(n_1115),
.B(n_1110),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1135),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1088),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1181),
.A2(n_1098),
.B(n_1130),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1126),
.A2(n_1074),
.B(n_1110),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1190),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1074),
.A2(n_1142),
.B(n_1098),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1070),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1074),
.A2(n_1142),
.B(n_1130),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1142),
.A2(n_1123),
.A3(n_1127),
.B1(n_1147),
.B2(n_1183),
.Y(n_1274)
);

AND2x6_ASAP7_75t_L g1275 ( 
.A(n_1123),
.B(n_1127),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1147),
.A2(n_1190),
.B1(n_1183),
.B2(n_1184),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1184),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1184),
.A2(n_832),
.B1(n_1179),
.B2(n_1173),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1167),
.A2(n_832),
.B(n_965),
.C(n_607),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1173),
.A2(n_832),
.B1(n_1179),
.B2(n_853),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1167),
.A2(n_832),
.B(n_1173),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1082),
.Y(n_1282)
);

AOI22x1_ASAP7_75t_L g1283 ( 
.A1(n_1138),
.A2(n_1191),
.B1(n_1185),
.B2(n_1112),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1075),
.A2(n_1180),
.B(n_1172),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1167),
.A2(n_1103),
.B(n_1169),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1176),
.B(n_1201),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1113),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_SL g1288 ( 
.A(n_1124),
.B(n_592),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1168),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1075),
.A2(n_1180),
.B(n_1172),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1075),
.A2(n_1180),
.B(n_1172),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1171),
.A2(n_996),
.B(n_1000),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1167),
.A2(n_1103),
.B(n_1169),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1167),
.A2(n_832),
.B(n_1173),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1089),
.B(n_1161),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1075),
.A2(n_1180),
.B(n_1172),
.Y(n_1296)
);

AOI221xp5_ASAP7_75t_L g1297 ( 
.A1(n_1167),
.A2(n_832),
.B1(n_853),
.B2(n_607),
.C(n_486),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_1194),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1078),
.B(n_1161),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1137),
.B(n_1166),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1075),
.A2(n_1180),
.B(n_1172),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1082),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1113),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1082),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1137),
.B(n_1166),
.Y(n_1305)
);

AND2x4_ASAP7_75t_SL g1306 ( 
.A(n_1094),
.B(n_1203),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1188),
.B(n_1194),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1168),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1078),
.B(n_1161),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1098),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1075),
.A2(n_1180),
.B(n_1172),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1168),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1124),
.B(n_592),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1168),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_L g1315 ( 
.A(n_1167),
.B(n_1077),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1167),
.A2(n_832),
.B(n_1173),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1113),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1188),
.B(n_1194),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1188),
.B(n_1194),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1124),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1168),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1103),
.A2(n_1167),
.A3(n_1206),
.B(n_1205),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1114),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1082),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1098),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1082),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1167),
.A2(n_832),
.B(n_1173),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1173),
.A2(n_832),
.B1(n_1179),
.B2(n_853),
.Y(n_1328)
);

AOI221x1_ASAP7_75t_SL g1329 ( 
.A1(n_1237),
.A2(n_1222),
.B1(n_1214),
.B2(n_1220),
.C(n_1319),
.Y(n_1329)
);

AOI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1297),
.A2(n_1328),
.B1(n_1280),
.B2(n_1279),
.C(n_1327),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1225),
.B(n_1286),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1214),
.B(n_1223),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1278),
.A2(n_1261),
.B(n_1238),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1227),
.A2(n_1224),
.B(n_1261),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1287),
.Y(n_1335)
);

AOI211xp5_ASAP7_75t_L g1336 ( 
.A1(n_1237),
.A2(n_1207),
.B(n_1216),
.C(n_1315),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1228),
.A2(n_1265),
.B(n_1263),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1280),
.A2(n_1328),
.B(n_1293),
.C(n_1285),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1253),
.B(n_1219),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1209),
.A2(n_1307),
.B1(n_1298),
.B2(n_1318),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1245),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1315),
.A2(n_1224),
.B(n_1208),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1215),
.B(n_1299),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1253),
.B(n_1251),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1253),
.B(n_1300),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1216),
.A2(n_1212),
.B(n_1243),
.C(n_1271),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1305),
.B(n_1244),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1242),
.B(n_1210),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1209),
.A2(n_1248),
.B1(n_1262),
.B2(n_1254),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1239),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1211),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1265),
.A2(n_1258),
.B(n_1235),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1254),
.A2(n_1257),
.B(n_1266),
.C(n_1312),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1317),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1218),
.A2(n_1303),
.B1(n_1255),
.B2(n_1211),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1306),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1250),
.B(n_1218),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1211),
.A2(n_1259),
.B1(n_1306),
.B2(n_1272),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1282),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1272),
.A2(n_1246),
.B1(n_1213),
.B2(n_1323),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1269),
.A2(n_1229),
.B(n_1256),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1252),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1247),
.A2(n_1326),
.B(n_1302),
.C(n_1304),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1213),
.A2(n_1323),
.B1(n_1324),
.B2(n_1276),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1247),
.A2(n_1234),
.B(n_1260),
.C(n_1232),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1283),
.A2(n_1295),
.B1(n_1252),
.B2(n_1299),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1277),
.B(n_1215),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1217),
.B(n_1312),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1295),
.A2(n_1309),
.B1(n_1320),
.B2(n_1270),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1309),
.B(n_1230),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1233),
.A2(n_1264),
.B(n_1271),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1320),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1310),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1239),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1240),
.B(n_1236),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1217),
.B(n_1308),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1226),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1226),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1273),
.A2(n_1241),
.B(n_1274),
.C(n_1249),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1241),
.A2(n_1274),
.B(n_1267),
.C(n_1268),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1274),
.A2(n_1230),
.B(n_1275),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1289),
.B(n_1321),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1230),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1288),
.A2(n_1313),
.B(n_1314),
.C(n_1321),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1230),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1310),
.A2(n_1325),
.B1(n_1292),
.B2(n_1322),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_1310),
.B(n_1325),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1322),
.A2(n_1275),
.B1(n_1231),
.B2(n_1221),
.Y(n_1388)
);

AOI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1275),
.A2(n_1284),
.B(n_1290),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1291),
.B(n_1301),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1296),
.B(n_1311),
.Y(n_1391)
);

OA22x2_ASAP7_75t_L g1392 ( 
.A1(n_1311),
.A2(n_1219),
.B1(n_1243),
.B2(n_1179),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1225),
.B(n_1286),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1279),
.A2(n_1167),
.B(n_832),
.C(n_965),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1215),
.B(n_1299),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1214),
.B(n_1223),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1306),
.Y(n_1397)
);

OA22x2_ASAP7_75t_L g1398 ( 
.A1(n_1219),
.A2(n_1243),
.B1(n_1179),
.B2(n_1173),
.Y(n_1398)
);

AOI221x1_ASAP7_75t_SL g1399 ( 
.A1(n_1237),
.A2(n_1119),
.B1(n_607),
.B2(n_853),
.C(n_447),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1280),
.A2(n_832),
.B1(n_1328),
.B2(n_1179),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1214),
.B(n_1223),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1281),
.A2(n_1167),
.B(n_1316),
.C(n_1294),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1280),
.A2(n_832),
.B1(n_1328),
.B2(n_1179),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1279),
.A2(n_1179),
.B(n_1173),
.C(n_832),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1214),
.B(n_1223),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1280),
.A2(n_832),
.B1(n_1328),
.B2(n_1179),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1280),
.A2(n_832),
.B1(n_1328),
.B2(n_1179),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1370),
.B(n_1383),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1391),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1389),
.A2(n_1388),
.B(n_1342),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1343),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1394),
.A2(n_1402),
.B(n_1404),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1350),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1404),
.A2(n_1407),
.B(n_1406),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1341),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1371),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1340),
.B(n_1333),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1332),
.B(n_1396),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1353),
.A2(n_1379),
.B(n_1380),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1401),
.B(n_1405),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1343),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1374),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1343),
.B(n_1395),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1400),
.A2(n_1403),
.B1(n_1330),
.B2(n_1398),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1385),
.B(n_1395),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1367),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1353),
.A2(n_1379),
.B(n_1380),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1337),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1395),
.B(n_1337),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1337),
.B(n_1361),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1338),
.A2(n_1346),
.B(n_1386),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1338),
.A2(n_1365),
.B(n_1390),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1361),
.B(n_1352),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1398),
.A2(n_1336),
.B1(n_1349),
.B2(n_1355),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1375),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1352),
.B(n_1375),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1363),
.A2(n_1366),
.B(n_1334),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1375),
.B(n_1359),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1334),
.A2(n_1369),
.B(n_1348),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_SL g1440 ( 
.A(n_1372),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1329),
.B(n_1347),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1372),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1399),
.A2(n_1392),
.B1(n_1357),
.B2(n_1331),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1339),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1392),
.B(n_1345),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1368),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1376),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1429),
.B(n_1344),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1416),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1447),
.B(n_1393),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_L g1451 ( 
.A(n_1410),
.B(n_1381),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1429),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1428),
.B(n_1354),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1413),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1413),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1447),
.B(n_1335),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_SL g1457 ( 
.A1(n_1412),
.A2(n_1424),
.B(n_1434),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1428),
.B(n_1358),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1435),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1422),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1409),
.B(n_1351),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1422),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1409),
.B(n_1433),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1409),
.B(n_1382),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1437),
.B(n_1384),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1446),
.B(n_1364),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1425),
.B(n_1436),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1438),
.B(n_1373),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1414),
.B(n_1435),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1360),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1408),
.B(n_1356),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_SL g1472 ( 
.A(n_1415),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1454),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1457),
.A2(n_1424),
.B1(n_1412),
.B2(n_1434),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1449),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1456),
.B(n_1417),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1457),
.A2(n_1417),
.B1(n_1439),
.B2(n_1431),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1454),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1453),
.B(n_1426),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1456),
.B(n_1442),
.C(n_1441),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1472),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1455),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1465),
.A2(n_1441),
.B(n_1443),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1460),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1472),
.A2(n_1443),
.B1(n_1418),
.B2(n_1420),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_1461),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1449),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1448),
.B(n_1423),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1460),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1462),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1469),
.A2(n_1439),
.B1(n_1431),
.B2(n_1437),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1449),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1465),
.A2(n_1431),
.B1(n_1439),
.B2(n_1437),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1469),
.A2(n_1418),
.B1(n_1420),
.B2(n_1440),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1448),
.B(n_1423),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1453),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1462),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1469),
.A2(n_1440),
.B1(n_1378),
.B2(n_1377),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1469),
.A2(n_1439),
.B1(n_1432),
.B2(n_1419),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1469),
.A2(n_1415),
.B1(n_1444),
.B2(n_1426),
.Y(n_1501)
);

OAI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1469),
.A2(n_1362),
.B1(n_1444),
.B2(n_1445),
.C(n_1421),
.Y(n_1502)
);

AOI31xp33_ASAP7_75t_L g1503 ( 
.A1(n_1471),
.A2(n_1445),
.A3(n_1377),
.B(n_1421),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1450),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1471),
.B(n_1408),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1471),
.B(n_1408),
.Y(n_1507)
);

OR2x6_ASAP7_75t_L g1508 ( 
.A(n_1469),
.B(n_1410),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1469),
.A2(n_1439),
.B1(n_1432),
.B2(n_1419),
.Y(n_1509)
);

NAND2x1_ASAP7_75t_SL g1510 ( 
.A(n_1484),
.B(n_1463),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1484),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1459),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1475),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1486),
.B(n_1467),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1473),
.Y(n_1515)
);

AOI211x1_ASAP7_75t_L g1516 ( 
.A1(n_1483),
.A2(n_1450),
.B(n_1466),
.C(n_1445),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1487),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1506),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1478),
.Y(n_1519)
);

NOR2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1480),
.B(n_1397),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1500),
.A2(n_1451),
.B(n_1430),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1504),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1499),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1507),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1482),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

AND2x6_ASAP7_75t_SL g1527 ( 
.A(n_1476),
.B(n_1378),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1491),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1481),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1504),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1481),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1488),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1494),
.A2(n_1427),
.B(n_1419),
.Y(n_1534)
);

AND2x6_ASAP7_75t_SL g1535 ( 
.A(n_1476),
.B(n_1362),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1497),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1488),
.Y(n_1537)
);

INVx4_ASAP7_75t_SL g1538 ( 
.A(n_1508),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1508),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1493),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1522),
.B(n_1489),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1516),
.B(n_1477),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1543)
);

AND3x1_ASAP7_75t_L g1544 ( 
.A(n_1527),
.B(n_1474),
.C(n_1535),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1518),
.B(n_1485),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1531),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1531),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1518),
.B(n_1505),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1522),
.B(n_1496),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1524),
.B(n_1479),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1535),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1530),
.B(n_1467),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1528),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1510),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1510),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1513),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1528),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1536),
.B(n_1505),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1531),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1513),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1512),
.B(n_1452),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1520),
.A2(n_1474),
.B1(n_1492),
.B2(n_1494),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1536),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1515),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1527),
.B(n_1448),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1520),
.A2(n_1509),
.B1(n_1500),
.B2(n_1495),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1512),
.B(n_1452),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_1470),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1515),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1519),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1513),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1464),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1529),
.B(n_1464),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1519),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1523),
.A2(n_1509),
.B1(n_1503),
.B2(n_1502),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1511),
.B(n_1470),
.Y(n_1577)
);

OAI33xp33_ASAP7_75t_L g1578 ( 
.A1(n_1525),
.A2(n_1495),
.A3(n_1501),
.B1(n_1466),
.B2(n_1470),
.B3(n_1458),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_L g1579 ( 
.A(n_1517),
.B(n_1501),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1544),
.B(n_1539),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1564),
.B(n_1526),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1565),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1553),
.B(n_1526),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1532),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1544),
.B(n_1539),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1541),
.B(n_1538),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1549),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1556),
.A2(n_1534),
.B(n_1521),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1551),
.B(n_1546),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1557),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1565),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1558),
.B(n_1532),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1538),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1533),
.Y(n_1594)
);

INVxp33_ASAP7_75t_L g1595 ( 
.A(n_1548),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1551),
.B(n_1534),
.C(n_1521),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1570),
.B(n_1533),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1570),
.B(n_1537),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1571),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1557),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1537),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1556),
.B(n_1554),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1561),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1560),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1575),
.B(n_1540),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1559),
.B(n_1514),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1560),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1561),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1561),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1547),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1575),
.B(n_1540),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1569),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1569),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1588),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1579),
.Y(n_1616)
);

AOI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1589),
.A2(n_1547),
.B(n_1543),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1586),
.B(n_1579),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1593),
.B(n_1562),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1593),
.B(n_1562),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1611),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1608),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1605),
.B(n_1542),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1580),
.A2(n_1563),
.B1(n_1576),
.B2(n_1567),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1596),
.A2(n_1545),
.B1(n_1566),
.B2(n_1574),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1587),
.B(n_1538),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1603),
.B(n_1568),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1603),
.B(n_1587),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1585),
.A2(n_1597),
.B(n_1590),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1611),
.B(n_1577),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1581),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1588),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1595),
.A2(n_1573),
.B1(n_1539),
.B2(n_1432),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1613),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1607),
.B(n_1550),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1588),
.B(n_1568),
.Y(n_1639)
);

AOI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1626),
.A2(n_1584),
.B(n_1592),
.Y(n_1640)
);

O2A1O1Ixp33_ASAP7_75t_SL g1641 ( 
.A1(n_1624),
.A2(n_1592),
.B(n_1584),
.C(n_1581),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1624),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_SL g1643 ( 
.A1(n_1617),
.A2(n_1594),
.B(n_1600),
.C(n_1591),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1637),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1631),
.B(n_1613),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1616),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1637),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1627),
.A2(n_1588),
.B1(n_1614),
.B2(n_1583),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1626),
.A2(n_1614),
.B1(n_1539),
.B2(n_1538),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1623),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1623),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1616),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1627),
.A2(n_1583),
.B1(n_1594),
.B2(n_1539),
.C(n_1598),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1631),
.B(n_1552),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1552),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1623),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1616),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1617),
.B(n_1582),
.C(n_1591),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1628),
.A2(n_1625),
.B1(n_1638),
.B2(n_1634),
.C(n_1618),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1657),
.B(n_1634),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1651),
.Y(n_1661)
);

OAI321xp33_ASAP7_75t_L g1662 ( 
.A1(n_1649),
.A2(n_1618),
.A3(n_1625),
.B1(n_1636),
.B2(n_1633),
.C(n_1630),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1645),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1619),
.Y(n_1664)
);

CKINVDCx6p67_ASAP7_75t_R g1665 ( 
.A(n_1642),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1646),
.B(n_1630),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1655),
.B(n_1619),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1652),
.B(n_1618),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1630),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1651),
.Y(n_1670)
);

NAND4xp75_ASAP7_75t_L g1671 ( 
.A(n_1669),
.B(n_1640),
.C(n_1656),
.D(n_1650),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1662),
.A2(n_1641),
.B1(n_1643),
.B2(n_1648),
.C(n_1653),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1663),
.A2(n_1641),
.B(n_1643),
.C(n_1658),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1660),
.A2(n_1648),
.B(n_1647),
.Y(n_1674)
);

AOI211xp5_ASAP7_75t_L g1675 ( 
.A1(n_1668),
.A2(n_1644),
.B(n_1620),
.C(n_1629),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1668),
.A2(n_1633),
.B1(n_1632),
.B2(n_1620),
.C(n_1619),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1665),
.B(n_1621),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1664),
.B(n_1621),
.Y(n_1678)
);

AOI221x1_ASAP7_75t_L g1679 ( 
.A1(n_1661),
.A2(n_1622),
.B1(n_1635),
.B2(n_1615),
.C(n_1629),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1677),
.B(n_1665),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1673),
.A2(n_1666),
.B1(n_1667),
.B2(n_1629),
.Y(n_1681)
);

NAND5xp2_ASAP7_75t_L g1682 ( 
.A(n_1672),
.B(n_1670),
.C(n_1621),
.D(n_1639),
.E(n_1632),
.Y(n_1682)
);

XOR2xp5_ASAP7_75t_L g1683 ( 
.A(n_1671),
.B(n_1629),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1678),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1680),
.B(n_1674),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1683),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1684),
.B(n_1675),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1681),
.B(n_1676),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1682),
.B(n_1629),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1684),
.B(n_1679),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1685),
.A2(n_1632),
.B1(n_1622),
.B2(n_1635),
.C(n_1615),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1686),
.A2(n_1632),
.B(n_1635),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1689),
.A2(n_1639),
.B(n_1622),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1687),
.B(n_1582),
.Y(n_1694)
);

XNOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1688),
.B(n_1397),
.Y(n_1695)
);

AOI322xp5_ASAP7_75t_L g1696 ( 
.A1(n_1694),
.A2(n_1690),
.A3(n_1622),
.B1(n_1615),
.B2(n_1639),
.C1(n_1600),
.C2(n_1604),
.Y(n_1696)
);

NOR3x1_ASAP7_75t_L g1697 ( 
.A(n_1693),
.B(n_1598),
.C(n_1602),
.Y(n_1697)
);

CKINVDCx16_ASAP7_75t_R g1698 ( 
.A(n_1695),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_SL g1699 ( 
.A(n_1698),
.B(n_1692),
.C(n_1691),
.Y(n_1699)
);

OAI211xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1699),
.A2(n_1696),
.B(n_1697),
.C(n_1601),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1700),
.A2(n_1590),
.B1(n_1610),
.B2(n_1609),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1700),
.B(n_1590),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1702),
.B(n_1597),
.Y(n_1703)
);

AOI21xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1701),
.A2(n_1597),
.B(n_1610),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1703),
.A2(n_1601),
.B(n_1610),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_SL g1706 ( 
.A1(n_1704),
.A2(n_1609),
.B1(n_1601),
.B2(n_1604),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1705),
.B(n_1604),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1707),
.A2(n_1706),
.B1(n_1609),
.B2(n_1612),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1606),
.B(n_1602),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1612),
.B1(n_1606),
.B2(n_1599),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1599),
.B1(n_1572),
.B2(n_1555),
.Y(n_1711)
);

AOI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1387),
.B(n_1572),
.C(n_1539),
.Y(n_1712)
);


endmodule