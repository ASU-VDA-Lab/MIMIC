module fake_ibex_1987_n_3139 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_658, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3139);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_658;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3139;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3105;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_1636;
wire n_939;
wire n_1687;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2846;
wire n_2685;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_2723;
wire n_1616;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2646;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_1395;
wire n_998;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_961;
wire n_991;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_3104;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_980;
wire n_1193;
wire n_849;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2148;
wire n_949;
wire n_704;
wire n_2104;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_267),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_417),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_48),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_317),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_237),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_405),
.Y(n_669)
);

CKINVDCx14_ASAP7_75t_R g670 ( 
.A(n_470),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_235),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_273),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_246),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_658),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_47),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_77),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_552),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_486),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_77),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_363),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_483),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_162),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_115),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_126),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_200),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_235),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_472),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_98),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_551),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_412),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_602),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_449),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_144),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_344),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_586),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_598),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_123),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_534),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_628),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_489),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_371),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_534),
.Y(n_702)
);

CKINVDCx14_ASAP7_75t_R g703 ( 
.A(n_596),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_3),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_547),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_186),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_149),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_374),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_656),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_146),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_634),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_194),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_248),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_549),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_92),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_127),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_396),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_491),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_589),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_274),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_67),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_73),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_617),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_497),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_281),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_378),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_560),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_190),
.Y(n_728)
);

INVx4_ASAP7_75t_R g729 ( 
.A(n_655),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_83),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_265),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_291),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_574),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_315),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_29),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_48),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_228),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_143),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_335),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_59),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_228),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_501),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_196),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_303),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_613),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_281),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_564),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_445),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_113),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_398),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_610),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_413),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_527),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_258),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_620),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_146),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_645),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_188),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_392),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_288),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_568),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_265),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_149),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_252),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_70),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_341),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_161),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_153),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_88),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_23),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_524),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_657),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_258),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_240),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_465),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_173),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_379),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_469),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_352),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_614),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_466),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_590),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_388),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_293),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_279),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_653),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_322),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_449),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_477),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_260),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_61),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_547),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_619),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_188),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_663),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_129),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_489),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_22),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_40),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_271),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_564),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_384),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_608),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_508),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_343),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_375),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_137),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_520),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_633),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_539),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_360),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_403),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_300),
.Y(n_814)
);

CKINVDCx16_ASAP7_75t_R g815 ( 
.A(n_213),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_623),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_543),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_197),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_618),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_487),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_135),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_296),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_147),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_636),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_136),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_557),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_192),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_287),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_371),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_71),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_13),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_573),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_51),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_626),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_212),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_142),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_408),
.Y(n_837)
);

CKINVDCx14_ASAP7_75t_R g838 ( 
.A(n_124),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_322),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_68),
.Y(n_840)
);

INVxp33_ASAP7_75t_R g841 ( 
.A(n_219),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_304),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_39),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_240),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_276),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_62),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_186),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_182),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_116),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_503),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_12),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_347),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_269),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_287),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_652),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_320),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_316),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_6),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_60),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_368),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_462),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_144),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_600),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_528),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_430),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_294),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_638),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_168),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_412),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_587),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_276),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_515),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_261),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_585),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_65),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_137),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_518),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_30),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_94),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_649),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_436),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_470),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_364),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_330),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_551),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_298),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_58),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_185),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_318),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_642),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_109),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_659),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_27),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_402),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_124),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_210),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_64),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_171),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_79),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_426),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_329),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_392),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_251),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_382),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_430),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_589),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_13),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_327),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_108),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_346),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_305),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_211),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_382),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_593),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_478),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_400),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_374),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_140),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_278),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_152),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_661),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_579),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_458),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_625),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_573),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_390),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_413),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_64),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_588),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_611),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_651),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_57),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_601),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_138),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_539),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_447),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_85),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_459),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_225),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_454),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_288),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_566),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_365),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_495),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_294),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_581),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_174),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_121),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_615),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_562),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_538),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_92),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_97),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_548),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_179),
.Y(n_955)
);

BUFx5_ASAP7_75t_L g956 ( 
.A(n_234),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_400),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_575),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_290),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_109),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_190),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_90),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_511),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_296),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_203),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_343),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_313),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_262),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_517),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_120),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_195),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_485),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_604),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_532),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_465),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_59),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_662),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_369),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_641),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_233),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_567),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_493),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_175),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_518),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_148),
.Y(n_985)
);

CKINVDCx16_ASAP7_75t_R g986 ( 
.A(n_174),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_378),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_69),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_479),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_167),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_321),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_219),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_444),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_425),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_558),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_128),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_71),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_527),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_14),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_208),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_650),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_168),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_200),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_159),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_603),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_2),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_578),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_277),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_358),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_25),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_380),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_632),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_275),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_492),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_212),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_488),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_191),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_46),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_445),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_182),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_555),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_441),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_612),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_504),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_338),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_494),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_377),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_38),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_55),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_577),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_229),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_243),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_598),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_424),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_631),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_509),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_648),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_29),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_119),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_615),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_428),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_166),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_131),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_291),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_654),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_365),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_603),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_411),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_204),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_39),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_660),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_443),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_218),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_70),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_431),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_646),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_187),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_787),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_978),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_711),
.B(n_0),
.Y(n_1060)
);

CKINVDCx16_ASAP7_75t_R g1061 ( 
.A(n_815),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_978),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1035),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_688),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_734),
.B(n_0),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_978),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_736),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_808),
.Y(n_1068)
);

INVxp33_ASAP7_75t_SL g1069 ( 
.A(n_788),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_670),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_711),
.B(n_1),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_703),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_838),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_840),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_808),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_809),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_674),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_739),
.B(n_1),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_809),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_951),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_986),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_956),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_699),
.B(n_2),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_665),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_723),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_821),
.B(n_917),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_917),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_667),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_880),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_935),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_935),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_956),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_867),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_867),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1045),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_675),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1045),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_974),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_681),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_682),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_816),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_826),
.Y(n_1102)
);

INVxp33_ASAP7_75t_SL g1103 ( 
.A(n_913),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1051),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1051),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_696),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_747),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_747),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_797),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_698),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_664),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_664),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_666),
.Y(n_1113)
);

CKINVDCx16_ASAP7_75t_R g1114 ( 
.A(n_712),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_797),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_666),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_823),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_816),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_669),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_835),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_669),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_673),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_853),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_894),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_894),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_709),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_904),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_770),
.B(n_4),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_904),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_676),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_733),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_908),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_740),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_676),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_744),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_819),
.B(n_824),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_750),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_678),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_914),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_759),
.Y(n_1140)
);

CKINVDCx16_ASAP7_75t_R g1141 ( 
.A(n_712),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_680),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_918),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_962),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_680),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_789),
.Y(n_1146)
);

CKINVDCx16_ASAP7_75t_R g1147 ( 
.A(n_789),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_683),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_777),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_791),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_683),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_921),
.B(n_5),
.Y(n_1152)
);

INVxp33_ASAP7_75t_SL g1153 ( 
.A(n_687),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_950),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_687),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_950),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_960),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_689),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1067),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1082),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1089),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1101),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1089),
.B(n_980),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_1077),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1068),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1075),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1076),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1102),
.B(n_789),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1079),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1082),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1069),
.A2(n_690),
.B1(n_691),
.B2(n_689),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1062),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1086),
.B(n_980),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1107),
.B(n_924),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1066),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1092),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1087),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1090),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1091),
.B(n_1010),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1098),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1144),
.B(n_850),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1129),
.B(n_1001),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1118),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1139),
.B(n_1012),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1126),
.B(n_1037),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1065),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1108),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1109),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1115),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1117),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1120),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1126),
.B(n_1056),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1078),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1123),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1124),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1125),
.B(n_956),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1060),
.A2(n_684),
.B(n_671),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1127),
.B(n_956),
.Y(n_1198)
);

AND2x6_ASAP7_75t_L g1199 ( 
.A(n_1071),
.B(n_931),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1132),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1143),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1146),
.B(n_964),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1158),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1064),
.B(n_1010),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1154),
.B(n_956),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1156),
.B(n_956),
.Y(n_1206)
);

AND2x6_ASAP7_75t_L g1207 ( 
.A(n_1136),
.B(n_931),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1157),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1128),
.A2(n_684),
.B(n_671),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1152),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1083),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1112),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1103),
.B(n_956),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1113),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1114),
.A2(n_1050),
.B1(n_1048),
.B2(n_814),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1085),
.A2(n_765),
.B(n_710),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1093),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1094),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1095),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1097),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1116),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1104),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1105),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1119),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1070),
.B(n_668),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1121),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1122),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1130),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1134),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1138),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1142),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1145),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1148),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1151),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1155),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1072),
.B(n_1011),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1153),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1141),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1147),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1061),
.B(n_975),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1073),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1058),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1074),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1080),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1080),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1063),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1081),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1081),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1088),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1096),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1099),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1084),
.B(n_931),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1100),
.B(n_755),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1106),
.B(n_850),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1106),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1110),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1131),
.B(n_1011),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1131),
.B(n_952),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1133),
.B(n_710),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1135),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1135),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1137),
.B(n_765),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1137),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1140),
.A2(n_822),
.B1(n_843),
.B2(n_805),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1140),
.A2(n_851),
.B1(n_879),
.B2(n_864),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1149),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1150),
.B(n_931),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1067),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1082),
.Y(n_1269)
);

XOR2xp5_ASAP7_75t_L g1270 ( 
.A(n_1080),
.B(n_884),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1082),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_SL g1272 ( 
.A(n_1078),
.B(n_668),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1089),
.B(n_785),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1082),
.A2(n_792),
.B(n_785),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_1114),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1067),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1102),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1059),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1067),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1107),
.B(n_757),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1059),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1059),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1101),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1059),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1101),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1082),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1089),
.B(n_792),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1082),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1082),
.A2(n_875),
.B(n_856),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1059),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1082),
.A2(n_875),
.B(n_856),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1067),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1101),
.Y(n_1293)
);

NAND2x1_ASAP7_75t_L g1294 ( 
.A(n_1078),
.B(n_729),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1102),
.B(n_952),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1067),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1059),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1059),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1067),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1067),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1059),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1067),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1102),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1082),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1059),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1084),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1082),
.B(n_794),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1067),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1082),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1067),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1102),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1082),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1107),
.B(n_773),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1107),
.B(n_796),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1059),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1101),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1102),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1111),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1102),
.B(n_952),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1101),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1077),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1107),
.B(n_810),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1111),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1101),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1084),
.A2(n_885),
.B1(n_919),
.B2(n_910),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1067),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1067),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1210),
.B(n_1211),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1274),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1161),
.B(n_794),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1274),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1280),
.B(n_834),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1216),
.A2(n_672),
.B1(n_679),
.B2(n_677),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1207),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1210),
.B(n_794),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1277),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1183),
.Y(n_1337)
);

AND2x6_ASAP7_75t_L g1338 ( 
.A(n_1217),
.B(n_947),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1289),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1289),
.Y(n_1340)
);

AO22x2_ASAP7_75t_L g1341 ( 
.A1(n_1215),
.A2(n_841),
.B1(n_741),
.B2(n_746),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1180),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1162),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1226),
.B(n_685),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1303),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1303),
.B(n_693),
.Y(n_1346)
);

AND3x1_ASAP7_75t_L g1347 ( 
.A(n_1247),
.B(n_692),
.C(n_686),
.Y(n_1347)
);

AND2x6_ASAP7_75t_L g1348 ( 
.A(n_1217),
.B(n_947),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1311),
.B(n_727),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1186),
.B(n_1227),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1164),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1311),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1208),
.Y(n_1353)
);

INVxp33_ASAP7_75t_SL g1354 ( 
.A(n_1317),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1162),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1283),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1283),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1280),
.B(n_855),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1275),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1285),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1186),
.B(n_1228),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1317),
.B(n_727),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1285),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1230),
.B(n_890),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1313),
.B(n_892),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1314),
.B(n_977),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1314),
.B(n_979),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1291),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1291),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1293),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1232),
.B(n_694),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1293),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1316),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1316),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1320),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1320),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1207),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1324),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1324),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1171),
.B(n_1319),
.Y(n_1380)
);

AND2x6_ASAP7_75t_L g1381 ( 
.A(n_1220),
.B(n_1017),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1168),
.B(n_700),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1210),
.B(n_668),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1159),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1295),
.B(n_700),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1165),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1193),
.B(n_714),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1216),
.A2(n_695),
.B1(n_702),
.B2(n_697),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1166),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1163),
.B(n_705),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1210),
.A2(n_707),
.B1(n_716),
.B2(n_706),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1167),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1169),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1213),
.B(n_668),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1163),
.B(n_718),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1214),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1207),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1322),
.B(n_704),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1181),
.B(n_713),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1177),
.Y(n_1400)
);

INVx4_ASAP7_75t_SL g1401 ( 
.A(n_1207),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1306),
.A2(n_955),
.B1(n_965),
.B2(n_927),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1224),
.B(n_721),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1318),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_1238),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1178),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1323),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1196),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1203),
.Y(n_1409)
);

AND2x6_ASAP7_75t_L g1410 ( 
.A(n_1220),
.B(n_1017),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1207),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1321),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1231),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1321),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1253),
.B(n_708),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1253),
.B(n_713),
.Y(n_1416)
);

BUFx10_ASAP7_75t_L g1417 ( 
.A(n_1239),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1326),
.Y(n_1418)
);

AND3x2_ASAP7_75t_L g1419 ( 
.A(n_1263),
.B(n_1004),
.C(n_973),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1220),
.B(n_720),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1174),
.B(n_1182),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1244),
.B(n_715),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1197),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1198),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1198),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1251),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1229),
.B(n_701),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1212),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1254),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1205),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1205),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1206),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1174),
.B(n_717),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1234),
.B(n_701),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1221),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1231),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1235),
.B(n_735),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1182),
.B(n_719),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1221),
.B(n_725),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1206),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1209),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1233),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1170),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1202),
.B(n_737),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1272),
.B(n_725),
.C(n_722),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1251),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1170),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1184),
.B(n_726),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1218),
.B(n_724),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1172),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1219),
.B(n_742),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1201),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1179),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1160),
.Y(n_1454)
);

AND2x2_ASAP7_75t_SL g1455 ( 
.A(n_1258),
.B(n_1042),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1223),
.B(n_751),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1272),
.A2(n_752),
.B1(n_760),
.B2(n_758),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1236),
.B(n_701),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1265),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1204),
.B(n_730),
.Y(n_1460)
);

AND2x6_ASAP7_75t_L g1461 ( 
.A(n_1220),
.B(n_701),
.Y(n_1461)
);

AND2x6_ASAP7_75t_L g1462 ( 
.A(n_1222),
.B(n_756),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1233),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1170),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1237),
.B(n_761),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1184),
.B(n_726),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_SL g1467 ( 
.A(n_1242),
.B(n_728),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1204),
.B(n_1192),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1175),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1233),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1247),
.B(n_763),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1268),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1257),
.B(n_732),
.Y(n_1473)
);

INVx5_ASAP7_75t_L g1474 ( 
.A(n_1269),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1294),
.B(n_738),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1325),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1278),
.Y(n_1477)
);

AND2x2_ASAP7_75t_SL g1478 ( 
.A(n_1257),
.B(n_1055),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1276),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1279),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1292),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1192),
.B(n_728),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1246),
.A2(n_1245),
.B1(n_1248),
.B2(n_1243),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1273),
.B(n_1008),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1222),
.B(n_756),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1270),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1269),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1296),
.B(n_1299),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1250),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1281),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1273),
.B(n_1008),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1300),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1282),
.Y(n_1493)
);

INVx6_ASAP7_75t_L g1494 ( 
.A(n_1287),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1302),
.B(n_731),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1287),
.B(n_999),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1269),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1308),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1264),
.A2(n_866),
.B1(n_997),
.B2(n_732),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1250),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1310),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1269),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1173),
.B(n_764),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1327),
.B(n_866),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1307),
.B(n_756),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1284),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1249),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1290),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1297),
.Y(n_1509)
);

BUFx4f_ASAP7_75t_L g1510 ( 
.A(n_1259),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1298),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1301),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1199),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1199),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1305),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1307),
.B(n_997),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1199),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1315),
.Y(n_1518)
);

AND2x6_ASAP7_75t_L g1519 ( 
.A(n_1187),
.B(n_756),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1271),
.Y(n_1520)
);

AND2x6_ASAP7_75t_L g1521 ( 
.A(n_1188),
.B(n_756),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1189),
.B(n_836),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1185),
.B(n_1000),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1240),
.A2(n_1002),
.B1(n_1005),
.B2(n_1000),
.Y(n_1524)
);

BUFx10_ASAP7_75t_L g1525 ( 
.A(n_1259),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1190),
.B(n_1191),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1199),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1271),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1262),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1194),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1249),
.Y(n_1531)
);

BUFx10_ASAP7_75t_L g1532 ( 
.A(n_1262),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1195),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1252),
.B(n_769),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1200),
.B(n_1002),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1160),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1176),
.B(n_1006),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1384),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1421),
.B(n_1468),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1386),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1354),
.A2(n_1267),
.B1(n_1022),
.B2(n_1241),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1359),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1482),
.B(n_1006),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1389),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1392),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1393),
.Y(n_1546)
);

OAI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1524),
.A2(n_1225),
.B1(n_1255),
.B2(n_1260),
.C(n_1256),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1536),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1400),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1406),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1345),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1336),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1351),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1408),
.B(n_1007),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1472),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1479),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1480),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1407),
.B(n_1412),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1352),
.A2(n_1013),
.B1(n_1014),
.B2(n_1007),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1536),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1341),
.A2(n_1261),
.B1(n_1266),
.B2(n_1029),
.Y(n_1561)
);

AO22x2_ASAP7_75t_L g1562 ( 
.A1(n_1441),
.A2(n_825),
.B1(n_849),
.B2(n_799),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1408),
.B(n_1013),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1481),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1412),
.B(n_1261),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1492),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1529),
.A2(n_1018),
.B1(n_1023),
.B2(n_1016),
.C(n_1014),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1414),
.B(n_772),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_1396),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1414),
.B(n_778),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1498),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1423),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1501),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1346),
.B(n_1018),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1344),
.B(n_781),
.Y(n_1575)
);

NAND3x1_ASAP7_75t_L g1576 ( 
.A(n_1402),
.B(n_783),
.C(n_782),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1435),
.B(n_1404),
.Y(n_1577)
);

AO22x2_ASAP7_75t_L g1578 ( 
.A1(n_1329),
.A2(n_793),
.B1(n_795),
.B2(n_790),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1349),
.B(n_1023),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1344),
.B(n_800),
.Y(n_1580)
);

AO22x2_ASAP7_75t_L g1581 ( 
.A1(n_1329),
.A2(n_807),
.B1(n_817),
.B2(n_804),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1409),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1530),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1382),
.B(n_1024),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1533),
.Y(n_1585)
);

OAI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1510),
.A2(n_1025),
.B1(n_1026),
.B2(n_1024),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1533),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1362),
.B(n_1025),
.Y(n_1588)
);

AO22x2_ASAP7_75t_L g1589 ( 
.A1(n_1331),
.A2(n_820),
.B1(n_827),
.B2(n_818),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1424),
.A2(n_1028),
.B1(n_1029),
.B2(n_1027),
.Y(n_1590)
);

AO22x2_ASAP7_75t_L g1591 ( 
.A1(n_1331),
.A2(n_830),
.B1(n_839),
.B2(n_828),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1467),
.B(n_1028),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1424),
.B(n_1030),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1428),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1425),
.B(n_1030),
.Y(n_1595)
);

AO22x2_ASAP7_75t_L g1596 ( 
.A1(n_1339),
.A2(n_847),
.B1(n_854),
.B2(n_842),
.Y(n_1596)
);

AO22x2_ASAP7_75t_L g1597 ( 
.A1(n_1339),
.A2(n_860),
.B1(n_862),
.B2(n_859),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1387),
.B(n_1031),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1380),
.A2(n_1033),
.B1(n_1036),
.B2(n_1032),
.C(n_1031),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1371),
.B(n_865),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1489),
.Y(n_1601)
);

AO22x2_ASAP7_75t_L g1602 ( 
.A1(n_1340),
.A2(n_870),
.B1(n_873),
.B2(n_869),
.Y(n_1602)
);

CKINVDCx14_ASAP7_75t_R g1603 ( 
.A(n_1500),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_SL g1604 ( 
.A(n_1471),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1439),
.Y(n_1605)
);

NAND3xp33_ASAP7_75t_SL g1606 ( 
.A(n_1426),
.B(n_1036),
.C(n_1033),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1350),
.A2(n_1039),
.B1(n_1040),
.B2(n_1038),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1471),
.B(n_882),
.Y(n_1608)
);

OAI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1429),
.A2(n_1510),
.B1(n_1361),
.B2(n_1416),
.C(n_1415),
.Y(n_1609)
);

AO22x2_ASAP7_75t_L g1610 ( 
.A1(n_1340),
.A2(n_886),
.B1(n_888),
.B2(n_883),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1385),
.B(n_1038),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1453),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1422),
.A2(n_1041),
.B1(n_1047),
.B2(n_1040),
.C(n_1039),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1425),
.B(n_1041),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1430),
.B(n_1049),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1433),
.A2(n_1053),
.B1(n_1054),
.B2(n_1052),
.C(n_1049),
.Y(n_1616)
);

NAND2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1347),
.B(n_889),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1453),
.Y(n_1618)
);

AO22x2_ASAP7_75t_L g1619 ( 
.A1(n_1368),
.A2(n_896),
.B1(n_898),
.B2(n_891),
.Y(n_1619)
);

AO22x2_ASAP7_75t_L g1620 ( 
.A1(n_1368),
.A2(n_923),
.B1(n_925),
.B2(n_899),
.Y(n_1620)
);

AO22x2_ASAP7_75t_L g1621 ( 
.A1(n_1369),
.A2(n_934),
.B1(n_937),
.B2(n_928),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1488),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1342),
.Y(n_1623)
);

AO22x2_ASAP7_75t_L g1624 ( 
.A1(n_1369),
.A2(n_945),
.B1(n_946),
.B2(n_944),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1450),
.Y(n_1625)
);

NAND2x1p5_ASAP7_75t_L g1626 ( 
.A(n_1436),
.B(n_957),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1399),
.A2(n_745),
.B1(n_748),
.B2(n_743),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1413),
.Y(n_1628)
);

AO22x2_ASAP7_75t_L g1629 ( 
.A1(n_1534),
.A2(n_1341),
.B1(n_1499),
.B2(n_1371),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1490),
.Y(n_1630)
);

NAND2x1p5_ASAP7_75t_L g1631 ( 
.A(n_1436),
.B(n_959),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1506),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1403),
.B(n_967),
.Y(n_1633)
);

AO22x2_ASAP7_75t_L g1634 ( 
.A1(n_1534),
.A2(n_982),
.B1(n_983),
.B2(n_981),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1508),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1405),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1477),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1431),
.B(n_749),
.Y(n_1638)
);

AO22x2_ASAP7_75t_L g1639 ( 
.A1(n_1473),
.A2(n_989),
.B1(n_1003),
.B2(n_984),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1403),
.A2(n_754),
.B1(n_762),
.B2(n_753),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1442),
.B(n_1009),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1509),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1512),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1432),
.B(n_766),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1515),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1518),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1449),
.A2(n_1456),
.B1(n_1451),
.B2(n_1444),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1449),
.A2(n_768),
.B1(n_771),
.B2(n_767),
.Y(n_1648)
);

AO22x2_ASAP7_75t_L g1649 ( 
.A1(n_1390),
.A2(n_1019),
.B1(n_1020),
.B2(n_1015),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1469),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1478),
.B(n_774),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1440),
.B(n_775),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1493),
.Y(n_1653)
);

CKINVDCx11_ASAP7_75t_R g1654 ( 
.A(n_1405),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1511),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1440),
.A2(n_1034),
.B1(n_1046),
.B2(n_1021),
.Y(n_1656)
);

CKINVDCx16_ASAP7_75t_R g1657 ( 
.A(n_1417),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1333),
.A2(n_1057),
.B1(n_779),
.B2(n_780),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1452),
.Y(n_1659)
);

AO22x2_ASAP7_75t_L g1660 ( 
.A1(n_1390),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1455),
.B(n_776),
.Y(n_1661)
);

AO22x2_ASAP7_75t_L g1662 ( 
.A1(n_1395),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1460),
.Y(n_1663)
);

AO22x2_ASAP7_75t_L g1664 ( 
.A1(n_1395),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1417),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1494),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1494),
.Y(n_1667)
);

OR2x2_ASAP7_75t_SL g1668 ( 
.A(n_1486),
.B(n_836),
.Y(n_1668)
);

AO22x2_ASAP7_75t_L g1669 ( 
.A1(n_1503),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1669)
);

CKINVDCx14_ASAP7_75t_R g1670 ( 
.A(n_1446),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1438),
.B(n_784),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1484),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1448),
.B(n_786),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1526),
.Y(n_1674)
);

AO22x2_ASAP7_75t_L g1675 ( 
.A1(n_1503),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1537),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1328),
.Y(n_1677)
);

AO22x2_ASAP7_75t_L g1678 ( 
.A1(n_1491),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1678)
);

AO22x2_ASAP7_75t_L g1679 ( 
.A1(n_1496),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1343),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1466),
.B(n_798),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1459),
.A2(n_802),
.B1(n_803),
.B2(n_801),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1355),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1356),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1357),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1334),
.B(n_1286),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1465),
.A2(n_811),
.B1(n_812),
.B2(n_806),
.Y(n_1687)
);

AO22x2_ASAP7_75t_L g1688 ( 
.A1(n_1419),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1360),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1363),
.Y(n_1690)
);

AO22x2_ASAP7_75t_L g1691 ( 
.A1(n_1445),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1525),
.B(n_813),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1372),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1525),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1373),
.Y(n_1695)
);

AO22x2_ASAP7_75t_L g1696 ( 
.A1(n_1458),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1374),
.Y(n_1697)
);

AO22x2_ASAP7_75t_L g1698 ( 
.A1(n_1401),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1375),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1507),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1376),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1379),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1418),
.Y(n_1703)
);

AO22x2_ASAP7_75t_L g1704 ( 
.A1(n_1401),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1531),
.Y(n_1705)
);

AO22x2_ASAP7_75t_L g1706 ( 
.A1(n_1398),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1483),
.B(n_829),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1532),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1495),
.Y(n_1709)
);

NAND2x1p5_ASAP7_75t_L g1710 ( 
.A(n_1463),
.B(n_1470),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1504),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1338),
.A2(n_832),
.B1(n_833),
.B2(n_831),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1535),
.Y(n_1713)
);

HAxp5_ASAP7_75t_SL g1714 ( 
.A(n_1476),
.B(n_31),
.CON(n_1714),
.SN(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1475),
.B(n_837),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1454),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_L g1717 ( 
.A(n_1348),
.B(n_1288),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1420),
.B(n_837),
.Y(n_1718)
);

AO22x2_ASAP7_75t_L g1719 ( 
.A1(n_1335),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1348),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1348),
.Y(n_1721)
);

AO22x2_ASAP7_75t_L g1722 ( 
.A1(n_1514),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1388),
.A2(n_844),
.B1(n_846),
.B2(n_845),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1514),
.B(n_837),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_L g1725 ( 
.A(n_1377),
.B(n_1288),
.Y(n_1725)
);

AO22x2_ASAP7_75t_L g1726 ( 
.A1(n_1527),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1332),
.B(n_1358),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1381),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1370),
.Y(n_1729)
);

AO22x2_ASAP7_75t_L g1730 ( 
.A1(n_1527),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1370),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1378),
.B(n_900),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1523),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1516),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1394),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1381),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_L g1737 ( 
.A(n_1377),
.B(n_1288),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1391),
.A2(n_857),
.B1(n_858),
.B2(n_852),
.C(n_848),
.Y(n_1738)
);

AO22x2_ASAP7_75t_L g1739 ( 
.A1(n_1513),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_1739)
);

AND2x6_ASAP7_75t_SL g1740 ( 
.A(n_1437),
.B(n_861),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1457),
.A2(n_871),
.B1(n_872),
.B2(n_868),
.C(n_863),
.Y(n_1741)
);

AO22x2_ASAP7_75t_L g1742 ( 
.A1(n_1517),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1505),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1381),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1427),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1434),
.Y(n_1747)
);

AO22x2_ASAP7_75t_L g1748 ( 
.A1(n_1367),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1330),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1410),
.Y(n_1750)
);

AO22x2_ASAP7_75t_L g1751 ( 
.A1(n_1410),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1522),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1383),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1485),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1364),
.B(n_874),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1353),
.Y(n_1756)
);

AO22x2_ASAP7_75t_L g1757 ( 
.A1(n_1337),
.A2(n_49),
.B1(n_45),
.B2(n_47),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1397),
.A2(n_877),
.B1(n_878),
.B2(n_876),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1353),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_1397),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1461),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_L g1762 ( 
.A(n_1411),
.B(n_1461),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1411),
.B(n_881),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1657),
.B(n_1411),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1552),
.B(n_1443),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1569),
.B(n_887),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1594),
.B(n_1443),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1539),
.B(n_893),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1760),
.B(n_895),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1636),
.B(n_1474),
.Y(n_1770)
);

NAND2xp33_ASAP7_75t_SL g1771 ( 
.A(n_1604),
.B(n_897),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1665),
.B(n_1474),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1601),
.B(n_1474),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1577),
.B(n_1520),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1582),
.B(n_1520),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1744),
.B(n_901),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1647),
.B(n_1520),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1551),
.B(n_902),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1559),
.B(n_903),
.Y(n_1779)
);

NAND2xp33_ASAP7_75t_SL g1780 ( 
.A(n_1750),
.B(n_905),
.Y(n_1780)
);

NAND2xp33_ASAP7_75t_SL g1781 ( 
.A(n_1750),
.B(n_906),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1712),
.B(n_907),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1590),
.B(n_909),
.Y(n_1783)
);

NAND2xp33_ASAP7_75t_SL g1784 ( 
.A(n_1721),
.B(n_911),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1694),
.B(n_912),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1758),
.B(n_915),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1700),
.B(n_916),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_SL g1788 ( 
.A(n_1720),
.B(n_920),
.Y(n_1788)
);

NAND2xp33_ASAP7_75t_SL g1789 ( 
.A(n_1727),
.B(n_922),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1705),
.B(n_926),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1574),
.B(n_929),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1583),
.B(n_1585),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1579),
.B(n_930),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1587),
.B(n_932),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1588),
.B(n_933),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1553),
.B(n_936),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1605),
.B(n_938),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1640),
.B(n_939),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1648),
.B(n_940),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1745),
.B(n_941),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1554),
.B(n_942),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1563),
.B(n_943),
.Y(n_1803)
);

NAND2xp33_ASAP7_75t_SL g1804 ( 
.A(n_1593),
.B(n_948),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1709),
.B(n_949),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1595),
.B(n_953),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1538),
.B(n_1528),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1614),
.B(n_954),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1615),
.B(n_958),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1708),
.B(n_1611),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1598),
.B(n_961),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1541),
.B(n_963),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1711),
.B(n_1713),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1626),
.B(n_966),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1631),
.B(n_968),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1540),
.B(n_969),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1641),
.B(n_970),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1716),
.B(n_971),
.Y(n_1818)
);

NAND2xp33_ASAP7_75t_SL g1819 ( 
.A(n_1638),
.B(n_972),
.Y(n_1819)
);

NAND2xp33_ASAP7_75t_SL g1820 ( 
.A(n_1644),
.B(n_976),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1627),
.B(n_985),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1652),
.B(n_987),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1544),
.B(n_988),
.Y(n_1823)
);

NAND2xp33_ASAP7_75t_SL g1824 ( 
.A(n_1572),
.B(n_990),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1607),
.B(n_991),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1584),
.B(n_992),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1692),
.B(n_1548),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1560),
.B(n_993),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1545),
.B(n_994),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1633),
.B(n_995),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1633),
.B(n_996),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1546),
.B(n_1462),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1676),
.B(n_1447),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1592),
.B(n_1628),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1555),
.B(n_1464),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1556),
.B(n_1487),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1557),
.B(n_1487),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1736),
.B(n_1497),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1568),
.B(n_1570),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1609),
.B(n_1502),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1617),
.B(n_1502),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1575),
.B(n_1580),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1575),
.B(n_1304),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1580),
.B(n_1304),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1600),
.B(n_1304),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1564),
.B(n_998),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1566),
.B(n_1309),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1723),
.B(n_1312),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1571),
.B(n_998),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1663),
.B(n_1672),
.Y(n_1851)
);

XNOR2xp5_ASAP7_75t_L g1852 ( 
.A(n_1629),
.B(n_49),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1651),
.B(n_1312),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1573),
.B(n_1734),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1661),
.B(n_998),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_SL g1856 ( 
.A(n_1749),
.B(n_1043),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1634),
.B(n_1043),
.Y(n_1857)
);

NAND2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1654),
.B(n_1043),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1687),
.B(n_1044),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1733),
.B(n_1519),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1625),
.B(n_1519),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1707),
.B(n_1521),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1543),
.B(n_1521),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1634),
.B(n_50),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1561),
.B(n_50),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1729),
.B(n_52),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1731),
.B(n_52),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1639),
.B(n_53),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1639),
.B(n_54),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1658),
.B(n_54),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1542),
.B(n_1565),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1623),
.B(n_55),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1578),
.B(n_56),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1763),
.B(n_57),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1671),
.B(n_58),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1673),
.B(n_61),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1632),
.B(n_62),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1681),
.B(n_63),
.Y(n_1878)
);

NAND2xp33_ASAP7_75t_SL g1879 ( 
.A(n_1630),
.B(n_63),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1715),
.B(n_65),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1715),
.B(n_66),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1682),
.B(n_66),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1635),
.B(n_67),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1710),
.B(n_72),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1732),
.B(n_74),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1732),
.B(n_75),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1656),
.B(n_75),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1578),
.B(n_76),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1642),
.B(n_78),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1581),
.B(n_78),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1643),
.B(n_79),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1645),
.B(n_80),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1646),
.B(n_80),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1724),
.B(n_81),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1581),
.B(n_81),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1724),
.B(n_82),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1650),
.B(n_82),
.Y(n_1897)
);

NAND2xp33_ASAP7_75t_SL g1898 ( 
.A(n_1653),
.B(n_84),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1655),
.B(n_86),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1589),
.B(n_86),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1659),
.B(n_87),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1589),
.B(n_89),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1666),
.B(n_89),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1667),
.B(n_90),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1755),
.B(n_91),
.Y(n_1905)
);

NAND2xp33_ASAP7_75t_SL g1906 ( 
.A(n_1637),
.B(n_93),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1591),
.B(n_95),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1674),
.B(n_95),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1703),
.B(n_96),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1591),
.B(n_96),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1699),
.B(n_99),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_SL g1912 ( 
.A(n_1701),
.B(n_100),
.Y(n_1912)
);

NAND2xp33_ASAP7_75t_SL g1913 ( 
.A(n_1702),
.B(n_100),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1612),
.B(n_101),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1618),
.B(n_101),
.Y(n_1915)
);

NAND2xp33_ASAP7_75t_SL g1916 ( 
.A(n_1608),
.B(n_102),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1596),
.B(n_103),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1597),
.B(n_103),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1608),
.B(n_104),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1680),
.B(n_105),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1683),
.B(n_105),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1684),
.B(n_106),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1685),
.B(n_106),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1602),
.B(n_107),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1689),
.B(n_108),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1668),
.B(n_1690),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1693),
.B(n_110),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1610),
.B(n_111),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1695),
.B(n_112),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1697),
.B(n_112),
.Y(n_1931)
);

NAND2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1677),
.B(n_113),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1718),
.B(n_114),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1619),
.B(n_114),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1756),
.B(n_115),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1759),
.B(n_116),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1735),
.B(n_117),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1603),
.B(n_118),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1743),
.B(n_118),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1746),
.B(n_1747),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1718),
.B(n_120),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1753),
.B(n_1754),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1619),
.B(n_122),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1620),
.B(n_1624),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1620),
.B(n_122),
.Y(n_1945)
);

NAND2xp33_ASAP7_75t_SL g1946 ( 
.A(n_1761),
.B(n_125),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1752),
.B(n_126),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1621),
.B(n_129),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1606),
.B(n_1686),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1670),
.B(n_130),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1567),
.B(n_132),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1624),
.B(n_132),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1649),
.B(n_1562),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1629),
.B(n_133),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1649),
.B(n_134),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1616),
.B(n_138),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1740),
.B(n_139),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1613),
.B(n_1717),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1678),
.B(n_141),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1547),
.B(n_145),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1576),
.B(n_147),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1738),
.B(n_148),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1599),
.B(n_150),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1714),
.B(n_150),
.Y(n_1964)
);

NAND2xp33_ASAP7_75t_SL g1965 ( 
.A(n_1739),
.B(n_151),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1739),
.B(n_151),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1742),
.B(n_152),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1742),
.B(n_153),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1741),
.B(n_1751),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1751),
.B(n_154),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1698),
.B(n_154),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1698),
.B(n_155),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1678),
.B(n_155),
.Y(n_1973)
);

NAND2xp33_ASAP7_75t_SL g1974 ( 
.A(n_1704),
.B(n_156),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1704),
.B(n_156),
.Y(n_1975)
);

NAND2xp33_ASAP7_75t_SL g1976 ( 
.A(n_1722),
.B(n_157),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_SL g1977 ( 
.A(n_1722),
.B(n_157),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1726),
.B(n_158),
.Y(n_1978)
);

NAND2xp33_ASAP7_75t_SL g1979 ( 
.A(n_1726),
.B(n_158),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1679),
.B(n_159),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1679),
.B(n_1660),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1730),
.B(n_160),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1730),
.B(n_160),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1660),
.B(n_161),
.Y(n_1984)
);

AND3x1_ASAP7_75t_L g1985 ( 
.A(n_1688),
.B(n_162),
.C(n_163),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1662),
.B(n_164),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1748),
.B(n_164),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_SL g1988 ( 
.A(n_1662),
.B(n_165),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_SL g1989 ( 
.A(n_1664),
.B(n_166),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1757),
.B(n_167),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1664),
.B(n_169),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1669),
.B(n_169),
.Y(n_1992)
);

NAND2xp33_ASAP7_75t_SL g1993 ( 
.A(n_1669),
.B(n_170),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1706),
.B(n_171),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_SL g1995 ( 
.A(n_1675),
.B(n_172),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1675),
.B(n_172),
.Y(n_1996)
);

NAND2xp33_ASAP7_75t_SL g1997 ( 
.A(n_1762),
.B(n_173),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1688),
.B(n_1696),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1696),
.B(n_175),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1719),
.B(n_176),
.Y(n_2000)
);

AND2x2_ASAP7_75t_SL g2001 ( 
.A(n_1725),
.B(n_177),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1691),
.B(n_178),
.Y(n_2002)
);

NAND2xp33_ASAP7_75t_SL g2003 ( 
.A(n_1737),
.B(n_178),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1657),
.B(n_179),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1601),
.B(n_180),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1539),
.B(n_180),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1657),
.B(n_181),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1657),
.B(n_181),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1657),
.B(n_183),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1657),
.B(n_184),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1657),
.B(n_184),
.Y(n_2011)
);

NAND2xp33_ASAP7_75t_SL g2012 ( 
.A(n_1539),
.B(n_185),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1657),
.B(n_187),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1539),
.B(n_189),
.Y(n_2014)
);

NAND2xp33_ASAP7_75t_SL g2015 ( 
.A(n_1539),
.B(n_189),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1657),
.B(n_191),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1657),
.B(n_192),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1657),
.B(n_193),
.Y(n_2018)
);

NAND2xp33_ASAP7_75t_SL g2019 ( 
.A(n_1539),
.B(n_194),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1601),
.B(n_197),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1539),
.B(n_198),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1657),
.B(n_199),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1657),
.B(n_201),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1657),
.B(n_201),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1657),
.B(n_202),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1657),
.B(n_202),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1657),
.B(n_203),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1657),
.B(n_204),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1657),
.B(n_205),
.Y(n_2029)
);

NAND2xp33_ASAP7_75t_SL g2030 ( 
.A(n_1539),
.B(n_206),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1657),
.B(n_207),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1657),
.B(n_207),
.Y(n_2032)
);

XNOR2x2_ASAP7_75t_L g2033 ( 
.A(n_1562),
.B(n_208),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1657),
.B(n_209),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1539),
.B(n_209),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1657),
.B(n_210),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1657),
.B(n_211),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_SL g2038 ( 
.A(n_1539),
.B(n_213),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1539),
.B(n_214),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1657),
.B(n_215),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1657),
.B(n_215),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1539),
.B(n_216),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1539),
.B(n_216),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1539),
.B(n_217),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1657),
.B(n_217),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1657),
.B(n_218),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1657),
.B(n_220),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1539),
.B(n_220),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1657),
.B(n_221),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1657),
.B(n_221),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1657),
.B(n_222),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1657),
.B(n_222),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1657),
.B(n_223),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1657),
.B(n_223),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1657),
.B(n_224),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1539),
.B(n_225),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1622),
.B(n_226),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1539),
.B(n_226),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1539),
.B(n_227),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1657),
.B(n_227),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1539),
.B(n_229),
.Y(n_2061)
);

NAND2xp33_ASAP7_75t_SL g2062 ( 
.A(n_1539),
.B(n_230),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1657),
.B(n_230),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1657),
.B(n_231),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_SL g2065 ( 
.A(n_1728),
.B(n_616),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1657),
.B(n_231),
.Y(n_2066)
);

NAND2xp33_ASAP7_75t_SL g2067 ( 
.A(n_1539),
.B(n_232),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1657),
.B(n_232),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1657),
.B(n_233),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_1657),
.B(n_236),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1539),
.B(n_236),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1657),
.B(n_237),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1657),
.B(n_238),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1657),
.B(n_238),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1657),
.B(n_239),
.Y(n_2075)
);

NAND2xp33_ASAP7_75t_SL g2076 ( 
.A(n_1539),
.B(n_241),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1657),
.B(n_241),
.Y(n_2077)
);

NAND2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1539),
.B(n_242),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1539),
.B(n_242),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1657),
.B(n_243),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_1622),
.B(n_244),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1657),
.B(n_244),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1657),
.B(n_245),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1657),
.B(n_245),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1657),
.B(n_247),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1539),
.B(n_247),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1657),
.B(n_248),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1657),
.B(n_249),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1657),
.B(n_249),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1657),
.B(n_250),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1986),
.A2(n_1973),
.B1(n_2081),
.B2(n_2057),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_1769),
.Y(n_2092)
);

AO21x1_ASAP7_75t_L g2093 ( 
.A1(n_1965),
.A2(n_250),
.B(n_251),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_L g2094 ( 
.A(n_1990),
.B(n_252),
.Y(n_2094)
);

OAI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_1813),
.A2(n_253),
.B(n_254),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1910),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1805),
.B(n_254),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_1847),
.A2(n_622),
.B(n_621),
.Y(n_2098)
);

A2O1A1Ixp33_ASAP7_75t_L g2099 ( 
.A1(n_1976),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_2099)
);

AOI221xp5_ASAP7_75t_SL g2100 ( 
.A1(n_1953),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.C(n_259),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1918),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1918),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1850),
.A2(n_627),
.B(n_624),
.Y(n_2103)
);

AOI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_1841),
.A2(n_263),
.B(n_266),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_1766),
.B(n_266),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1805),
.B(n_2043),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1829),
.B(n_268),
.Y(n_2107)
);

NAND2xp33_ASAP7_75t_R g2108 ( 
.A(n_1933),
.B(n_268),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2043),
.B(n_269),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_2057),
.Y(n_2110)
);

OAI22x1_ASAP7_75t_L g2111 ( 
.A1(n_1973),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1829),
.B(n_270),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2048),
.B(n_273),
.Y(n_2113)
);

OAI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2006),
.A2(n_274),
.B(n_275),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2048),
.B(n_277),
.Y(n_2115)
);

AOI21xp33_ASAP7_75t_L g2116 ( 
.A1(n_1958),
.A2(n_278),
.B(n_279),
.Y(n_2116)
);

BUFx4_ASAP7_75t_SL g2117 ( 
.A(n_1771),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1873),
.Y(n_2118)
);

OAI21x1_ASAP7_75t_L g2119 ( 
.A1(n_1836),
.A2(n_630),
.B(n_629),
.Y(n_2119)
);

AO22x2_ASAP7_75t_L g2120 ( 
.A1(n_1973),
.A2(n_283),
.B1(n_280),
.B2(n_282),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1910),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1919),
.Y(n_2122)
);

AOI221x1_ASAP7_75t_L g2123 ( 
.A1(n_2002),
.A2(n_283),
.B1(n_280),
.B2(n_282),
.C(n_284),
.Y(n_2123)
);

OAI21xp33_ASAP7_75t_SL g2124 ( 
.A1(n_1966),
.A2(n_1968),
.B(n_1967),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1856),
.B(n_284),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2058),
.B(n_285),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1849),
.A2(n_637),
.B(n_635),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_2057),
.B(n_286),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_2057),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1795),
.B(n_286),
.Y(n_2130)
);

CKINVDCx11_ASAP7_75t_R g2131 ( 
.A(n_1933),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1795),
.B(n_289),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_2081),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1848),
.Y(n_2134)
);

A2O1A1Ixp33_ASAP7_75t_L g2135 ( 
.A1(n_1977),
.A2(n_293),
.B(n_290),
.C(n_292),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1854),
.B(n_292),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_1832),
.A2(n_640),
.B(n_639),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1834),
.B(n_295),
.Y(n_2138)
);

AOI21xp33_ASAP7_75t_L g2139 ( 
.A1(n_2006),
.A2(n_295),
.B(n_297),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_SL g2140 ( 
.A1(n_1852),
.A2(n_298),
.B(n_299),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_1873),
.Y(n_2141)
);

OAI21x1_ASAP7_75t_L g2142 ( 
.A1(n_1863),
.A2(n_644),
.B(n_643),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1888),
.B(n_299),
.Y(n_2143)
);

OAI21xp33_ASAP7_75t_L g2144 ( 
.A1(n_1981),
.A2(n_300),
.B(n_301),
.Y(n_2144)
);

CKINVDCx8_ASAP7_75t_R g2145 ( 
.A(n_1986),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1919),
.Y(n_2146)
);

A2O1A1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_1979),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_2147)
);

OAI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2014),
.A2(n_302),
.B(n_304),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1925),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1944),
.A2(n_1986),
.B1(n_2081),
.B2(n_1973),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_1974),
.B(n_305),
.C(n_306),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1793),
.B(n_306),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1888),
.B(n_1890),
.Y(n_2153)
);

OAI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2014),
.A2(n_307),
.B(n_308),
.Y(n_2154)
);

A2O1A1Ixp33_ASAP7_75t_L g2155 ( 
.A1(n_1982),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1807),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1925),
.Y(n_2157)
);

AO32x2_ASAP7_75t_L g2158 ( 
.A1(n_2033),
.A2(n_311),
.A3(n_309),
.B1(n_310),
.B2(n_312),
.Y(n_2158)
);

OAI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_2021),
.A2(n_310),
.B(n_312),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1944),
.B(n_313),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_1843),
.B(n_314),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1768),
.B(n_314),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_1774),
.Y(n_2163)
);

BUFx2_ASAP7_75t_L g2164 ( 
.A(n_1933),
.Y(n_2164)
);

NAND3x1_ASAP7_75t_L g2165 ( 
.A(n_1959),
.B(n_319),
.C(n_320),
.Y(n_2165)
);

OAI21xp33_ASAP7_75t_L g2166 ( 
.A1(n_1986),
.A2(n_319),
.B(n_321),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_1840),
.B(n_323),
.Y(n_2167)
);

OAI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2081),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1810),
.B(n_1830),
.Y(n_2169)
);

OAI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_2035),
.A2(n_328),
.B(n_329),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1807),
.Y(n_2171)
);

CKINVDCx11_ASAP7_75t_R g2172 ( 
.A(n_1933),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2035),
.A2(n_331),
.B(n_332),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_SL g2174 ( 
.A1(n_1852),
.A2(n_332),
.B(n_333),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_1941),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2086),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1857),
.B(n_336),
.Y(n_2177)
);

BUFx2_ASAP7_75t_R g2178 ( 
.A(n_1964),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2039),
.A2(n_337),
.B(n_338),
.Y(n_2179)
);

BUFx10_ASAP7_75t_L g2180 ( 
.A(n_1941),
.Y(n_2180)
);

NOR2xp67_ASAP7_75t_L g2181 ( 
.A(n_1941),
.B(n_337),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_2042),
.A2(n_339),
.B(n_340),
.Y(n_2182)
);

OAI21xp5_ASAP7_75t_SL g2183 ( 
.A1(n_1959),
.A2(n_339),
.B(n_340),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2044),
.A2(n_341),
.B(n_342),
.Y(n_2184)
);

OR2x6_ASAP7_75t_L g2185 ( 
.A(n_1941),
.B(n_342),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_1764),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1831),
.B(n_345),
.Y(n_2187)
);

OAI21xp33_ASAP7_75t_L g2188 ( 
.A1(n_1998),
.A2(n_347),
.B(n_348),
.Y(n_2188)
);

AOI21xp33_ASAP7_75t_L g2189 ( 
.A1(n_2056),
.A2(n_349),
.B(n_350),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1943),
.Y(n_2190)
);

AOI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_2059),
.A2(n_350),
.B(n_351),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2061),
.A2(n_351),
.B(n_352),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1812),
.B(n_353),
.Y(n_2193)
);

OR2x6_ASAP7_75t_L g2194 ( 
.A(n_1923),
.B(n_354),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_2071),
.A2(n_355),
.B(n_356),
.Y(n_2195)
);

AOI221xp5_ASAP7_75t_L g2196 ( 
.A1(n_1988),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.C(n_358),
.Y(n_2196)
);

AO21x2_ASAP7_75t_L g2197 ( 
.A1(n_1999),
.A2(n_357),
.B(n_359),
.Y(n_2197)
);

NAND2x1p5_ASAP7_75t_L g2198 ( 
.A(n_1923),
.B(n_359),
.Y(n_2198)
);

NAND2xp33_ASAP7_75t_R g2199 ( 
.A(n_1890),
.B(n_361),
.Y(n_2199)
);

AOI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2079),
.A2(n_362),
.B(n_363),
.Y(n_2200)
);

NOR2x1_ASAP7_75t_SL g2201 ( 
.A(n_1842),
.B(n_1971),
.Y(n_2201)
);

AOI211x1_ASAP7_75t_L g2202 ( 
.A1(n_1987),
.A2(n_367),
.B(n_364),
.C(n_366),
.Y(n_2202)
);

AND3x4_ASAP7_75t_L g2203 ( 
.A(n_1923),
.B(n_368),
.C(n_370),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1989),
.A2(n_373),
.B1(n_370),
.B2(n_372),
.Y(n_2204)
);

INVx3_ASAP7_75t_L g2205 ( 
.A(n_1923),
.Y(n_2205)
);

OAI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_1956),
.A2(n_372),
.B(n_373),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_1993),
.A2(n_381),
.B1(n_376),
.B2(n_377),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1858),
.B(n_383),
.Y(n_2208)
);

AOI21x1_ASAP7_75t_SL g2209 ( 
.A1(n_1860),
.A2(n_385),
.B(n_386),
.Y(n_2209)
);

AND3x1_ASAP7_75t_L g2210 ( 
.A(n_1954),
.B(n_386),
.C(n_387),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_SL g2211 ( 
.A1(n_1972),
.A2(n_389),
.B(n_390),
.Y(n_2211)
);

AOI21xp33_ASAP7_75t_L g2212 ( 
.A1(n_1859),
.A2(n_1855),
.B(n_1962),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1963),
.B(n_391),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_1791),
.B(n_393),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_R g2215 ( 
.A(n_1917),
.B(n_393),
.Y(n_2215)
);

INVxp67_ASAP7_75t_SL g2216 ( 
.A(n_1917),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1833),
.Y(n_2217)
);

A2O1A1Ixp33_ASAP7_75t_L g2218 ( 
.A1(n_1995),
.A2(n_396),
.B(n_394),
.C(n_395),
.Y(n_2218)
);

AOI211x1_ASAP7_75t_L g2219 ( 
.A1(n_1994),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_1927),
.B(n_399),
.Y(n_2220)
);

AOI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_1929),
.A2(n_1948),
.B1(n_1934),
.B2(n_1954),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2001),
.B(n_401),
.Y(n_2222)
);

A2O1A1Ixp33_ASAP7_75t_L g2223 ( 
.A1(n_2012),
.A2(n_403),
.B(n_401),
.C(n_402),
.Y(n_2223)
);

NAND2xp33_ASAP7_75t_R g2224 ( 
.A(n_1929),
.B(n_404),
.Y(n_2224)
);

AND2x6_ASAP7_75t_L g2225 ( 
.A(n_2000),
.B(n_404),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_1934),
.Y(n_2226)
);

A2O1A1Ixp33_ASAP7_75t_L g2227 ( 
.A1(n_2015),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_1833),
.Y(n_2228)
);

AOI221xp5_ASAP7_75t_SL g2229 ( 
.A1(n_1975),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.C(n_414),
.Y(n_2229)
);

AOI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_1942),
.A2(n_410),
.B(n_414),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2001),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1851),
.B(n_416),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_1940),
.A2(n_418),
.B(n_419),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1945),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1969),
.B(n_419),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2000),
.B(n_420),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1827),
.B(n_420),
.Y(n_2237)
);

OAI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_1960),
.A2(n_421),
.B(n_422),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_1814),
.B(n_423),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1816),
.B(n_425),
.Y(n_2240)
);

OAI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_1872),
.A2(n_427),
.B(n_428),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_1823),
.B(n_429),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1868),
.B(n_429),
.Y(n_2243)
);

A2O1A1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_2019),
.A2(n_431),
.B(n_432),
.C(n_433),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_L g2245 ( 
.A(n_1970),
.B(n_432),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1801),
.B(n_434),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_1869),
.B(n_435),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1837),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2005),
.B(n_437),
.Y(n_2249)
);

OR2x2_ASAP7_75t_L g2250 ( 
.A(n_1789),
.B(n_437),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_1777),
.A2(n_438),
.B(n_439),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2020),
.B(n_438),
.Y(n_2252)
);

OAI21x1_ASAP7_75t_L g2253 ( 
.A1(n_1862),
.A2(n_439),
.B(n_440),
.Y(n_2253)
);

OA21x2_ASAP7_75t_L g2254 ( 
.A1(n_1978),
.A2(n_442),
.B(n_443),
.Y(n_2254)
);

AO31x2_ASAP7_75t_L g2255 ( 
.A1(n_1952),
.A2(n_1908),
.A3(n_1980),
.B(n_1900),
.Y(n_2255)
);

OR2x6_ASAP7_75t_L g2256 ( 
.A(n_1991),
.B(n_444),
.Y(n_2256)
);

NAND2x1p5_ASAP7_75t_L g2257 ( 
.A(n_2001),
.B(n_446),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1895),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1779),
.B(n_448),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1864),
.B(n_450),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1825),
.B(n_451),
.Y(n_2261)
);

INVx4_ASAP7_75t_L g2262 ( 
.A(n_1838),
.Y(n_2262)
);

O2A1O1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_1955),
.A2(n_451),
.B(n_452),
.C(n_453),
.Y(n_2263)
);

OAI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_1877),
.A2(n_455),
.B(n_456),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1902),
.Y(n_2265)
);

CKINVDCx6p67_ASAP7_75t_R g2266 ( 
.A(n_1957),
.Y(n_2266)
);

OR2x6_ASAP7_75t_L g2267 ( 
.A(n_1996),
.B(n_457),
.Y(n_2267)
);

INVx2_ASAP7_75t_SL g2268 ( 
.A(n_1775),
.Y(n_2268)
);

OAI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_1883),
.A2(n_457),
.B(n_458),
.Y(n_2269)
);

O2A1O1Ixp5_ASAP7_75t_L g2270 ( 
.A1(n_1874),
.A2(n_459),
.B(n_460),
.C(n_461),
.Y(n_2270)
);

INVxp67_ASAP7_75t_SL g2271 ( 
.A(n_2065),
.Y(n_2271)
);

OAI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_1951),
.A2(n_463),
.B(n_464),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1838),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1907),
.Y(n_2274)
);

AO21x1_ASAP7_75t_L g2275 ( 
.A1(n_1983),
.A2(n_466),
.B(n_467),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1783),
.B(n_468),
.Y(n_2276)
);

BUFx4f_ASAP7_75t_L g2277 ( 
.A(n_1860),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_1767),
.Y(n_2278)
);

OAI21x1_ASAP7_75t_SL g2279 ( 
.A1(n_1984),
.A2(n_468),
.B(n_469),
.Y(n_2279)
);

NOR2xp67_ASAP7_75t_SL g2280 ( 
.A(n_1992),
.B(n_471),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_SL g2281 ( 
.A(n_1916),
.B(n_472),
.C(n_473),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1908),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1815),
.B(n_473),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_1838),
.Y(n_2284)
);

OAI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_1870),
.A2(n_474),
.B(n_475),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1799),
.B(n_476),
.Y(n_2286)
);

INVxp67_ASAP7_75t_SL g2287 ( 
.A(n_2065),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_1817),
.B(n_478),
.Y(n_2288)
);

OR2x2_ASAP7_75t_L g2289 ( 
.A(n_1778),
.B(n_480),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1838),
.Y(n_2290)
);

AO31x2_ASAP7_75t_L g2291 ( 
.A1(n_2033),
.A2(n_1997),
.A3(n_1946),
.B(n_1898),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_SL g2292 ( 
.A1(n_1860),
.A2(n_481),
.B(n_482),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_1824),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1882),
.B(n_483),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1800),
.B(n_484),
.Y(n_2295)
);

CKINVDCx11_ASAP7_75t_R g2296 ( 
.A(n_1985),
.Y(n_2296)
);

OA22x2_ASAP7_75t_L g2297 ( 
.A1(n_1961),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_2297)
);

INVxp67_ASAP7_75t_SL g2298 ( 
.A(n_1880),
.Y(n_2298)
);

AOI21x1_ASAP7_75t_SL g2299 ( 
.A1(n_1861),
.A2(n_490),
.B(n_491),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1826),
.B(n_492),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_1881),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_2301)
);

BUFx2_ASAP7_75t_L g2302 ( 
.A(n_1920),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_1853),
.B(n_1835),
.Y(n_2303)
);

HB1xp67_ASAP7_75t_L g2304 ( 
.A(n_1885),
.Y(n_2304)
);

AND3x4_ASAP7_75t_L g2305 ( 
.A(n_1985),
.B(n_498),
.C(n_499),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_1770),
.Y(n_2306)
);

NAND3xp33_ASAP7_75t_L g2307 ( 
.A(n_2030),
.B(n_500),
.C(n_502),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1950),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1821),
.B(n_502),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1871),
.Y(n_2310)
);

O2A1O1Ixp33_ASAP7_75t_L g2311 ( 
.A1(n_1865),
.A2(n_503),
.B(n_504),
.C(n_505),
.Y(n_2311)
);

O2A1O1Ixp5_ASAP7_75t_L g2312 ( 
.A1(n_1905),
.A2(n_505),
.B(n_506),
.C(n_507),
.Y(n_2312)
);

AO21x2_ASAP7_75t_L g2313 ( 
.A1(n_1909),
.A2(n_506),
.B(n_507),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1811),
.B(n_508),
.Y(n_2314)
);

BUFx6f_ASAP7_75t_L g2315 ( 
.A(n_1772),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_1938),
.B(n_510),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_1887),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_2317)
);

A2O1A1Ixp33_ASAP7_75t_L g2318 ( 
.A1(n_2038),
.A2(n_512),
.B(n_513),
.C(n_514),
.Y(n_2318)
);

AO31x2_ASAP7_75t_L g2319 ( 
.A1(n_1879),
.A2(n_515),
.A3(n_516),
.B(n_517),
.Y(n_2319)
);

A2O1A1Ixp33_ASAP7_75t_L g2320 ( 
.A1(n_2062),
.A2(n_516),
.B(n_519),
.C(n_520),
.Y(n_2320)
);

HB1xp67_ASAP7_75t_L g2321 ( 
.A(n_1886),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_1875),
.A2(n_519),
.B(n_521),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1889),
.Y(n_2323)
);

AOI21xp33_ASAP7_75t_L g2324 ( 
.A1(n_1949),
.A2(n_522),
.B(n_523),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_1876),
.A2(n_525),
.B(n_526),
.Y(n_2325)
);

AO21x2_ASAP7_75t_L g2326 ( 
.A1(n_1897),
.A2(n_525),
.B(n_526),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_1878),
.A2(n_529),
.B(n_530),
.Y(n_2327)
);

A2O1A1Ixp33_ASAP7_75t_L g2328 ( 
.A1(n_2067),
.A2(n_529),
.B(n_530),
.C(n_531),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1891),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1802),
.B(n_533),
.Y(n_2330)
);

OR2x6_ASAP7_75t_L g2331 ( 
.A(n_2004),
.B(n_533),
.Y(n_2331)
);

NAND3xp33_ASAP7_75t_L g2332 ( 
.A(n_2076),
.B(n_2078),
.C(n_1932),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1803),
.B(n_535),
.Y(n_2333)
);

INVx1_ASAP7_75t_SL g2334 ( 
.A(n_1797),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_1930),
.A2(n_535),
.B1(n_536),
.B2(n_537),
.Y(n_2335)
);

INVxp67_ASAP7_75t_L g2336 ( 
.A(n_1792),
.Y(n_2336)
);

AND2x2_ASAP7_75t_SL g2337 ( 
.A(n_1780),
.B(n_614),
.Y(n_2337)
);

BUFx12f_ASAP7_75t_L g2338 ( 
.A(n_2007),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_1781),
.B(n_540),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_1788),
.Y(n_2340)
);

AO32x2_ASAP7_75t_L g2341 ( 
.A1(n_1911),
.A2(n_541),
.A3(n_542),
.B1(n_544),
.B2(n_545),
.Y(n_2341)
);

A2O1A1Ixp33_ASAP7_75t_L g2342 ( 
.A1(n_1912),
.A2(n_1913),
.B(n_1906),
.C(n_2003),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1899),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_1844),
.A2(n_546),
.B(n_550),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_1794),
.B(n_550),
.Y(n_2345)
);

NOR2x1_ASAP7_75t_L g2346 ( 
.A(n_1884),
.B(n_553),
.Y(n_2346)
);

A2O1A1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_1804),
.A2(n_554),
.B(n_555),
.C(n_556),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_1845),
.A2(n_554),
.B(n_556),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2008),
.B(n_557),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_1796),
.B(n_558),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_1892),
.A2(n_559),
.B1(n_560),
.B2(n_561),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_1784),
.B(n_561),
.Y(n_2352)
);

INVxp33_ASAP7_75t_SL g2353 ( 
.A(n_1787),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_1773),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2091),
.A2(n_1819),
.B(n_1820),
.C(n_1893),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2282),
.B(n_1894),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2156),
.B(n_1896),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2171),
.B(n_1921),
.Y(n_2358)
);

NAND3xp33_ASAP7_75t_L g2359 ( 
.A(n_2123),
.B(n_1901),
.C(n_1939),
.Y(n_2359)
);

OAI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2238),
.A2(n_1924),
.B(n_1922),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2145),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2118),
.B(n_2009),
.Y(n_2362)
);

NOR2x1_ASAP7_75t_SL g2363 ( 
.A(n_2185),
.B(n_2194),
.Y(n_2363)
);

O2A1O1Ixp33_ASAP7_75t_L g2364 ( 
.A1(n_2183),
.A2(n_2090),
.B(n_2089),
.C(n_2088),
.Y(n_2364)
);

CKINVDCx20_ASAP7_75t_R g2365 ( 
.A(n_2131),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2271),
.A2(n_1867),
.B(n_1866),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2248),
.Y(n_2367)
);

OAI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_2091),
.A2(n_1926),
.B1(n_1928),
.B2(n_1931),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2160),
.Y(n_2369)
);

INVx2_ASAP7_75t_SL g2370 ( 
.A(n_2117),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2120),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2134),
.Y(n_2372)
);

BUFx5_ASAP7_75t_L g2373 ( 
.A(n_2180),
.Y(n_2373)
);

OAI21x1_ASAP7_75t_L g2374 ( 
.A1(n_2119),
.A2(n_1936),
.B(n_1935),
.Y(n_2374)
);

OAI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_2140),
.A2(n_2087),
.B1(n_2085),
.B2(n_2084),
.Y(n_2375)
);

OAI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2194),
.A2(n_2083),
.B1(n_2082),
.B2(n_2080),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2225),
.A2(n_1903),
.B1(n_1904),
.B2(n_2074),
.Y(n_2377)
);

BUFx2_ASAP7_75t_L g2378 ( 
.A(n_2185),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2172),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_2185),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2194),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_L g2382 ( 
.A1(n_2142),
.A2(n_1914),
.B(n_1915),
.Y(n_2382)
);

OAI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2206),
.A2(n_1937),
.B(n_1947),
.Y(n_2383)
);

NAND2x1p5_ASAP7_75t_L g2384 ( 
.A(n_2128),
.B(n_2164),
.Y(n_2384)
);

INVx1_ASAP7_75t_SL g2385 ( 
.A(n_2175),
.Y(n_2385)
);

NAND2x1p5_ASAP7_75t_L g2386 ( 
.A(n_2128),
.B(n_1765),
.Y(n_2386)
);

NAND2x1p5_ASAP7_75t_L g2387 ( 
.A(n_2110),
.B(n_1846),
.Y(n_2387)
);

OAI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2299),
.A2(n_1828),
.B(n_1818),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_2153),
.B(n_2077),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2141),
.B(n_2010),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2108),
.A2(n_2075),
.B1(n_2073),
.B2(n_2072),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2225),
.A2(n_2070),
.B1(n_2069),
.B2(n_2068),
.Y(n_2392)
);

CKINVDCx16_ASAP7_75t_R g2393 ( 
.A(n_2199),
.Y(n_2393)
);

OAI22x1_ASAP7_75t_L g2394 ( 
.A1(n_2203),
.A2(n_2029),
.B1(n_2064),
.B2(n_2063),
.Y(n_2394)
);

INVx2_ASAP7_75t_SL g2395 ( 
.A(n_2293),
.Y(n_2395)
);

AOI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_2287),
.A2(n_1839),
.B(n_1822),
.Y(n_2396)
);

OAI21x1_ASAP7_75t_L g2397 ( 
.A1(n_2137),
.A2(n_1806),
.B(n_1808),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2337),
.B(n_1776),
.Y(n_2398)
);

NOR3xp33_ASAP7_75t_L g2399 ( 
.A(n_2183),
.B(n_2066),
.C(n_2060),
.Y(n_2399)
);

AOI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2140),
.A2(n_2106),
.B1(n_2210),
.B2(n_2150),
.C(n_2121),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2340),
.Y(n_2401)
);

BUFx12f_ASAP7_75t_L g2402 ( 
.A(n_2180),
.Y(n_2402)
);

INVx5_ASAP7_75t_L g2403 ( 
.A(n_2225),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2105),
.Y(n_2404)
);

OAI21x1_ASAP7_75t_L g2405 ( 
.A1(n_2098),
.A2(n_1809),
.B(n_1782),
.Y(n_2405)
);

BUFx3_ASAP7_75t_L g2406 ( 
.A(n_2353),
.Y(n_2406)
);

AOI22xp33_ASAP7_75t_L g2407 ( 
.A1(n_2225),
.A2(n_2055),
.B1(n_2054),
.B2(n_2053),
.Y(n_2407)
);

OAI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2221),
.A2(n_2052),
.B1(n_2051),
.B2(n_2050),
.Y(n_2408)
);

O2A1O1Ixp33_ASAP7_75t_SL g2409 ( 
.A1(n_2222),
.A2(n_2049),
.B(n_2047),
.C(n_2046),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2143),
.B(n_2045),
.Y(n_2410)
);

OAI22xp5_ASAP7_75t_SL g2411 ( 
.A1(n_2305),
.A2(n_2210),
.B1(n_2257),
.B2(n_2216),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2296),
.A2(n_2041),
.B1(n_2040),
.B2(n_2037),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2096),
.B(n_1786),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2115),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2103),
.A2(n_1785),
.B(n_1798),
.Y(n_2415)
);

AOI221xp5_ASAP7_75t_L g2416 ( 
.A1(n_2122),
.A2(n_2036),
.B1(n_2034),
.B2(n_2032),
.C(n_2031),
.Y(n_2416)
);

BUFx10_ASAP7_75t_L g2417 ( 
.A(n_2239),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_SL g2418 ( 
.A(n_2166),
.B(n_2011),
.Y(n_2418)
);

AO21x2_ASAP7_75t_L g2419 ( 
.A1(n_2279),
.A2(n_2028),
.B(n_2027),
.Y(n_2419)
);

OA21x2_ASAP7_75t_L g2420 ( 
.A1(n_2229),
.A2(n_2026),
.B(n_2025),
.Y(n_2420)
);

AOI22xp33_ASAP7_75t_L g2421 ( 
.A1(n_2256),
.A2(n_2024),
.B1(n_2023),
.B2(n_2022),
.Y(n_2421)
);

OAI21x1_ASAP7_75t_L g2422 ( 
.A1(n_2209),
.A2(n_2018),
.B(n_2017),
.Y(n_2422)
);

OR2x6_ASAP7_75t_L g2423 ( 
.A(n_2198),
.B(n_2016),
.Y(n_2423)
);

OAI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2272),
.A2(n_2013),
.B(n_1790),
.Y(n_2424)
);

OA21x2_ASAP7_75t_L g2425 ( 
.A1(n_2229),
.A2(n_2253),
.B(n_2100),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2226),
.B(n_562),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2236),
.B(n_563),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2107),
.B(n_563),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2092),
.Y(n_2429)
);

CKINVDCx11_ASAP7_75t_R g2430 ( 
.A(n_2338),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2146),
.B(n_2149),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2289),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2112),
.B(n_565),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2157),
.B(n_567),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2129),
.Y(n_2435)
);

INVxp67_ASAP7_75t_SL g2436 ( 
.A(n_2205),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2124),
.A2(n_569),
.B(n_570),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2262),
.B(n_570),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2124),
.A2(n_571),
.B(n_572),
.Y(n_2439)
);

AOI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_2342),
.A2(n_574),
.B(n_575),
.Y(n_2440)
);

INVx2_ASAP7_75t_SL g2441 ( 
.A(n_2310),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2115),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2332),
.A2(n_576),
.B(n_577),
.Y(n_2443)
);

OAI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2332),
.A2(n_580),
.B(n_581),
.Y(n_2444)
);

OAI21x1_ASAP7_75t_L g2445 ( 
.A1(n_2127),
.A2(n_582),
.B(n_583),
.Y(n_2445)
);

AOI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2256),
.A2(n_582),
.B1(n_583),
.B2(n_584),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_2266),
.Y(n_2447)
);

AOI22xp33_ASAP7_75t_L g2448 ( 
.A1(n_2256),
.A2(n_584),
.B1(n_585),
.B2(n_586),
.Y(n_2448)
);

NAND2x1p5_ASAP7_75t_L g2449 ( 
.A(n_2277),
.B(n_587),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2235),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2190),
.B(n_2234),
.Y(n_2451)
);

INVx1_ASAP7_75t_SL g2452 ( 
.A(n_2228),
.Y(n_2452)
);

NAND2x1p5_ASAP7_75t_L g2453 ( 
.A(n_2277),
.B(n_591),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2178),
.B(n_592),
.Y(n_2454)
);

OAI22xp33_ASAP7_75t_L g2455 ( 
.A1(n_2215),
.A2(n_594),
.B1(n_595),
.B2(n_596),
.Y(n_2455)
);

NAND2x1p5_ASAP7_75t_L g2456 ( 
.A(n_2133),
.B(n_2262),
.Y(n_2456)
);

OAI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_2213),
.A2(n_594),
.B(n_595),
.Y(n_2457)
);

AOI22xp33_ASAP7_75t_L g2458 ( 
.A1(n_2267),
.A2(n_597),
.B1(n_599),
.B2(n_600),
.Y(n_2458)
);

INVx6_ASAP7_75t_L g2459 ( 
.A(n_2273),
.Y(n_2459)
);

OAI21x1_ASAP7_75t_SL g2460 ( 
.A1(n_2201),
.A2(n_597),
.B(n_601),
.Y(n_2460)
);

O2A1O1Ixp33_ASAP7_75t_L g2461 ( 
.A1(n_2218),
.A2(n_605),
.B(n_606),
.C(n_607),
.Y(n_2461)
);

OAI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2258),
.A2(n_2274),
.B(n_2265),
.Y(n_2462)
);

INVx1_ASAP7_75t_SL g2463 ( 
.A(n_2302),
.Y(n_2463)
);

NOR2x1_ASAP7_75t_R g2464 ( 
.A(n_2308),
.B(n_609),
.Y(n_2464)
);

AOI22xp33_ASAP7_75t_SL g2465 ( 
.A1(n_2174),
.A2(n_609),
.B1(n_610),
.B2(n_611),
.Y(n_2465)
);

OR2x6_ASAP7_75t_L g2466 ( 
.A(n_2181),
.B(n_612),
.Y(n_2466)
);

OAI221xp5_ASAP7_75t_L g2467 ( 
.A1(n_2224),
.A2(n_2166),
.B1(n_2188),
.B2(n_2204),
.C(n_2144),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2284),
.B(n_2217),
.Y(n_2468)
);

AOI21x1_ASAP7_75t_L g2469 ( 
.A1(n_2280),
.A2(n_2220),
.B(n_2094),
.Y(n_2469)
);

CKINVDCx11_ASAP7_75t_R g2470 ( 
.A(n_2334),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2284),
.B(n_2217),
.Y(n_2471)
);

AOI22xp33_ASAP7_75t_SL g2472 ( 
.A1(n_2214),
.A2(n_2231),
.B1(n_2239),
.B2(n_2151),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2243),
.B(n_2247),
.Y(n_2473)
);

AOI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2267),
.A2(n_2165),
.B1(n_2204),
.B2(n_2168),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2255),
.B(n_2290),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2161),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2331),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2255),
.B(n_2273),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2255),
.B(n_2273),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2260),
.B(n_2294),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2267),
.A2(n_2214),
.B1(n_2281),
.B2(n_2304),
.Y(n_2481)
);

AOI21xp33_ASAP7_75t_L g2482 ( 
.A1(n_2094),
.A2(n_2298),
.B(n_2177),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2331),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2323),
.B(n_2329),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2152),
.B(n_2343),
.Y(n_2485)
);

BUFx2_ASAP7_75t_L g2486 ( 
.A(n_2303),
.Y(n_2486)
);

NAND2x1p5_ASAP7_75t_L g2487 ( 
.A(n_2208),
.B(n_2339),
.Y(n_2487)
);

OA21x2_ASAP7_75t_L g2488 ( 
.A1(n_2114),
.A2(n_2154),
.B(n_2148),
.Y(n_2488)
);

NAND2xp33_ASAP7_75t_R g2489 ( 
.A(n_2254),
.B(n_2250),
.Y(n_2489)
);

INVx4_ASAP7_75t_L g2490 ( 
.A(n_2306),
.Y(n_2490)
);

AO21x2_ASAP7_75t_L g2491 ( 
.A1(n_2093),
.A2(n_2170),
.B(n_2159),
.Y(n_2491)
);

OAI22xp33_ASAP7_75t_L g2492 ( 
.A1(n_2335),
.A2(n_2111),
.B1(n_2297),
.B2(n_2351),
.Y(n_2492)
);

BUFx12f_ASAP7_75t_L g2493 ( 
.A(n_2345),
.Y(n_2493)
);

CKINVDCx16_ASAP7_75t_R g2494 ( 
.A(n_2316),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2303),
.B(n_2245),
.Y(n_2495)
);

NAND2x1p5_ASAP7_75t_L g2496 ( 
.A(n_2125),
.B(n_2245),
.Y(n_2496)
);

BUFx12f_ASAP7_75t_L g2497 ( 
.A(n_2350),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2169),
.B(n_2336),
.Y(n_2498)
);

INVx5_ASAP7_75t_L g2499 ( 
.A(n_2306),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2232),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2167),
.Y(n_2501)
);

OAI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_2173),
.A2(n_2285),
.B(n_2126),
.Y(n_2502)
);

AOI21x1_ASAP7_75t_SL g2503 ( 
.A1(n_2249),
.A2(n_2252),
.B(n_2162),
.Y(n_2503)
);

INVx5_ASAP7_75t_L g2504 ( 
.A(n_2315),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2321),
.B(n_2109),
.Y(n_2505)
);

OAI21x1_ASAP7_75t_L g2506 ( 
.A1(n_2270),
.A2(n_2312),
.B(n_2251),
.Y(n_2506)
);

A2O1A1Ixp33_ASAP7_75t_L g2507 ( 
.A1(n_2307),
.A2(n_2095),
.B(n_2335),
.C(n_2263),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2346),
.B(n_2186),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_SL g2509 ( 
.A(n_2099),
.B(n_2135),
.Y(n_2509)
);

AO31x2_ASAP7_75t_L g2510 ( 
.A1(n_2275),
.A2(n_2155),
.A3(n_2147),
.B(n_2328),
.Y(n_2510)
);

INVx1_ASAP7_75t_SL g2511 ( 
.A(n_2268),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2283),
.B(n_2288),
.Y(n_2512)
);

OA21x2_ASAP7_75t_L g2513 ( 
.A1(n_2241),
.A2(n_2269),
.B(n_2264),
.Y(n_2513)
);

AOI221xp5_ASAP7_75t_L g2514 ( 
.A1(n_2101),
.A2(n_2102),
.B1(n_2187),
.B2(n_2219),
.C(n_2202),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2349),
.B(n_2097),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2319),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2130),
.B(n_2132),
.Y(n_2517)
);

OA21x2_ASAP7_75t_L g2518 ( 
.A1(n_2184),
.A2(n_2212),
.B(n_2227),
.Y(n_2518)
);

AO32x2_ASAP7_75t_L g2519 ( 
.A1(n_2176),
.A2(n_2317),
.A3(n_2301),
.B1(n_2354),
.B2(n_2278),
.Y(n_2519)
);

OAI21x1_ASAP7_75t_L g2520 ( 
.A1(n_2179),
.A2(n_2200),
.B(n_2195),
.Y(n_2520)
);

OAI21x1_ASAP7_75t_SL g2521 ( 
.A1(n_2207),
.A2(n_2196),
.B(n_2351),
.Y(n_2521)
);

OAI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2182),
.A2(n_2192),
.B(n_2191),
.Y(n_2522)
);

AO21x2_ASAP7_75t_L g2523 ( 
.A1(n_2197),
.A2(n_2104),
.B(n_2313),
.Y(n_2523)
);

OR2x6_ASAP7_75t_L g2524 ( 
.A(n_2292),
.B(n_2211),
.Y(n_2524)
);

O2A1O1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2223),
.A2(n_2320),
.B(n_2318),
.C(n_2244),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2315),
.Y(n_2526)
);

OAI21xp33_ASAP7_75t_L g2527 ( 
.A1(n_2113),
.A2(n_2347),
.B(n_2116),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2291),
.B(n_2136),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2319),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2138),
.Y(n_2530)
);

OAI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2202),
.A2(n_2219),
.B1(n_2242),
.B2(n_2240),
.Y(n_2531)
);

OAI21x1_ASAP7_75t_L g2532 ( 
.A1(n_2344),
.A2(n_2348),
.B(n_2322),
.Y(n_2532)
);

AO21x2_ASAP7_75t_L g2533 ( 
.A1(n_2197),
.A2(n_2313),
.B(n_2326),
.Y(n_2533)
);

OAI21x1_ASAP7_75t_L g2534 ( 
.A1(n_2325),
.A2(n_2327),
.B(n_2233),
.Y(n_2534)
);

OAI21x1_ASAP7_75t_L g2535 ( 
.A1(n_2230),
.A2(n_2237),
.B(n_2311),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2314),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2193),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2163),
.B(n_2291),
.Y(n_2538)
);

INVxp67_ASAP7_75t_SL g2539 ( 
.A(n_2352),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2246),
.Y(n_2540)
);

INVx1_ASAP7_75t_SL g2541 ( 
.A(n_2261),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_2291),
.Y(n_2542)
);

OAI21x1_ASAP7_75t_L g2543 ( 
.A1(n_2309),
.A2(n_2295),
.B(n_2286),
.Y(n_2543)
);

OA21x2_ASAP7_75t_L g2544 ( 
.A1(n_2139),
.A2(n_2189),
.B(n_2259),
.Y(n_2544)
);

OR3x4_ASAP7_75t_SL g2545 ( 
.A(n_2158),
.B(n_2341),
.C(n_2324),
.Y(n_2545)
);

OR2x2_ASAP7_75t_L g2546 ( 
.A(n_2276),
.B(n_2333),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2158),
.B(n_2330),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2367),
.Y(n_2548)
);

INVxp33_ASAP7_75t_L g2549 ( 
.A(n_2363),
.Y(n_2549)
);

BUFx3_ASAP7_75t_L g2550 ( 
.A(n_2402),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2375),
.B(n_2408),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2432),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2372),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_2370),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2434),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2431),
.B(n_2300),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2427),
.B(n_2341),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2428),
.B(n_2433),
.Y(n_2558)
);

OAI21xp5_ASAP7_75t_L g2559 ( 
.A1(n_2507),
.A2(n_2525),
.B(n_2359),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2451),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2451),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2473),
.B(n_2512),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2438),
.Y(n_2563)
);

AND2x4_ASAP7_75t_L g2564 ( 
.A(n_2403),
.B(n_2495),
.Y(n_2564)
);

INVxp67_ASAP7_75t_SL g2565 ( 
.A(n_2478),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2369),
.B(n_2371),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2403),
.Y(n_2567)
);

INVx8_ASAP7_75t_L g2568 ( 
.A(n_2365),
.Y(n_2568)
);

INVxp67_ASAP7_75t_L g2569 ( 
.A(n_2381),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2484),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2438),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_2495),
.B(n_2468),
.Y(n_2572)
);

INVx4_ASAP7_75t_SL g2573 ( 
.A(n_2466),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2501),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2450),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_SL g2576 ( 
.A1(n_2467),
.A2(n_2378),
.B1(n_2411),
.B2(n_2393),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2480),
.B(n_2515),
.Y(n_2577)
);

OAI21xp33_ASAP7_75t_SL g2578 ( 
.A1(n_2400),
.A2(n_2474),
.B(n_2439),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2494),
.B(n_2426),
.Y(n_2579)
);

BUFx4f_ASAP7_75t_L g2580 ( 
.A(n_2449),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2414),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2442),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2404),
.B(n_2410),
.Y(n_2583)
);

CKINVDCx20_ASAP7_75t_R g2584 ( 
.A(n_2430),
.Y(n_2584)
);

NOR2xp67_ASAP7_75t_SL g2585 ( 
.A(n_2477),
.B(n_2483),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2408),
.B(n_2389),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2478),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_2468),
.B(n_2471),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2413),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2498),
.B(n_2476),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2362),
.B(n_2390),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2511),
.B(n_2441),
.Y(n_2592)
);

OR2x2_ASAP7_75t_L g2593 ( 
.A(n_2401),
.B(n_2429),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2516),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2380),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2358),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2529),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2452),
.Y(n_2598)
);

HB1xp67_ASAP7_75t_SL g2599 ( 
.A(n_2373),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2537),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2479),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2462),
.B(n_2547),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2511),
.B(n_2417),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2406),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2417),
.B(n_2536),
.Y(n_2605)
);

OR2x6_ASAP7_75t_L g2606 ( 
.A(n_2384),
.B(n_2466),
.Y(n_2606)
);

INVx4_ASAP7_75t_L g2607 ( 
.A(n_2466),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2479),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2357),
.Y(n_2609)
);

INVx4_ASAP7_75t_L g2610 ( 
.A(n_2449),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_2411),
.B(n_2376),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2357),
.Y(n_2612)
);

INVx2_ASAP7_75t_SL g2613 ( 
.A(n_2447),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2462),
.B(n_2528),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2505),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2505),
.Y(n_2616)
);

BUFx2_ASAP7_75t_L g2617 ( 
.A(n_2373),
.Y(n_2617)
);

BUFx2_ASAP7_75t_L g2618 ( 
.A(n_2373),
.Y(n_2618)
);

HB1xp67_ASAP7_75t_L g2619 ( 
.A(n_2475),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2475),
.Y(n_2620)
);

OAI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2525),
.A2(n_2359),
.B(n_2461),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2540),
.B(n_2500),
.Y(n_2622)
);

INVx1_ASAP7_75t_SL g2623 ( 
.A(n_2452),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2530),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2400),
.B(n_2531),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2356),
.Y(n_2626)
);

INVx3_ASAP7_75t_L g2627 ( 
.A(n_2373),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2356),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2385),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2485),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2384),
.B(n_2486),
.Y(n_2631)
);

OAI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2474),
.A2(n_2467),
.B1(n_2472),
.B2(n_2481),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2395),
.B(n_2463),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2531),
.B(n_2538),
.Y(n_2634)
);

HB1xp67_ASAP7_75t_L g2635 ( 
.A(n_2385),
.Y(n_2635)
);

OAI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2437),
.A2(n_2439),
.B1(n_2492),
.B2(n_2458),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2373),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2399),
.B(n_2541),
.Y(n_2638)
);

HB1xp67_ASAP7_75t_L g2639 ( 
.A(n_2538),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_2526),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2456),
.Y(n_2641)
);

OR2x6_ASAP7_75t_L g2642 ( 
.A(n_2437),
.B(n_2453),
.Y(n_2642)
);

A2O1A1Ixp33_ASAP7_75t_L g2643 ( 
.A1(n_2443),
.A2(n_2444),
.B(n_2355),
.C(n_2440),
.Y(n_2643)
);

AOI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2376),
.A2(n_2455),
.B1(n_2391),
.B2(n_2418),
.Y(n_2644)
);

INVx4_ASAP7_75t_L g2645 ( 
.A(n_2499),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2541),
.B(n_2470),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2386),
.Y(n_2647)
);

INVxp33_ASAP7_75t_L g2648 ( 
.A(n_2464),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2508),
.Y(n_2649)
);

INVx3_ASAP7_75t_L g2650 ( 
.A(n_2456),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2508),
.Y(n_2651)
);

INVx4_ASAP7_75t_L g2652 ( 
.A(n_2499),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2420),
.Y(n_2653)
);

AO21x2_ASAP7_75t_L g2654 ( 
.A1(n_2482),
.A2(n_2533),
.B(n_2523),
.Y(n_2654)
);

AND2x4_ASAP7_75t_L g2655 ( 
.A(n_2471),
.B(n_2361),
.Y(n_2655)
);

OAI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2440),
.A2(n_2444),
.B(n_2443),
.Y(n_2656)
);

INVx4_ASAP7_75t_SL g2657 ( 
.A(n_2524),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2542),
.Y(n_2658)
);

HB1xp67_ASAP7_75t_L g2659 ( 
.A(n_2489),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_SL g2660 ( 
.A(n_2418),
.B(n_2524),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2460),
.Y(n_2661)
);

OAI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2502),
.A2(n_2514),
.B(n_2457),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2539),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2457),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2361),
.Y(n_2665)
);

AO21x2_ASAP7_75t_L g2666 ( 
.A1(n_2523),
.A2(n_2366),
.B(n_2521),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2499),
.Y(n_2667)
);

OAI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2509),
.A2(n_2423),
.B1(n_2391),
.B2(n_2524),
.Y(n_2668)
);

AND2x4_ASAP7_75t_L g2669 ( 
.A(n_2435),
.B(n_2436),
.Y(n_2669)
);

HB1xp67_ASAP7_75t_L g2670 ( 
.A(n_2425),
.Y(n_2670)
);

AND2x4_ASAP7_75t_L g2671 ( 
.A(n_2435),
.B(n_2504),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2491),
.B(n_2488),
.Y(n_2672)
);

INVx4_ASAP7_75t_L g2673 ( 
.A(n_2504),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2493),
.B(n_2497),
.Y(n_2674)
);

HB1xp67_ASAP7_75t_L g2675 ( 
.A(n_2425),
.Y(n_2675)
);

BUFx2_ASAP7_75t_L g2676 ( 
.A(n_2490),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2504),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2446),
.B(n_2448),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2490),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2459),
.Y(n_2680)
);

OR2x6_ASAP7_75t_L g2681 ( 
.A(n_2423),
.B(n_2496),
.Y(n_2681)
);

OR2x6_ASAP7_75t_L g2682 ( 
.A(n_2606),
.B(n_2423),
.Y(n_2682)
);

NAND2xp33_ASAP7_75t_R g2683 ( 
.A(n_2606),
.B(n_2379),
.Y(n_2683)
);

CKINVDCx20_ASAP7_75t_R g2684 ( 
.A(n_2584),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_2558),
.Y(n_2685)
);

NAND2xp33_ASAP7_75t_R g2686 ( 
.A(n_2606),
.B(n_2454),
.Y(n_2686)
);

BUFx10_ASAP7_75t_L g2687 ( 
.A(n_2554),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2552),
.Y(n_2688)
);

NAND2xp33_ASAP7_75t_R g2689 ( 
.A(n_2611),
.B(n_2464),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_R g2690 ( 
.A(n_2584),
.B(n_2469),
.Y(n_2690)
);

NAND2xp33_ASAP7_75t_R g2691 ( 
.A(n_2611),
.B(n_2513),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2615),
.B(n_2517),
.Y(n_2692)
);

NAND2xp33_ASAP7_75t_R g2693 ( 
.A(n_2676),
.B(n_2518),
.Y(n_2693)
);

CKINVDCx8_ASAP7_75t_R g2694 ( 
.A(n_2568),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2616),
.B(n_2514),
.Y(n_2695)
);

NAND2xp33_ASAP7_75t_R g2696 ( 
.A(n_2617),
.B(n_2518),
.Y(n_2696)
);

AND2x4_ASAP7_75t_L g2697 ( 
.A(n_2573),
.B(n_2419),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2574),
.B(n_2546),
.Y(n_2698)
);

INVxp67_ASAP7_75t_L g2699 ( 
.A(n_2593),
.Y(n_2699)
);

AND2x4_ASAP7_75t_L g2700 ( 
.A(n_2573),
.B(n_2419),
.Y(n_2700)
);

OR2x6_ASAP7_75t_L g2701 ( 
.A(n_2607),
.B(n_2398),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2575),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_R g2703 ( 
.A(n_2599),
.B(n_2550),
.Y(n_2703)
);

BUFx2_ASAP7_75t_R g2704 ( 
.A(n_2550),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2577),
.B(n_2562),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_L g2706 ( 
.A(n_2648),
.B(n_2364),
.Y(n_2706)
);

BUFx3_ASAP7_75t_L g2707 ( 
.A(n_2568),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_R g2708 ( 
.A(n_2568),
.B(n_2580),
.Y(n_2708)
);

AND2x4_ASAP7_75t_L g2709 ( 
.A(n_2573),
.B(n_2396),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_R g2710 ( 
.A(n_2580),
.B(n_2607),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2583),
.B(n_2633),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_R g2712 ( 
.A(n_2613),
.B(n_2421),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2600),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2638),
.B(n_2543),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2592),
.B(n_2544),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_R g2716 ( 
.A(n_2660),
.B(n_2412),
.Y(n_2716)
);

NAND2xp33_ASAP7_75t_R g2717 ( 
.A(n_2618),
.B(n_2544),
.Y(n_2717)
);

INVxp67_ASAP7_75t_L g2718 ( 
.A(n_2590),
.Y(n_2718)
);

NAND2xp33_ASAP7_75t_R g2719 ( 
.A(n_2642),
.B(n_2677),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2560),
.B(n_2394),
.Y(n_2720)
);

NAND2xp33_ASAP7_75t_R g2721 ( 
.A(n_2642),
.B(n_2424),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2624),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2622),
.Y(n_2723)
);

OR2x4_ASAP7_75t_L g2724 ( 
.A(n_2551),
.B(n_2545),
.Y(n_2724)
);

NAND2xp33_ASAP7_75t_R g2725 ( 
.A(n_2642),
.B(n_2424),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_R g2726 ( 
.A(n_2660),
.B(n_2392),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2561),
.B(n_2630),
.Y(n_2727)
);

XNOR2xp5_ASAP7_75t_L g2728 ( 
.A(n_2648),
.B(n_2407),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2566),
.Y(n_2729)
);

NAND2xp33_ASAP7_75t_R g2730 ( 
.A(n_2677),
.B(n_2422),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2604),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2591),
.B(n_2519),
.Y(n_2732)
);

BUFx3_ASAP7_75t_L g2733 ( 
.A(n_2667),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2674),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_R g2735 ( 
.A(n_2627),
.B(n_2637),
.Y(n_2735)
);

NAND2xp33_ASAP7_75t_R g2736 ( 
.A(n_2567),
.B(n_2646),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_R g2737 ( 
.A(n_2627),
.B(n_2509),
.Y(n_2737)
);

CKINVDCx16_ASAP7_75t_R g2738 ( 
.A(n_2579),
.Y(n_2738)
);

XNOR2xp5_ASAP7_75t_L g2739 ( 
.A(n_2576),
.B(n_2416),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2586),
.B(n_2589),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2657),
.B(n_2388),
.Y(n_2741)
);

INVxp67_ASAP7_75t_L g2742 ( 
.A(n_2598),
.Y(n_2742)
);

XNOR2xp5_ASAP7_75t_L g2743 ( 
.A(n_2576),
.B(n_2416),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2595),
.B(n_2519),
.Y(n_2744)
);

AND2x4_ASAP7_75t_L g2745 ( 
.A(n_2639),
.B(n_2520),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_R g2746 ( 
.A(n_2637),
.B(n_2610),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2581),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2586),
.B(n_2465),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2598),
.B(n_2496),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_R g2750 ( 
.A(n_2610),
.B(n_2377),
.Y(n_2750)
);

AND2x4_ASAP7_75t_L g2751 ( 
.A(n_2639),
.B(n_2522),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2667),
.Y(n_2752)
);

NAND2xp33_ASAP7_75t_R g2753 ( 
.A(n_2679),
.B(n_2383),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2582),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2681),
.B(n_2534),
.Y(n_2755)
);

NAND2xp33_ASAP7_75t_R g2756 ( 
.A(n_2679),
.B(n_2360),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_R g2757 ( 
.A(n_2641),
.B(n_2409),
.Y(n_2757)
);

CKINVDCx20_ASAP7_75t_R g2758 ( 
.A(n_2603),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_R g2759 ( 
.A(n_2641),
.B(n_2503),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2548),
.B(n_2368),
.Y(n_2760)
);

BUFx24_ASAP7_75t_SL g2761 ( 
.A(n_2644),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_R g2762 ( 
.A(n_2650),
.B(n_2487),
.Y(n_2762)
);

OR2x4_ASAP7_75t_L g2763 ( 
.A(n_2551),
.B(n_2527),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2564),
.B(n_2532),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2629),
.Y(n_2765)
);

NAND2xp33_ASAP7_75t_R g2766 ( 
.A(n_2650),
.B(n_2360),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2553),
.B(n_2527),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2564),
.B(n_2535),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2555),
.B(n_2510),
.Y(n_2769)
);

XNOR2xp5_ASAP7_75t_L g2770 ( 
.A(n_2632),
.B(n_2487),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_SL g2771 ( 
.A(n_2585),
.B(n_2387),
.Y(n_2771)
);

BUFx2_ASAP7_75t_L g2772 ( 
.A(n_2623),
.Y(n_2772)
);

INVxp67_ASAP7_75t_L g2773 ( 
.A(n_2629),
.Y(n_2773)
);

XNOR2xp5_ASAP7_75t_L g2774 ( 
.A(n_2632),
.B(n_2415),
.Y(n_2774)
);

INVxp67_ASAP7_75t_L g2775 ( 
.A(n_2635),
.Y(n_2775)
);

AND2x4_ASAP7_75t_L g2776 ( 
.A(n_2649),
.B(n_2510),
.Y(n_2776)
);

NAND2xp33_ASAP7_75t_R g2777 ( 
.A(n_2625),
.B(n_2445),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2651),
.B(n_2405),
.Y(n_2778)
);

NAND2xp33_ASAP7_75t_R g2779 ( 
.A(n_2625),
.B(n_2397),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2570),
.B(n_2374),
.Y(n_2780)
);

XNOR2xp5_ASAP7_75t_L g2781 ( 
.A(n_2668),
.B(n_2506),
.Y(n_2781)
);

BUFx10_ASAP7_75t_L g2782 ( 
.A(n_2671),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2569),
.B(n_2382),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2587),
.B(n_2601),
.Y(n_2784)
);

XNOR2xp5_ASAP7_75t_L g2785 ( 
.A(n_2668),
.B(n_2549),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2626),
.B(n_2628),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_R g2787 ( 
.A(n_2645),
.B(n_2652),
.Y(n_2787)
);

AND2x2_ASAP7_75t_L g2788 ( 
.A(n_2569),
.B(n_2640),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2609),
.B(n_2612),
.Y(n_2789)
);

NAND2xp33_ASAP7_75t_R g2790 ( 
.A(n_2605),
.B(n_2557),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_R g2791 ( 
.A(n_2645),
.B(n_2652),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_R g2792 ( 
.A(n_2673),
.B(n_2631),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2640),
.B(n_2588),
.Y(n_2793)
);

NAND2xp33_ASAP7_75t_R g2794 ( 
.A(n_2655),
.B(n_2669),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2596),
.Y(n_2795)
);

XNOR2xp5_ASAP7_75t_L g2796 ( 
.A(n_2549),
.B(n_2636),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2673),
.Y(n_2797)
);

XNOR2xp5_ASAP7_75t_L g2798 ( 
.A(n_2636),
.B(n_2588),
.Y(n_2798)
);

BUFx3_ASAP7_75t_L g2799 ( 
.A(n_2655),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2556),
.B(n_2602),
.Y(n_2800)
);

NAND2xp33_ASAP7_75t_R g2801 ( 
.A(n_2669),
.B(n_2563),
.Y(n_2801)
);

BUFx3_ASAP7_75t_L g2802 ( 
.A(n_2680),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2587),
.B(n_2601),
.Y(n_2803)
);

INVxp67_ASAP7_75t_L g2804 ( 
.A(n_2635),
.Y(n_2804)
);

INVxp67_ASAP7_75t_L g2805 ( 
.A(n_2665),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2608),
.B(n_2572),
.Y(n_2806)
);

AND2x4_ASAP7_75t_L g2807 ( 
.A(n_2608),
.B(n_2572),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_R g2808 ( 
.A(n_2659),
.B(n_2647),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2715),
.B(n_2619),
.Y(n_2809)
);

OR2x2_ASAP7_75t_L g2810 ( 
.A(n_2765),
.B(n_2619),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2708),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_SL g2812 ( 
.A(n_2703),
.B(n_2578),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2714),
.B(n_2634),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2702),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2713),
.Y(n_2815)
);

NOR2x1_ASAP7_75t_L g2816 ( 
.A(n_2733),
.B(n_2559),
.Y(n_2816)
);

CKINVDCx5p33_ASAP7_75t_R g2817 ( 
.A(n_2683),
.Y(n_2817)
);

OR2x2_ASAP7_75t_L g2818 ( 
.A(n_2773),
.B(n_2620),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2795),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2732),
.B(n_2664),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2776),
.B(n_2744),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2776),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2800),
.B(n_2634),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2745),
.B(n_2565),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2745),
.B(n_2565),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2722),
.Y(n_2826)
);

INVx2_ASAP7_75t_SL g2827 ( 
.A(n_2792),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2784),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2751),
.B(n_2666),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2697),
.B(n_2659),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2688),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2723),
.B(n_2662),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2751),
.B(n_2666),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2780),
.Y(n_2834)
);

NAND3xp33_ASAP7_75t_L g2835 ( 
.A(n_2691),
.B(n_2706),
.C(n_2739),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2783),
.B(n_2620),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2740),
.B(n_2662),
.Y(n_2837)
);

INVxp33_ASAP7_75t_L g2838 ( 
.A(n_2808),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2769),
.B(n_2653),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2747),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2789),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2743),
.A2(n_2678),
.B1(n_2656),
.B2(n_2661),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2803),
.B(n_2658),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2803),
.B(n_2658),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2729),
.B(n_2654),
.Y(n_2845)
);

AOI22xp33_ASAP7_75t_L g2846 ( 
.A1(n_2796),
.A2(n_2656),
.B1(n_2559),
.B2(n_2621),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2778),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2786),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2806),
.B(n_2654),
.Y(n_2849)
);

BUFx2_ASAP7_75t_L g2850 ( 
.A(n_2735),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2806),
.B(n_2594),
.Y(n_2851)
);

INVx1_ASAP7_75t_SL g2852 ( 
.A(n_2704),
.Y(n_2852)
);

OR2x2_ASAP7_75t_L g2853 ( 
.A(n_2775),
.B(n_2614),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_2804),
.B(n_2614),
.Y(n_2854)
);

NAND2x1p5_ASAP7_75t_L g2855 ( 
.A(n_2741),
.B(n_2571),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2727),
.Y(n_2856)
);

NOR2x1_ASAP7_75t_L g2857 ( 
.A(n_2707),
.B(n_2682),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2807),
.B(n_2597),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2807),
.B(n_2670),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2705),
.B(n_2663),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2767),
.Y(n_2861)
);

INVx2_ASAP7_75t_SL g2862 ( 
.A(n_2782),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2754),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2711),
.B(n_2670),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2768),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2698),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2760),
.Y(n_2867)
);

NAND3xp33_ASAP7_75t_SL g2868 ( 
.A(n_2694),
.B(n_2643),
.C(n_2621),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2834),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2829),
.B(n_2697),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2823),
.B(n_2788),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_SL g2872 ( 
.A(n_2827),
.B(n_2746),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2813),
.B(n_2700),
.Y(n_2873)
);

INVx3_ASAP7_75t_L g2874 ( 
.A(n_2830),
.Y(n_2874)
);

OAI221xp5_ASAP7_75t_L g2875 ( 
.A1(n_2842),
.A2(n_2846),
.B1(n_2835),
.B2(n_2689),
.C(n_2812),
.Y(n_2875)
);

OR2x2_ASAP7_75t_L g2876 ( 
.A(n_2809),
.B(n_2699),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_R g2877 ( 
.A(n_2811),
.B(n_2736),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2827),
.Y(n_2878)
);

BUFx3_ASAP7_75t_L g2879 ( 
.A(n_2811),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2813),
.B(n_2700),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2823),
.B(n_2720),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2826),
.Y(n_2882)
);

NAND2xp33_ASAP7_75t_SL g2883 ( 
.A(n_2838),
.B(n_2737),
.Y(n_2883)
);

HB1xp67_ASAP7_75t_L g2884 ( 
.A(n_2828),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2826),
.Y(n_2885)
);

INVx3_ASAP7_75t_L g2886 ( 
.A(n_2830),
.Y(n_2886)
);

BUFx3_ASAP7_75t_L g2887 ( 
.A(n_2862),
.Y(n_2887)
);

BUFx6f_ASAP7_75t_L g2888 ( 
.A(n_2830),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2850),
.Y(n_2889)
);

INVx4_ASAP7_75t_L g2890 ( 
.A(n_2850),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2821),
.B(n_2793),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2821),
.B(n_2675),
.Y(n_2892)
);

AOI221xp5_ASAP7_75t_SL g2893 ( 
.A1(n_2852),
.A2(n_2798),
.B1(n_2685),
.B2(n_2770),
.C(n_2718),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2868),
.A2(n_2774),
.B1(n_2716),
.B2(n_2785),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2864),
.B(n_2675),
.Y(n_2895)
);

BUFx2_ASAP7_75t_L g2896 ( 
.A(n_2857),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2864),
.B(n_2772),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2809),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2849),
.B(n_2749),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2853),
.B(n_2742),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2853),
.B(n_2672),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2816),
.Y(n_2902)
);

OR2x2_ASAP7_75t_L g2903 ( 
.A(n_2854),
.B(n_2672),
.Y(n_2903)
);

INVxp67_ASAP7_75t_L g2904 ( 
.A(n_2862),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2855),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2831),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2849),
.B(n_2764),
.Y(n_2907)
);

HB1xp67_ASAP7_75t_L g2908 ( 
.A(n_2810),
.Y(n_2908)
);

INVx1_ASAP7_75t_SL g2909 ( 
.A(n_2817),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2824),
.B(n_2764),
.Y(n_2910)
);

OAI221xp5_ASAP7_75t_L g2911 ( 
.A1(n_2837),
.A2(n_2728),
.B1(n_2686),
.B2(n_2725),
.C(n_2721),
.Y(n_2911)
);

INVx1_ASAP7_75t_SL g2912 ( 
.A(n_2817),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2819),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2899),
.B(n_2833),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2898),
.B(n_2854),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2908),
.B(n_2867),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2899),
.B(n_2833),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2907),
.B(n_2824),
.Y(n_2918)
);

INVxp67_ASAP7_75t_L g2919 ( 
.A(n_2889),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2901),
.B(n_2867),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_2890),
.B(n_2865),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2900),
.Y(n_2922)
);

OR2x2_ASAP7_75t_L g2923 ( 
.A(n_2900),
.B(n_2860),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2901),
.B(n_2820),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2907),
.B(n_2825),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2891),
.B(n_2825),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2891),
.B(n_2836),
.Y(n_2927)
);

OR2x2_ASAP7_75t_L g2928 ( 
.A(n_2903),
.B(n_2810),
.Y(n_2928)
);

AOI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2875),
.A2(n_2763),
.B1(n_2790),
.B2(n_2724),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2903),
.B(n_2861),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2882),
.Y(n_2931)
);

HB1xp67_ASAP7_75t_L g2932 ( 
.A(n_2884),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2897),
.B(n_2836),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2897),
.B(n_2859),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2882),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2881),
.B(n_2861),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2885),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2895),
.B(n_2845),
.Y(n_2938)
);

OR2x2_ASAP7_75t_L g2939 ( 
.A(n_2876),
.B(n_2818),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2892),
.B(n_2859),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2892),
.B(n_2843),
.Y(n_2941)
);

INVx2_ASAP7_75t_SL g2942 ( 
.A(n_2890),
.Y(n_2942)
);

HB1xp67_ASAP7_75t_L g2943 ( 
.A(n_2890),
.Y(n_2943)
);

INVxp67_ASAP7_75t_L g2944 ( 
.A(n_2889),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2887),
.Y(n_2945)
);

AND2x4_ASAP7_75t_L g2946 ( 
.A(n_2870),
.B(n_2865),
.Y(n_2946)
);

INVx2_ASAP7_75t_SL g2947 ( 
.A(n_2887),
.Y(n_2947)
);

NAND2xp67_ASAP7_75t_L g2948 ( 
.A(n_2877),
.B(n_2845),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2895),
.B(n_2843),
.Y(n_2949)
);

INVx1_ASAP7_75t_SL g2950 ( 
.A(n_2879),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2873),
.B(n_2844),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2869),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2873),
.B(n_2844),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2879),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2880),
.B(n_2822),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2885),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2880),
.B(n_2822),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2910),
.B(n_2851),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2870),
.B(n_2847),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2871),
.B(n_2839),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2910),
.B(n_2851),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2870),
.B(n_2858),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2914),
.B(n_2896),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2950),
.B(n_2909),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2932),
.B(n_2902),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2922),
.B(n_2841),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_2954),
.Y(n_2967)
);

OAI221xp5_ASAP7_75t_L g2968 ( 
.A1(n_2929),
.A2(n_2893),
.B1(n_2911),
.B2(n_2894),
.C(n_2896),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2915),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2927),
.B(n_2841),
.Y(n_2970)
);

OAI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2942),
.A2(n_2878),
.B1(n_2794),
.B2(n_2874),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_SL g2972 ( 
.A(n_2942),
.B(n_2893),
.Y(n_2972)
);

OAI221xp5_ASAP7_75t_L g2973 ( 
.A1(n_2943),
.A2(n_2883),
.B1(n_2878),
.B2(n_2872),
.C(n_2904),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_R g2974 ( 
.A(n_2954),
.B(n_2684),
.Y(n_2974)
);

CKINVDCx14_ASAP7_75t_R g2975 ( 
.A(n_2923),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2927),
.B(n_2848),
.Y(n_2976)
);

INVxp33_ASAP7_75t_SL g2977 ( 
.A(n_2962),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2920),
.B(n_2916),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2924),
.B(n_2848),
.Y(n_2979)
);

OR2x2_ASAP7_75t_L g2980 ( 
.A(n_2928),
.B(n_2876),
.Y(n_2980)
);

AO221x2_ASAP7_75t_L g2981 ( 
.A1(n_2948),
.A2(n_2738),
.B1(n_2710),
.B2(n_2866),
.C(n_2719),
.Y(n_2981)
);

AOI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2945),
.A2(n_2870),
.B1(n_2912),
.B2(n_2693),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2915),
.B(n_2856),
.Y(n_2983)
);

AO221x2_ASAP7_75t_L g2984 ( 
.A1(n_2948),
.A2(n_2731),
.B1(n_2801),
.B2(n_2687),
.C(n_2758),
.Y(n_2984)
);

NOR2x1_ASAP7_75t_L g2985 ( 
.A(n_2921),
.B(n_2682),
.Y(n_2985)
);

NAND2xp33_ASAP7_75t_SL g2986 ( 
.A(n_2945),
.B(n_2787),
.Y(n_2986)
);

AND2x4_ASAP7_75t_L g2987 ( 
.A(n_2947),
.B(n_2874),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2933),
.B(n_2856),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_2947),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2933),
.B(n_2906),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2919),
.B(n_2734),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2936),
.B(n_2913),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2939),
.B(n_2928),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2939),
.B(n_2913),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2963),
.B(n_2914),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2972),
.B(n_2975),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2994),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2993),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2969),
.B(n_2960),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2978),
.B(n_2926),
.Y(n_3000)
);

AOI22xp33_ASAP7_75t_L g3001 ( 
.A1(n_2968),
.A2(n_2726),
.B1(n_2781),
.B2(n_2946),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2980),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2970),
.B(n_2926),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2983),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2976),
.B(n_2917),
.Y(n_3005)
);

AND2x2_ASAP7_75t_L g3006 ( 
.A(n_2987),
.B(n_2917),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2987),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2982),
.B(n_2940),
.Y(n_3008)
);

INVx1_ASAP7_75t_SL g3009 ( 
.A(n_2967),
.Y(n_3009)
);

OR2x2_ASAP7_75t_L g3010 ( 
.A(n_2992),
.B(n_2930),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_2974),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2981),
.B(n_2940),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2988),
.B(n_2949),
.Y(n_3013)
);

AOI21xp5_ASAP7_75t_L g3014 ( 
.A1(n_2986),
.A2(n_2984),
.B(n_2981),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2985),
.B(n_2962),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2965),
.B(n_2918),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2984),
.B(n_2918),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2966),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2990),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2979),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2977),
.B(n_2949),
.Y(n_3021)
);

AND2x4_ASAP7_75t_L g3022 ( 
.A(n_2989),
.B(n_2944),
.Y(n_3022)
);

HB1xp67_ASAP7_75t_L g3023 ( 
.A(n_2964),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2971),
.B(n_2923),
.Y(n_3024)
);

OR2x2_ASAP7_75t_L g3025 ( 
.A(n_2973),
.B(n_2938),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2991),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2969),
.B(n_2941),
.Y(n_3027)
);

BUFx2_ASAP7_75t_L g3028 ( 
.A(n_2986),
.Y(n_3028)
);

OR2x2_ASAP7_75t_L g3029 ( 
.A(n_2993),
.B(n_2952),
.Y(n_3029)
);

A2O1A1Ixp33_ASAP7_75t_L g3030 ( 
.A1(n_3014),
.A2(n_2886),
.B(n_2874),
.C(n_2921),
.Y(n_3030)
);

NOR3xp33_ASAP7_75t_SL g3031 ( 
.A(n_3011),
.B(n_2766),
.C(n_2756),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_3011),
.B(n_2888),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_3023),
.B(n_2941),
.Y(n_3033)
);

OAI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_3028),
.A2(n_2886),
.B1(n_2888),
.B2(n_2905),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2998),
.B(n_3020),
.Y(n_3035)
);

OAI22xp33_ASAP7_75t_SL g3036 ( 
.A1(n_3028),
.A2(n_2701),
.B1(n_2886),
.B2(n_2921),
.Y(n_3036)
);

AOI21xp33_ASAP7_75t_L g3037 ( 
.A1(n_2996),
.A2(n_2717),
.B(n_2753),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2996),
.A2(n_2701),
.B(n_2748),
.Y(n_3038)
);

AOI211xp5_ASAP7_75t_L g3039 ( 
.A1(n_3017),
.A2(n_2712),
.B(n_2690),
.C(n_2750),
.Y(n_3039)
);

NOR3xp33_ASAP7_75t_L g3040 ( 
.A(n_3009),
.B(n_2832),
.C(n_2805),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_3002),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_3012),
.B(n_3017),
.Y(n_3042)
);

CKINVDCx20_ASAP7_75t_R g3043 ( 
.A(n_3026),
.Y(n_3043)
);

AND3x1_ASAP7_75t_L g3044 ( 
.A(n_3001),
.B(n_3012),
.C(n_3026),
.Y(n_3044)
);

OAI22xp5_ASAP7_75t_L g3045 ( 
.A1(n_3025),
.A2(n_2888),
.B1(n_2959),
.B2(n_2934),
.Y(n_3045)
);

OAI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_3025),
.A2(n_3024),
.B1(n_3021),
.B2(n_3015),
.Y(n_3046)
);

INVxp33_ASAP7_75t_L g3047 ( 
.A(n_3022),
.Y(n_3047)
);

HB1xp67_ASAP7_75t_L g3048 ( 
.A(n_3029),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_3018),
.B(n_2934),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2999),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_3019),
.Y(n_3051)
);

INVxp67_ASAP7_75t_L g3052 ( 
.A(n_3022),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_3027),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_3015),
.B(n_2925),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_3004),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_3048),
.B(n_2997),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_3050),
.B(n_2997),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_3047),
.B(n_3008),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3033),
.Y(n_3059)
);

INVx2_ASAP7_75t_SL g3060 ( 
.A(n_3032),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_3052),
.B(n_3008),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_3043),
.Y(n_3062)
);

NOR2x1_ASAP7_75t_L g3063 ( 
.A(n_3030),
.B(n_3022),
.Y(n_3063)
);

NOR3xp33_ASAP7_75t_L g3064 ( 
.A(n_3052),
.B(n_3007),
.C(n_3016),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_3054),
.B(n_3006),
.Y(n_3065)
);

OR2x2_ASAP7_75t_L g3066 ( 
.A(n_3041),
.B(n_3035),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_3051),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_3042),
.B(n_3006),
.Y(n_3068)
);

AOI221xp5_ASAP7_75t_L g3069 ( 
.A1(n_3044),
.A2(n_3007),
.B1(n_3016),
.B2(n_3000),
.C(n_2995),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_3055),
.B(n_3010),
.Y(n_3070)
);

OR2x2_ASAP7_75t_L g3071 ( 
.A(n_3053),
.B(n_3029),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_3046),
.B(n_3010),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_3039),
.B(n_2995),
.Y(n_3073)
);

OAI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_3031),
.A2(n_3003),
.B1(n_3013),
.B2(n_3005),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_3040),
.B(n_2925),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3071),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_3062),
.Y(n_3077)
);

INVx2_ASAP7_75t_SL g3078 ( 
.A(n_3060),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_3072),
.B(n_3036),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_3058),
.Y(n_3080)
);

INVx2_ASAP7_75t_SL g3081 ( 
.A(n_3063),
.Y(n_3081)
);

HB1xp67_ASAP7_75t_L g3082 ( 
.A(n_3067),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3061),
.B(n_3040),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_3056),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3056),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3064),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3070),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_3070),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3066),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_3057),
.Y(n_3090)
);

INVx2_ASAP7_75t_SL g3091 ( 
.A(n_3073),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_L g3092 ( 
.A(n_3059),
.B(n_3045),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3057),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3068),
.Y(n_3094)
);

OAI22xp5_ASAP7_75t_SL g3095 ( 
.A1(n_3078),
.A2(n_3074),
.B1(n_3069),
.B2(n_3049),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3077),
.B(n_3075),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_SL g3097 ( 
.A1(n_3081),
.A2(n_3074),
.B(n_3038),
.Y(n_3097)
);

NAND3xp33_ASAP7_75t_L g3098 ( 
.A(n_3086),
.B(n_3037),
.C(n_3065),
.Y(n_3098)
);

NAND3xp33_ASAP7_75t_L g3099 ( 
.A(n_3084),
.B(n_3034),
.C(n_2730),
.Y(n_3099)
);

NOR2x1_ASAP7_75t_L g3100 ( 
.A(n_3085),
.B(n_2905),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_3091),
.B(n_2931),
.Y(n_3101)
);

AOI221xp5_ASAP7_75t_L g3102 ( 
.A1(n_3076),
.A2(n_3083),
.B1(n_3087),
.B2(n_3088),
.C(n_3094),
.Y(n_3102)
);

NAND4xp25_ASAP7_75t_L g3103 ( 
.A(n_3079),
.B(n_2771),
.C(n_2777),
.D(n_2799),
.Y(n_3103)
);

OAI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_3083),
.A2(n_2888),
.B1(n_2905),
.B2(n_2752),
.Y(n_3104)
);

AOI221xp5_ASAP7_75t_L g3105 ( 
.A1(n_3080),
.A2(n_2759),
.B1(n_2840),
.B2(n_2814),
.C(n_2815),
.Y(n_3105)
);

NOR3xp33_ASAP7_75t_L g3106 ( 
.A(n_3089),
.B(n_2695),
.C(n_2643),
.Y(n_3106)
);

NAND4xp25_ASAP7_75t_L g3107 ( 
.A(n_3092),
.B(n_3093),
.C(n_3090),
.D(n_3082),
.Y(n_3107)
);

OAI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_3098),
.A2(n_3092),
.B(n_3082),
.Y(n_3108)
);

AOI22xp5_ASAP7_75t_L g3109 ( 
.A1(n_3095),
.A2(n_2959),
.B1(n_2946),
.B2(n_2752),
.Y(n_3109)
);

AOI211xp5_ASAP7_75t_L g3110 ( 
.A1(n_3107),
.A2(n_2757),
.B(n_2762),
.C(n_2797),
.Y(n_3110)
);

OAI221xp5_ASAP7_75t_L g3111 ( 
.A1(n_3103),
.A2(n_2696),
.B1(n_2797),
.B2(n_2779),
.C(n_2888),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_3097),
.A2(n_2692),
.B(n_2556),
.Y(n_3112)
);

XNOR2xp5_ASAP7_75t_L g3113 ( 
.A(n_3096),
.B(n_2959),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_3106),
.A2(n_2946),
.B1(n_2755),
.B2(n_2802),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_3102),
.A2(n_2937),
.B(n_2935),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_3105),
.B(n_3101),
.Y(n_3116)
);

NAND2x1p5_ASAP7_75t_SL g3117 ( 
.A(n_3108),
.B(n_3100),
.Y(n_3117)
);

INVxp67_ASAP7_75t_L g3118 ( 
.A(n_3116),
.Y(n_3118)
);

OR2x2_ASAP7_75t_L g3119 ( 
.A(n_3112),
.B(n_3109),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_3113),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_3115),
.B(n_3104),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_R g3122 ( 
.A(n_3120),
.B(n_3110),
.Y(n_3122)
);

NAND3xp33_ASAP7_75t_L g3123 ( 
.A(n_3118),
.B(n_3111),
.C(n_3099),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_R g3124 ( 
.A(n_3119),
.B(n_3114),
.Y(n_3124)
);

NAND3xp33_ASAP7_75t_L g3125 ( 
.A(n_3121),
.B(n_2956),
.C(n_2863),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_3117),
.B(n_2863),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_3126),
.Y(n_3127)
);

OAI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_3123),
.A2(n_2961),
.B(n_2958),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_3124),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_3122),
.B(n_2906),
.Y(n_3130)
);

OAI21xp5_ASAP7_75t_SL g3131 ( 
.A1(n_3129),
.A2(n_3127),
.B(n_3130),
.Y(n_3131)
);

OAI31xp33_ASAP7_75t_L g3132 ( 
.A1(n_3128),
.A2(n_3125),
.A3(n_2709),
.B(n_2958),
.Y(n_3132)
);

HB1xp67_ASAP7_75t_L g3133 ( 
.A(n_3131),
.Y(n_3133)
);

AOI31xp33_ASAP7_75t_L g3134 ( 
.A1(n_3133),
.A2(n_3132),
.A3(n_2961),
.B(n_2855),
.Y(n_3134)
);

INVx1_ASAP7_75t_SL g3135 ( 
.A(n_3134),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_SL g3136 ( 
.A1(n_3135),
.A2(n_2951),
.B1(n_2953),
.B2(n_2791),
.Y(n_3136)
);

INVx4_ASAP7_75t_L g3137 ( 
.A(n_3136),
.Y(n_3137)
);

AOI221xp5_ASAP7_75t_L g3138 ( 
.A1(n_3137),
.A2(n_2953),
.B1(n_2951),
.B2(n_2957),
.C(n_2955),
.Y(n_3138)
);

AOI211xp5_ASAP7_75t_L g3139 ( 
.A1(n_3138),
.A2(n_2957),
.B(n_2955),
.C(n_2761),
.Y(n_3139)
);


endmodule