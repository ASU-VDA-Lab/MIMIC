module fake_netlist_6_2794_n_1926 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1926);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1926;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_131),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_67),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_36),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_38),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_72),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_82),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_74),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_33),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_9),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_12),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_23),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_25),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_53),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_157),
.Y(n_216)
);

BUFx8_ASAP7_75t_SL g217 ( 
.A(n_140),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_76),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_88),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_66),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_122),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_91),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_105),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_51),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_70),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_126),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_28),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_113),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_169),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_26),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_53),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_2),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_161),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_176),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_84),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_103),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_142),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_114),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_69),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_79),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_124),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_57),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_181),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_125),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_25),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_107),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_46),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_185),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_94),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_56),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_12),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_75),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_166),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_95),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_36),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_63),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_28),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_31),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_96),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_151),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_115),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_137),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_42),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_98),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_89),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_167),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_49),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_170),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_16),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_62),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_59),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_153),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_13),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_56),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_31),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_64),
.Y(n_299)
);

BUFx2_ASAP7_75t_SL g300 ( 
.A(n_147),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_15),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_18),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_152),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_106),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_80),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_42),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_104),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_78),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_112),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_68),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_180),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_130),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_58),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_16),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_173),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_24),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_159),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_138),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_27),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_148),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_143),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_86),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_97),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_13),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_24),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_83),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_99),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_60),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_155),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_61),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_150),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_116),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_39),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_63),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_44),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_149),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_43),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_144),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_183),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_108),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_46),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_17),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_43),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_189),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_77),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_168),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_57),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_8),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_21),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_100),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_120),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_8),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_133),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_58),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_85),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_101),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_45),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_90),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_30),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_172),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_49),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_165),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_3),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_29),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_123),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_4),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_154),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_188),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_158),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_178),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_21),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_135),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_5),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_26),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_48),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_145),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_7),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_110),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_111),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_61),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_9),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_121),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_129),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_7),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_1),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_40),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_39),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_54),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_40),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_214),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_214),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_293),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_214),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_214),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_259),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_214),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_214),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_363),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_223),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_297),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_203),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_214),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_209),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_209),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_259),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_203),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_206),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_209),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_209),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_275),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_230),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_239),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_299),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_275),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_275),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_275),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_284),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_284),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_284),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_284),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_306),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_242),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_244),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_259),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_270),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_306),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_276),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_301),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_299),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_237),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_237),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_206),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_279),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_269),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_294),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_213),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_296),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_296),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_198),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_236),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_306),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_333),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_333),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_329),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_329),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_306),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_197),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_199),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_229),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_207),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_235),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_325),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_252),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_262),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_364),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_328),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_265),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_266),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_364),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_210),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_277),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_217),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_330),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_193),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_226),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_290),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_207),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_208),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_292),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_298),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_213),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_226),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_198),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_302),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_208),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_313),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_344),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_221),
.Y(n_482)
);

INVxp33_ASAP7_75t_SL g483 ( 
.A(n_221),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_344),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_308),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_210),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_316),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_336),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_331),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_319),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_308),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_196),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_466),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_432),
.A2(n_377),
.B1(n_379),
.B2(n_319),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_445),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_445),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_412),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_399),
.B(n_268),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_412),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_497),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_443),
.B(n_196),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_268),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_396),
.A2(n_243),
.B1(n_324),
.B2(n_274),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_405),
.A2(n_274),
.B1(n_324),
.B2(n_243),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_468),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_414),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_418),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_418),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_464),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_410),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_464),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_464),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_403),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_273),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_402),
.B(n_273),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_420),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_487),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_417),
.A2(n_353),
.B1(n_361),
.B2(n_345),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_444),
.B(n_196),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_409),
.B(n_201),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_487),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_411),
.B(n_241),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_454),
.B(n_303),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_487),
.B(n_210),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_398),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_497),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_415),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_R g555 ( 
.A(n_415),
.B(n_194),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_433),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_416),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_416),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_426),
.B(n_427),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_401),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_424),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_404),
.A2(n_377),
.B1(n_379),
.B2(n_381),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_401),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_472),
.B(n_238),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_479),
.A2(n_345),
.B1(n_353),
.B2(n_361),
.Y(n_569)
);

OA21x2_ASAP7_75t_L g570 ( 
.A1(n_394),
.A2(n_256),
.B(n_255),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_428),
.B(n_255),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_425),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_427),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_486),
.B(n_201),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_448),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_406),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_449),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_434),
.B(n_256),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_425),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_430),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_430),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_450),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_550),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_300),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_550),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_507),
.A2(n_380),
.B1(n_278),
.B2(n_368),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_505),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_516),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_507),
.B(n_469),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_561),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_561),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_547),
.B(n_429),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_561),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_561),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_566),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_566),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_548),
.A2(n_431),
.B1(n_437),
.B2(n_429),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_550),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_511),
.B(n_552),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_566),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_566),
.Y(n_605)
);

CKINVDCx6p67_ASAP7_75t_R g606 ( 
.A(n_556),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_513),
.A2(n_338),
.B1(n_340),
.B2(n_337),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_507),
.B(n_533),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_509),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_394),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_549),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_518),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_525),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_568),
.B(n_483),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_553),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_507),
.B(n_395),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_501),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_501),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_552),
.B(n_494),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_278),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_529),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_529),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_502),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_550),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_526),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_550),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_518),
.B(n_431),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_560),
.Y(n_636)
);

AO21x2_ASAP7_75t_L g637 ( 
.A1(n_532),
.A2(n_200),
.B(n_192),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_512),
.B(n_397),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_560),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_570),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_543),
.A2(n_439),
.B1(n_456),
.B2(n_437),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_504),
.Y(n_643)
);

BUFx4f_ASAP7_75t_L g644 ( 
.A(n_570),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_543),
.B(n_400),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_504),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_570),
.A2(n_400),
.B(n_406),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_516),
.B(n_475),
.C(n_440),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_555),
.B(n_439),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_R g651 ( 
.A(n_499),
.B(n_517),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_559),
.B(n_456),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_542),
.B(n_460),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_556),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_574),
.B(n_460),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_506),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_560),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_574),
.B(n_467),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_510),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_560),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_531),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_557),
.B(n_467),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_571),
.A2(n_385),
.B1(n_389),
.B2(n_380),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_560),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_523),
.B(n_492),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_546),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_523),
.B(n_492),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_578),
.A2(n_212),
.B(n_204),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_536),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_576),
.B(n_195),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_558),
.B(n_436),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_536),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_526),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_508),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g678 ( 
.A(n_569),
.B(n_459),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_563),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_571),
.B(n_469),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_575),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_571),
.B(n_582),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_526),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_526),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_538),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_573),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_576),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_576),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_565),
.B(n_201),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_515),
.A2(n_482),
.B1(n_471),
.B2(n_452),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_538),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_515),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_500),
.B(n_225),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_549),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_577),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_576),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_519),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_514),
.B(n_225),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_519),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_576),
.B(n_202),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_508),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_551),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_562),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_562),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_564),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_564),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_582),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_520),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_520),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_581),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_521),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_581),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_SL g716 ( 
.A(n_540),
.B(n_365),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_521),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_528),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_527),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_527),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_527),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_528),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_527),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_508),
.B(n_224),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_535),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_535),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_539),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_508),
.B(n_227),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_544),
.B(n_476),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_544),
.B(n_476),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_527),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_524),
.B(n_231),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_608),
.B(n_291),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_646),
.B(n_524),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_621),
.B(n_291),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_621),
.B(n_291),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_614),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_616),
.B(n_569),
.C(n_514),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_677),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_614),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_653),
.B(n_435),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_639),
.A2(n_453),
.B(n_455),
.C(n_451),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_614),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_619),
.A2(n_458),
.B(n_461),
.C(n_457),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_617),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_592),
.B(n_524),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_625),
.A2(n_232),
.B1(n_222),
.B2(n_463),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_592),
.B(n_524),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_621),
.B(n_291),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_680),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_710),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_644),
.A2(n_233),
.B(n_228),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_682),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_711),
.B(n_541),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_682),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_662),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_641),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_662),
.B(n_438),
.Y(n_759)
);

OAI22xp33_ASAP7_75t_L g760 ( 
.A1(n_716),
.A2(n_378),
.B1(n_365),
.B2(n_381),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_668),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_711),
.B(n_541),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_596),
.B(n_642),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_674),
.Y(n_765)
);

INVx8_ASAP7_75t_L g766 ( 
.A(n_586),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_611),
.B(n_541),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_624),
.B(n_601),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_641),
.A2(n_447),
.B(n_441),
.C(n_442),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_668),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_644),
.A2(n_537),
.B(n_534),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_679),
.B(n_446),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_717),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_611),
.B(n_541),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_611),
.B(n_554),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_679),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_644),
.B(n_371),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_718),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_611),
.B(n_554),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_656),
.B(n_205),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_659),
.B(n_205),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_686),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_641),
.B(n_371),
.Y(n_783)
);

NOR2x1p5_ASAP7_75t_L g784 ( 
.A(n_606),
.B(n_346),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_729),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_625),
.A2(n_287),
.B1(n_387),
.B2(n_386),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_625),
.A2(n_286),
.B1(n_383),
.B2(n_382),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_730),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_625),
.B(n_567),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_686),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_663),
.B(n_462),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_594),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_594),
.Y(n_793)
);

INVx5_ASAP7_75t_L g794 ( 
.A(n_645),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_635),
.B(n_572),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_595),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_730),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_689),
.B(n_694),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_718),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_595),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_615),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_625),
.B(n_579),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_591),
.A2(n_378),
.B1(n_347),
.B2(n_351),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_598),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_648),
.B(n_371),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_617),
.B(n_213),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_588),
.A2(n_250),
.B1(n_251),
.B2(n_234),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_586),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_650),
.B(n_211),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_645),
.B(n_245),
.Y(n_810)
);

AO221x1_ASAP7_75t_L g811 ( 
.A1(n_607),
.A2(n_371),
.B1(n_240),
.B2(n_247),
.C(n_248),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_609),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_612),
.B(n_692),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_652),
.B(n_211),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_612),
.B(n_253),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_609),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_701),
.B(n_215),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_617),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_645),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_598),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_618),
.B(n_579),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_654),
.B(n_580),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_617),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_618),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_677),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_620),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_588),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_645),
.B(n_246),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_585),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_620),
.B(n_622),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_599),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_588),
.A2(n_288),
.B1(n_280),
.B2(n_282),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_588),
.A2(n_637),
.B1(n_628),
.B2(n_630),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_612),
.B(n_692),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_622),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_628),
.B(n_580),
.Y(n_836)
);

BUFx6f_ASAP7_75t_SL g837 ( 
.A(n_586),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_586),
.B(n_215),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_645),
.B(n_249),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_630),
.B(n_285),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_643),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_599),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_681),
.B(n_465),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_643),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_654),
.B(n_470),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_612),
.B(n_307),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_647),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_647),
.B(n_318),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_655),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_655),
.B(n_322),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_657),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_657),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_660),
.B(n_254),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_660),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_586),
.B(n_216),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_612),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_603),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_600),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_693),
.B(n_366),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_693),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_704),
.A2(n_374),
.B1(n_315),
.B2(n_220),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_700),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_700),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_585),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_667),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_637),
.A2(n_272),
.B1(n_258),
.B2(n_260),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_702),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_712),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_712),
.B(n_530),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_692),
.B(n_261),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_714),
.B(n_216),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_714),
.B(n_530),
.Y(n_872)
);

AOI221xp5_ASAP7_75t_L g873 ( 
.A1(n_699),
.A2(n_358),
.B1(n_356),
.B2(n_352),
.C(n_370),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_692),
.B(n_263),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_589),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_589),
.Y(n_876)
);

BUFx5_ASAP7_75t_L g877 ( 
.A(n_597),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_722),
.B(n_530),
.Y(n_878)
);

BUFx6f_ASAP7_75t_SL g879 ( 
.A(n_606),
.Y(n_879)
);

CKINVDCx16_ASAP7_75t_R g880 ( 
.A(n_651),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_637),
.A2(n_314),
.B1(n_264),
.B2(n_478),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_722),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_725),
.B(n_530),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_696),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_725),
.B(n_267),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_726),
.B(n_530),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_726),
.B(n_530),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_605),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_690),
.B(n_264),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_692),
.B(n_271),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_669),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_727),
.B(n_218),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_727),
.B(n_545),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_649),
.B(n_264),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_863),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_863),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_754),
.B(n_719),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_764),
.A2(n_732),
.B1(n_728),
.B2(n_724),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_773),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_760),
.B(n_678),
.C(n_696),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_776),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_758),
.B(n_673),
.Y(n_902)
);

INVx5_ASAP7_75t_L g903 ( 
.A(n_794),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_765),
.B(n_678),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_812),
.B(n_703),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_818),
.B(n_823),
.Y(n_906)
);

BUFx4f_ASAP7_75t_L g907 ( 
.A(n_766),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_782),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_829),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_756),
.B(n_719),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_740),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_770),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_753),
.B(n_695),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_829),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_790),
.Y(n_915)
);

AND3x1_ASAP7_75t_SL g916 ( 
.A(n_873),
.B(n_474),
.C(n_473),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_770),
.Y(n_917)
);

OAI22xp33_ASAP7_75t_L g918 ( 
.A1(n_738),
.A2(n_391),
.B1(n_384),
.B2(n_388),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_778),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_880),
.B(n_225),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_864),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_764),
.B(n_695),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_799),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_733),
.A2(n_670),
.B(n_638),
.C(n_665),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_799),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_739),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_748),
.Y(n_927)
);

OAI22xp33_ASAP7_75t_L g928 ( 
.A1(n_768),
.A2(n_375),
.B1(n_715),
.B2(n_713),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_751),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_816),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_739),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_824),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_801),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_794),
.B(n_695),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_826),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_843),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_768),
.A2(n_658),
.B1(n_666),
.B2(n_602),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_827),
.A2(n_664),
.B1(n_671),
.B2(n_706),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_865),
.B(n_602),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_801),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_891),
.B(n_670),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_827),
.A2(n_623),
.B1(n_715),
.B2(n_713),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_752),
.B(n_602),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_835),
.B(n_597),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_864),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_757),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_759),
.B(n_314),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_740),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_841),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_844),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_794),
.B(n_695),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_772),
.B(n_602),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_798),
.B(n_631),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_847),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_875),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_794),
.A2(n_587),
.B(n_583),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_811),
.A2(n_626),
.B1(n_675),
.B2(n_685),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_849),
.Y(n_958)
);

INVx8_ASAP7_75t_L g959 ( 
.A(n_766),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_851),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_852),
.B(n_604),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_854),
.B(n_604),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_875),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_761),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_798),
.B(n_631),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_806),
.B(n_314),
.Y(n_966)
);

AO22x1_ASAP7_75t_L g967 ( 
.A1(n_817),
.A2(n_220),
.B1(n_219),
.B2(n_218),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_876),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_763),
.A2(n_633),
.B1(n_658),
.B2(n_665),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_860),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_884),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_785),
.A2(n_666),
.B1(n_631),
.B2(n_633),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_788),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_862),
.B(n_631),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_871),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_735),
.A2(n_731),
.B(n_719),
.C(n_721),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_817),
.B(n_315),
.C(n_219),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_867),
.B(n_633),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_868),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_877),
.B(n_633),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_882),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_805),
.A2(n_807),
.B1(n_832),
.B2(n_760),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_775),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_791),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_797),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_825),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_830),
.B(n_795),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_803),
.B(n_317),
.C(n_480),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_877),
.B(n_638),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_871),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_805),
.A2(n_629),
.B1(n_675),
.B2(n_685),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_780),
.B(n_638),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_745),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_892),
.B(n_741),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_876),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_792),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_793),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_779),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_796),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_892),
.B(n_638),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_877),
.B(n_658),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_800),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_746),
.Y(n_1003)
);

NAND2x2_ASAP7_75t_L g1004 ( 
.A(n_784),
.B(n_257),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_804),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_749),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_877),
.B(n_658),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_737),
.B(n_665),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_821),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_836),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_820),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_743),
.B(n_665),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_791),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_831),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_780),
.B(n_666),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_879),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_842),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_889),
.B(n_495),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_879),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_783),
.B(n_687),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_791),
.Y(n_1021)
);

AND2x6_ASAP7_75t_SL g1022 ( 
.A(n_894),
.B(n_489),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_766),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_869),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_858),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_747),
.B(n_789),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_845),
.B(n_489),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_819),
.A2(n_587),
.B(n_583),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_781),
.B(n_687),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_808),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_872),
.Y(n_1031)
);

OR2x2_ASAP7_75t_SL g1032 ( 
.A(n_803),
.B(n_490),
.Y(n_1032)
);

BUFx8_ASAP7_75t_L g1033 ( 
.A(n_837),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_823),
.B(n_490),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_888),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_767),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_734),
.B(n_687),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_857),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_781),
.B(n_687),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_807),
.A2(n_626),
.B1(n_629),
.B2(n_671),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_878),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_809),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_883),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_809),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_814),
.B(n_491),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_822),
.B(n_774),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_755),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_832),
.A2(n_623),
.B1(n_627),
.B2(n_698),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_814),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_833),
.B(n_697),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_819),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_886),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_802),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_840),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_848),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_887),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_893),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_762),
.Y(n_1058)
);

AND2x6_ASAP7_75t_L g1059 ( 
.A(n_838),
.B(n_720),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_850),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_855),
.B(n_697),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_833),
.B(n_697),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_837),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_859),
.B(n_697),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_866),
.B(n_583),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_881),
.B(n_735),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_881),
.B(n_723),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_736),
.B(n_723),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_769),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_SL g1070 ( 
.A(n_1042),
.B(n_988),
.C(n_994),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1009),
.B(n_736),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_975),
.A2(n_769),
.B(n_733),
.C(n_742),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_973),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1010),
.B(n_750),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_903),
.A2(n_777),
.B(n_750),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_904),
.A2(n_853),
.B1(n_885),
.B2(n_787),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1044),
.B(n_861),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_988),
.A2(n_777),
.B1(n_874),
.B2(n_870),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_904),
.A2(n_786),
.B1(n_874),
.B2(n_870),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_903),
.A2(n_856),
.B(n_828),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_901),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1049),
.B(n_744),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1028),
.A2(n_771),
.B(n_890),
.Y(n_1083)
);

CKINVDCx14_ASAP7_75t_R g1084 ( 
.A(n_971),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_SL g1085 ( 
.A1(n_975),
.A2(n_990),
.B(n_922),
.C(n_1065),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_903),
.A2(n_856),
.B(n_839),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_990),
.B(n_610),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_992),
.A2(n_810),
.B(n_627),
.C(n_691),
.Y(n_1088)
);

NAND3xp33_ASAP7_75t_SL g1089 ( 
.A(n_920),
.B(n_317),
.C(n_283),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_903),
.A2(n_834),
.B(n_813),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1046),
.A2(n_321),
.B1(n_281),
.B2(n_289),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_908),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_912),
.B(n_583),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1051),
.A2(n_834),
.B(n_813),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1066),
.A2(n_983),
.B(n_998),
.C(n_982),
.Y(n_1095)
);

AO22x1_ASAP7_75t_L g1096 ( 
.A1(n_966),
.A2(n_933),
.B1(n_915),
.B2(n_917),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1050),
.A2(n_846),
.B(n_815),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_987),
.A2(n_691),
.B(n_613),
.C(n_698),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_973),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_985),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_909),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_982),
.A2(n_846),
.B(n_815),
.C(n_731),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_985),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_930),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_895),
.B(n_295),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_R g1106 ( 
.A(n_993),
.B(n_304),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_940),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_912),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_928),
.A2(n_706),
.B(n_705),
.C(n_707),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_953),
.A2(n_731),
.B(n_721),
.C(n_720),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_917),
.B(n_587),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_928),
.A2(n_705),
.B(n_707),
.C(n_708),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1054),
.B(n_305),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_947),
.B(n_493),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1045),
.A2(n_707),
.B(n_708),
.C(n_709),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1055),
.B(n_309),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_911),
.B(n_310),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_902),
.A2(n_640),
.B(n_661),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1003),
.B(n_709),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_953),
.A2(n_721),
.B(n_720),
.C(n_605),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1065),
.A2(n_593),
.B(n_590),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1006),
.B(n_590),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_1038),
.B(n_311),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_913),
.A2(n_640),
.B(n_634),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1060),
.B(n_723),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_911),
.B(n_312),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_932),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1021),
.B(n_636),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_986),
.Y(n_1130)
);

AO22x1_ASAP7_75t_L g1131 ( 
.A1(n_984),
.A2(n_327),
.B1(n_326),
.B2(n_323),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_946),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1046),
.A2(n_369),
.B1(n_320),
.B2(n_334),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_977),
.B(n_335),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_1016),
.B(n_339),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_913),
.A2(n_688),
.B(n_636),
.Y(n_1136)
);

AOI22x1_ASAP7_75t_L g1137 ( 
.A1(n_1069),
.A2(n_661),
.B1(n_688),
.B2(n_372),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_986),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_946),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_911),
.B(n_343),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1015),
.A2(n_1029),
.B1(n_1039),
.B2(n_965),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_914),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_948),
.B(n_348),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_948),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1019),
.B(n_257),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_921),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1026),
.A2(n_688),
.B(n_684),
.Y(n_1147)
);

AO22x1_ASAP7_75t_L g1148 ( 
.A1(n_1013),
.A2(n_359),
.B1(n_376),
.B2(n_373),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1047),
.B(n_349),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_927),
.B(n_481),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_945),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_965),
.A2(n_1029),
.B(n_1039),
.C(n_1015),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_948),
.Y(n_1153)
);

BUFx5_ASAP7_75t_L g1154 ( 
.A(n_897),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1063),
.B(n_350),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1026),
.A2(n_684),
.B(n_683),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1061),
.A2(n_360),
.B(n_354),
.C(n_355),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_948),
.B(n_896),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_905),
.A2(n_481),
.B(n_485),
.C(n_484),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1021),
.A2(n_357),
.B1(n_362),
.B2(n_341),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_935),
.A2(n_485),
.B(n_488),
.C(n_341),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_1063),
.B(n_257),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_949),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_955),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1061),
.A2(n_1062),
.B1(n_1053),
.B2(n_1000),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_964),
.B(n_332),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1032),
.A2(n_488),
.B1(n_341),
.B2(n_342),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_950),
.A2(n_954),
.B(n_979),
.C(n_970),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1053),
.B(n_332),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1053),
.A2(n_937),
.B1(n_1067),
.B2(n_952),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1053),
.B(n_332),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_898),
.A2(n_684),
.B(n_683),
.C(n_676),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1030),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_939),
.A2(n_676),
.B(n_672),
.C(n_632),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_963),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_SL g1176 ( 
.A(n_907),
.B(n_342),
.Y(n_1176)
);

AND3x1_ASAP7_75t_SL g1177 ( 
.A(n_900),
.B(n_929),
.C(n_958),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_960),
.B(n_584),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_952),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1030),
.Y(n_1180)
);

OAI21xp33_ASAP7_75t_SL g1181 ( 
.A1(n_981),
.A2(n_342),
.B(n_3),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_939),
.B(n_676),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_918),
.B(n_676),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1023),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_907),
.B(n_672),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1034),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_672),
.B1(n_632),
.B2(n_584),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1020),
.A2(n_549),
.B(n_537),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_899),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_956),
.A2(n_632),
.B(n_584),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_SL g1191 ( 
.A1(n_980),
.A2(n_81),
.B(n_191),
.C(n_179),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_SL g1192 ( 
.A1(n_957),
.A2(n_632),
.B(n_584),
.C(n_65),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1058),
.B(n_584),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_918),
.B(n_1),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_944),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1022),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1036),
.B(n_545),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_SL g1198 ( 
.A(n_1023),
.B(n_545),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1033),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1034),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1023),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_919),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_943),
.A2(n_545),
.B(n_10),
.C(n_14),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_980),
.A2(n_537),
.B(n_534),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1107),
.B(n_1023),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1141),
.A2(n_1043),
.B(n_1024),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1172),
.A2(n_924),
.B(n_957),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1194),
.A2(n_916),
.B1(n_1059),
.B2(n_943),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1174),
.A2(n_1037),
.B(n_1064),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1070),
.B(n_967),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1081),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1152),
.A2(n_991),
.B(n_941),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1128),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1163),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1114),
.B(n_906),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1108),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1095),
.B(n_1031),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1085),
.A2(n_991),
.B(n_1068),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1121),
.A2(n_974),
.B(n_978),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1170),
.A2(n_1041),
.B(n_1057),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1092),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1189),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1083),
.A2(n_989),
.B(n_1001),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1165),
.A2(n_1056),
.A3(n_1052),
.B(n_925),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1101),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1110),
.A2(n_962),
.B(n_961),
.Y(n_1226)
);

AO32x2_ASAP7_75t_L g1227 ( 
.A1(n_1167),
.A2(n_916),
.A3(n_1059),
.B1(n_976),
.B2(n_942),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_R g1228 ( 
.A(n_1084),
.B(n_959),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_1183),
.A2(n_1008),
.B(n_1012),
.Y(n_1229)
);

AO21x1_ASAP7_75t_L g1230 ( 
.A1(n_1072),
.A2(n_1074),
.B(n_1071),
.Y(n_1230)
);

NAND2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1184),
.B(n_986),
.Y(n_1231)
);

OA21x2_ASAP7_75t_L g1232 ( 
.A1(n_1120),
.A2(n_923),
.B(n_972),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1179),
.B(n_1036),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1075),
.A2(n_951),
.B(n_934),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1070),
.A2(n_1036),
.B1(n_1002),
.B2(n_1025),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1147),
.A2(n_989),
.B(n_1007),
.Y(n_1236)
);

NAND2x2_ASAP7_75t_L g1237 ( 
.A(n_1173),
.B(n_1004),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1124),
.A2(n_1007),
.B(n_1001),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1199),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1076),
.A2(n_942),
.B1(n_931),
.B2(n_926),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1079),
.A2(n_969),
.B(n_1017),
.C(n_1035),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1184),
.B(n_986),
.Y(n_1242)
);

BUFx8_ASAP7_75t_L g1243 ( 
.A(n_1132),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1078),
.A2(n_938),
.B1(n_1048),
.B2(n_1040),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1144),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1139),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1139),
.B(n_1033),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1072),
.A2(n_1048),
.B(n_1040),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1136),
.A2(n_995),
.B(n_968),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1190),
.A2(n_926),
.B(n_931),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1102),
.A2(n_938),
.B(n_897),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1087),
.B(n_1077),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1082),
.A2(n_1014),
.B(n_1011),
.C(n_1005),
.Y(n_1253)
);

AOI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1182),
.A2(n_999),
.B(n_897),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1149),
.B(n_996),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1153),
.B(n_1180),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1073),
.B(n_997),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1112),
.A2(n_910),
.B(n_897),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1088),
.A2(n_1118),
.B(n_1086),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1168),
.A2(n_959),
.B(n_910),
.C(n_1004),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1168),
.A2(n_910),
.B(n_87),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1080),
.A2(n_537),
.B(n_534),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1099),
.B(n_910),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1197),
.A2(n_175),
.B(n_163),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1176),
.B(n_6),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1203),
.B(n_10),
.C(n_15),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1100),
.B(n_17),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1166),
.B(n_18),
.Y(n_1268)
);

OAI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_1145),
.A2(n_19),
.B(n_20),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1202),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1157),
.A2(n_19),
.A3(n_20),
.B(n_22),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1089),
.A2(n_22),
.B(n_23),
.C(n_27),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1103),
.B(n_30),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1186),
.B(n_32),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1201),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1109),
.A2(n_141),
.B(n_139),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_1161),
.B(n_32),
.C(n_34),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1119),
.A2(n_35),
.A3(n_37),
.B(n_38),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1097),
.A2(n_119),
.B(n_117),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1096),
.B(n_37),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1200),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1153),
.B(n_1150),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1093),
.B(n_41),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1094),
.A2(n_41),
.B(n_47),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1177),
.A2(n_1089),
.B1(n_1181),
.B2(n_1171),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1111),
.B(n_50),
.Y(n_1286)
);

NOR4xp25_ASAP7_75t_L g1287 ( 
.A(n_1195),
.B(n_52),
.C(n_54),
.D(n_55),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_SL g1288 ( 
.A(n_1201),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1162),
.B(n_55),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1193),
.A2(n_59),
.A3(n_62),
.B(n_1129),
.Y(n_1290)
);

AO22x2_ASAP7_75t_L g1291 ( 
.A1(n_1169),
.A2(n_1196),
.B1(n_1158),
.B2(n_1195),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1161),
.B(n_1160),
.C(n_1134),
.Y(n_1292)
);

AO21x1_ASAP7_75t_L g1293 ( 
.A1(n_1115),
.A2(n_1159),
.B(n_1098),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1192),
.A2(n_1090),
.B(n_1187),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1122),
.A2(n_1159),
.B(n_1126),
.Y(n_1296)
);

AOI221xp5_ASAP7_75t_L g1297 ( 
.A1(n_1131),
.A2(n_1148),
.B1(n_1106),
.B2(n_1135),
.C(n_1191),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1144),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1130),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1130),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1142),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1178),
.A2(n_1146),
.A3(n_1175),
.B(n_1164),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1151),
.B(n_1091),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1137),
.A2(n_1204),
.B(n_1188),
.Y(n_1304)
);

OAI22x1_ASAP7_75t_L g1305 ( 
.A1(n_1185),
.A2(n_1143),
.B1(n_1117),
.B2(n_1140),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1138),
.Y(n_1306)
);

NOR3xp33_ASAP7_75t_L g1307 ( 
.A(n_1127),
.B(n_1155),
.C(n_1105),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1138),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_L g1309 ( 
.A(n_1133),
.B(n_1123),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1154),
.B(n_1042),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1154),
.A2(n_1152),
.B(n_1141),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1154),
.A2(n_1042),
.B1(n_1152),
.B2(n_975),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1154),
.B(n_1042),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1121),
.A2(n_1083),
.B(n_1156),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1084),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1104),
.Y(n_1316)
);

AOI221x1_ASAP7_75t_L g1317 ( 
.A1(n_1141),
.A2(n_1152),
.B1(n_1194),
.B2(n_988),
.C(n_1172),
.Y(n_1317)
);

AO21x1_ASAP7_75t_L g1318 ( 
.A1(n_1141),
.A2(n_1066),
.B(n_1170),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1152),
.A2(n_1042),
.B1(n_975),
.B2(n_990),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1125),
.B(n_1114),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1199),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1194),
.B(n_768),
.C(n_764),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1144),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1152),
.A2(n_1141),
.B(n_1085),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1121),
.A2(n_1083),
.B(n_1156),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1070),
.B(n_936),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1081),
.B(n_681),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1125),
.B(n_975),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1201),
.Y(n_1329)
);

NAND2x1_ASAP7_75t_L g1330 ( 
.A(n_1184),
.B(n_1198),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1081),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1152),
.A2(n_1042),
.B1(n_975),
.B2(n_990),
.Y(n_1332)
);

NAND3xp33_ASAP7_75t_SL g1333 ( 
.A(n_1162),
.B(n_616),
.C(n_653),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1201),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1125),
.B(n_1042),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_SL g1336 ( 
.A(n_1194),
.B(n_880),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1121),
.A2(n_1083),
.B(n_1156),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1152),
.A2(n_1141),
.B(n_1085),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1125),
.B(n_975),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_L g1340 ( 
.A(n_1081),
.B(n_818),
.Y(n_1340)
);

NOR2xp67_ASAP7_75t_L g1341 ( 
.A(n_1070),
.B(n_936),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1125),
.B(n_1114),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1125),
.B(n_975),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1107),
.B(n_1023),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1324),
.A2(n_1338),
.B(n_1317),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1243),
.Y(n_1346)
);

AOI22x1_ASAP7_75t_L g1347 ( 
.A1(n_1305),
.A2(n_1291),
.B1(n_1284),
.B2(n_1276),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1320),
.B(n_1342),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1322),
.A2(n_1333),
.B1(n_1269),
.B2(n_1266),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1328),
.B(n_1339),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1282),
.B(n_1215),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1248),
.A2(n_1244),
.B(n_1212),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1322),
.A2(n_1292),
.B(n_1285),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1343),
.B(n_1335),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1287),
.A2(n_1266),
.B1(n_1269),
.B2(n_1268),
.C(n_1210),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1329),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1338),
.A2(n_1206),
.B(n_1220),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1216),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1205),
.B(n_1344),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1219),
.A2(n_1236),
.B(n_1249),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1336),
.A2(n_1277),
.B1(n_1318),
.B2(n_1289),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1312),
.B(n_1319),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1254),
.A2(n_1238),
.B(n_1304),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1239),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1246),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1251),
.A2(n_1311),
.B(n_1208),
.C(n_1272),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1205),
.B(n_1344),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1223),
.A2(n_1250),
.B(n_1234),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1252),
.B(n_1332),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1336),
.A2(n_1280),
.B1(n_1265),
.B2(n_1285),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1329),
.B(n_1245),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1326),
.A2(n_1341),
.B1(n_1208),
.B2(n_1294),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1292),
.A2(n_1217),
.B(n_1241),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1331),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1327),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1218),
.A2(n_1229),
.B(n_1311),
.Y(n_1378)
);

BUFx4_ASAP7_75t_SL g1379 ( 
.A(n_1315),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1302),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1251),
.A2(n_1277),
.B(n_1283),
.C(n_1286),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1213),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1218),
.A2(n_1293),
.B(n_1258),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1228),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1329),
.B(n_1245),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1256),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1243),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1233),
.B(n_1247),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1316),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1262),
.A2(n_1226),
.B(n_1296),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1226),
.A2(n_1296),
.B(n_1264),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1274),
.B(n_1301),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1209),
.A2(n_1207),
.B(n_1279),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1310),
.A2(n_1313),
.B(n_1230),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1222),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1209),
.A2(n_1207),
.B(n_1279),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1232),
.A2(n_1253),
.B(n_1240),
.Y(n_1397)
);

CKINVDCx8_ASAP7_75t_R g1398 ( 
.A(n_1221),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1302),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1270),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1281),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1211),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1255),
.A2(n_1303),
.B(n_1330),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1273),
.A2(n_1309),
.B1(n_1297),
.B2(n_1307),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1235),
.A2(n_1263),
.B(n_1300),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1300),
.A2(n_1308),
.B(n_1231),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1257),
.A2(n_1340),
.B1(n_1267),
.B2(n_1225),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1231),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1224),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1242),
.A2(n_1323),
.B(n_1224),
.Y(n_1410)
);

OAI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1287),
.A2(n_1237),
.B1(n_1260),
.B2(n_1299),
.C(n_1306),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1242),
.A2(n_1323),
.B(n_1224),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1227),
.A2(n_1290),
.B(n_1271),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1321),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1298),
.A2(n_1227),
.B(n_1271),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1227),
.A2(n_1271),
.B(n_1278),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1278),
.A2(n_1288),
.B(n_1298),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1278),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1334),
.A2(n_1333),
.B(n_768),
.C(n_1322),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1214),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1239),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1216),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1324),
.A2(n_1338),
.B(n_1317),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1322),
.A2(n_760),
.B1(n_768),
.B2(n_738),
.C(n_764),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1248),
.A2(n_753),
.B(n_1152),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1239),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1205),
.B(n_1344),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1324),
.A2(n_1338),
.B(n_1317),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1322),
.A2(n_653),
.B1(n_616),
.B2(n_768),
.C(n_764),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1214),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1214),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1214),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1329),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1214),
.Y(n_1435)
);

CKINVDCx6p67_ASAP7_75t_R g1436 ( 
.A(n_1239),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1239),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1322),
.B(n_616),
.C(n_768),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1328),
.B(n_1339),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1221),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1243),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1214),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1329),
.Y(n_1445)
);

OAI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1322),
.A2(n_653),
.B1(n_616),
.B2(n_768),
.C(n_764),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1239),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1322),
.A2(n_1333),
.B(n_768),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1231),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1322),
.A2(n_1333),
.B1(n_904),
.B2(n_1336),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1214),
.Y(n_1454)
);

AO31x2_ASAP7_75t_L g1455 ( 
.A1(n_1220),
.A2(n_1206),
.A3(n_1229),
.B(n_1318),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_SL g1456 ( 
.A1(n_1248),
.A2(n_1152),
.B(n_1276),
.C(n_1322),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_SL g1457 ( 
.A1(n_1261),
.A2(n_1220),
.B(n_1276),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1322),
.A2(n_1333),
.B(n_768),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1243),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1322),
.A2(n_1194),
.B1(n_988),
.B2(n_1333),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1322),
.B(n_904),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1322),
.A2(n_1333),
.B(n_768),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1243),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1320),
.B(n_1342),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1322),
.A2(n_768),
.B1(n_1042),
.B2(n_764),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1205),
.B(n_1344),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1216),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1322),
.A2(n_1194),
.B1(n_988),
.B2(n_1333),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1322),
.B(n_616),
.C(n_768),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1239),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1322),
.A2(n_768),
.B(n_764),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1314),
.A2(n_1337),
.B(n_1325),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1216),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1214),
.Y(n_1474)
);

BUFx4_ASAP7_75t_R g1475 ( 
.A(n_1275),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1216),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1259),
.A2(n_1295),
.B(n_1324),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1214),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1211),
.B(n_936),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1214),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1430),
.A2(n_1446),
.B(n_1465),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1360),
.B(n_1369),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1365),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1381),
.A2(n_1419),
.B(n_1426),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1439),
.A2(n_1469),
.B1(n_1425),
.B2(n_1349),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1354),
.B(n_1348),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1353),
.B(n_1352),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1471),
.A2(n_1458),
.B(n_1449),
.C(n_1462),
.Y(n_1488)
);

OAI31xp33_ASAP7_75t_L g1489 ( 
.A1(n_1461),
.A2(n_1372),
.A3(n_1468),
.B(n_1460),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1456),
.A2(n_1375),
.B(n_1368),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1381),
.B(n_1349),
.Y(n_1491)
);

OA22x2_ASAP7_75t_L g1492 ( 
.A1(n_1453),
.A2(n_1388),
.B1(n_1374),
.B2(n_1363),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1461),
.A2(n_1468),
.B(n_1460),
.C(n_1404),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1368),
.A2(n_1347),
.B(n_1363),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1356),
.B(n_1350),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1404),
.A2(n_1362),
.B1(n_1440),
.B2(n_1377),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1360),
.B(n_1369),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1359),
.B(n_1467),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1362),
.A2(n_1400),
.B1(n_1389),
.B2(n_1395),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1457),
.A2(n_1401),
.B1(n_1422),
.B2(n_1473),
.C(n_1407),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1393),
.A2(n_1396),
.B(n_1391),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1382),
.A2(n_1345),
.B1(n_1429),
.B2(n_1423),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1392),
.B(n_1386),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1345),
.A2(n_1429),
.B1(n_1423),
.B2(n_1388),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1393),
.A2(n_1396),
.B(n_1391),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1345),
.B(n_1423),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1476),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1442),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1369),
.B(n_1428),
.Y(n_1509)
);

AOI211xp5_ASAP7_75t_L g1510 ( 
.A1(n_1411),
.A2(n_1403),
.B(n_1479),
.C(n_1402),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1366),
.B(n_1376),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1429),
.B(n_1383),
.Y(n_1512)
);

INVx5_ASAP7_75t_L g1513 ( 
.A(n_1434),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1388),
.Y(n_1514)
);

INVx5_ASAP7_75t_L g1515 ( 
.A(n_1434),
.Y(n_1515)
);

CKINVDCx16_ASAP7_75t_R g1516 ( 
.A(n_1414),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1379),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1398),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1434),
.Y(n_1519)
);

CKINVDCx14_ASAP7_75t_R g1520 ( 
.A(n_1414),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1475),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1383),
.B(n_1378),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1420),
.A2(n_1480),
.B1(n_1478),
.B2(n_1431),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1466),
.B(n_1408),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1432),
.A2(n_1433),
.B(n_1454),
.C(n_1444),
.Y(n_1525)
);

AND2x2_ASAP7_75t_SL g1526 ( 
.A(n_1384),
.B(n_1475),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_R g1527 ( 
.A(n_1421),
.B(n_1470),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1435),
.A2(n_1474),
.B(n_1346),
.C(n_1477),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1387),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1451),
.B(n_1373),
.Y(n_1530)
);

O2A1O1Ixp5_ASAP7_75t_L g1531 ( 
.A1(n_1415),
.A2(n_1394),
.B(n_1409),
.C(n_1418),
.Y(n_1531)
);

NOR2xp67_ASAP7_75t_R g1532 ( 
.A(n_1427),
.B(n_1438),
.Y(n_1532)
);

NOR2xp67_ASAP7_75t_L g1533 ( 
.A(n_1427),
.B(n_1438),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1445),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1373),
.B(n_1385),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1421),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1406),
.B(n_1357),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1385),
.B(n_1417),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1417),
.B(n_1463),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1470),
.B(n_1448),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1445),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1448),
.B(n_1443),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1409),
.A2(n_1418),
.B(n_1358),
.C(n_1399),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1459),
.A2(n_1358),
.B1(n_1416),
.B2(n_1445),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1405),
.B(n_1357),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1358),
.A2(n_1416),
.B1(n_1357),
.B2(n_1436),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1397),
.A2(n_1390),
.B(n_1361),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1416),
.B(n_1413),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1397),
.A2(n_1361),
.B(n_1364),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1413),
.B(n_1455),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1367),
.A2(n_1399),
.B(n_1380),
.C(n_1455),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1380),
.A2(n_1455),
.B1(n_1412),
.B2(n_1410),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1370),
.B(n_1355),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1424),
.A2(n_1437),
.B1(n_1441),
.B2(n_1447),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1441),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1447),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1472),
.A2(n_745),
.B(n_1430),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1472),
.A2(n_1396),
.B(n_1393),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1359),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1371),
.B(n_1353),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1354),
.B(n_1348),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1351),
.B(n_1464),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1366),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1430),
.A2(n_1446),
.B(n_1333),
.C(n_1471),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1351),
.B(n_1464),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1371),
.B(n_1353),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1398),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1351),
.B(n_1464),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1430),
.A2(n_1322),
.B1(n_1446),
.B2(n_982),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1351),
.B(n_1464),
.Y(n_1571)
);

INVx3_ASAP7_75t_SL g1572 ( 
.A(n_1365),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1430),
.A2(n_1446),
.B(n_1322),
.C(n_1439),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1351),
.B(n_1464),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1351),
.B(n_1464),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1430),
.A2(n_745),
.B(n_1446),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1430),
.A2(n_745),
.B(n_1446),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1430),
.A2(n_745),
.B(n_1446),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1560),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1545),
.B(n_1537),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1538),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1555),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1489),
.A2(n_1485),
.B1(n_1570),
.B2(n_1492),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1484),
.B(n_1558),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1561),
.B(n_1567),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1522),
.B(n_1512),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1502),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1514),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1502),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1550),
.B(n_1548),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1512),
.B(n_1504),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1481),
.A2(n_1573),
.B(n_1565),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1561),
.B(n_1567),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1539),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1543),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1504),
.B(n_1487),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1506),
.B(n_1487),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1543),
.Y(n_1600)
);

INVxp67_ASAP7_75t_SL g1601 ( 
.A(n_1551),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1531),
.A2(n_1506),
.B(n_1494),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1570),
.A2(n_1492),
.B1(n_1491),
.B2(n_1490),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1501),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1535),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1505),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1546),
.B(n_1544),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1546),
.B(n_1544),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1530),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1552),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1490),
.B(n_1528),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1525),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1495),
.B(n_1491),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1495),
.B(n_1507),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1525),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1552),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1557),
.B(n_1556),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1553),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1563),
.B(n_1566),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1488),
.B(n_1499),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1554),
.A2(n_1549),
.B(n_1547),
.Y(n_1621)
);

AO21x2_ASAP7_75t_L g1622 ( 
.A1(n_1576),
.A2(n_1578),
.B(n_1577),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1498),
.B(n_1486),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1562),
.B(n_1511),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1499),
.A2(n_1488),
.B(n_1493),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1523),
.Y(n_1626)
);

BUFx12f_ASAP7_75t_L g1627 ( 
.A(n_1483),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1496),
.B(n_1500),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1547),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1564),
.B(n_1503),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1500),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1592),
.B(n_1575),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1582),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1582),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1582),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1585),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1587),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1594),
.A2(n_1526),
.B1(n_1529),
.B2(n_1524),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1593),
.B(n_1508),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1594),
.A2(n_1524),
.B1(n_1482),
.B2(n_1509),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1592),
.B(n_1598),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1510),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1593),
.B(n_1569),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1644)
);

INVx2_ASAP7_75t_R g1645 ( 
.A(n_1597),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1588),
.B(n_1571),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1618),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1583),
.A2(n_1482),
.B1(n_1497),
.B2(n_1509),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1590),
.Y(n_1649)
);

INVx4_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1580),
.B(n_1513),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1590),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1580),
.B(n_1534),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1589),
.B(n_1521),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1591),
.B(n_1516),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1586),
.B(n_1513),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1591),
.B(n_1541),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1643),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1642),
.A2(n_1628),
.B1(n_1625),
.B2(n_1622),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1638),
.A2(n_1603),
.B(n_1628),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1649),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

OAI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1655),
.A2(n_1620),
.B(n_1613),
.C(n_1631),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1648),
.A2(n_1584),
.B1(n_1631),
.B2(n_1613),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1635),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1650),
.A2(n_1625),
.B1(n_1584),
.B2(n_1620),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

OAI31xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1651),
.A2(n_1601),
.A3(n_1584),
.B(n_1619),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_SL g1669 ( 
.A(n_1655),
.B(n_1527),
.C(n_1614),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_SL g1670 ( 
.A(n_1655),
.B(n_1540),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1581),
.Y(n_1671)
);

NAND2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1632),
.B(n_1536),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1656),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1637),
.Y(n_1675)
);

AOI31xp33_ASAP7_75t_L g1676 ( 
.A1(n_1640),
.A2(n_1520),
.A3(n_1586),
.B(n_1595),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1646),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1633),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1623),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1650),
.B(n_1584),
.C(n_1614),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1634),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1641),
.B(n_1647),
.Y(n_1682)
);

AND4x1_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1542),
.C(n_1532),
.D(n_1595),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1634),
.Y(n_1684)
);

OAI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1643),
.A2(n_1611),
.B1(n_1607),
.B2(n_1608),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1650),
.B(n_1533),
.C(n_1615),
.D(n_1612),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1636),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1639),
.A2(n_1623),
.B1(n_1624),
.B2(n_1601),
.C(n_1611),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1651),
.B(n_1585),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1641),
.B(n_1581),
.Y(n_1690)
);

AOI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1644),
.A2(n_1626),
.B1(n_1579),
.B2(n_1600),
.C1(n_1610),
.C2(n_1616),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1647),
.B(n_1596),
.Y(n_1692)
);

OAI222xp33_ASAP7_75t_L g1693 ( 
.A1(n_1643),
.A2(n_1611),
.B1(n_1596),
.B2(n_1624),
.C1(n_1630),
.C2(n_1619),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1654),
.A2(n_1605),
.B1(n_1611),
.B2(n_1609),
.Y(n_1694)
);

OAI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1639),
.A2(n_1616),
.B1(n_1610),
.B2(n_1630),
.C(n_1572),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1649),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1647),
.B(n_1617),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1662),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1662),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1689),
.Y(n_1700)
);

OA21x2_ASAP7_75t_L g1701 ( 
.A1(n_1659),
.A2(n_1621),
.B(n_1629),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1696),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1695),
.Y(n_1704)
);

BUFx8_ASAP7_75t_L g1705 ( 
.A(n_1663),
.Y(n_1705)
);

BUFx8_ASAP7_75t_L g1706 ( 
.A(n_1687),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1665),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1667),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1661),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1682),
.B(n_1645),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1658),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1687),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1680),
.A2(n_1606),
.B(n_1604),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1674),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1682),
.B(n_1645),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1678),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1681),
.Y(n_1718)
);

INVx4_ASAP7_75t_SL g1719 ( 
.A(n_1689),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1681),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_L g1721 ( 
.A(n_1666),
.B(n_1639),
.C(n_1654),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1697),
.B(n_1632),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_L g1723 ( 
.A(n_1660),
.B(n_1602),
.C(n_1657),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1684),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1675),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1661),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1704),
.B(n_1691),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1698),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_L g1729 ( 
.A(n_1726),
.B(n_1669),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1679),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1719),
.B(n_1689),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1698),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1706),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1719),
.B(n_1689),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1712),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1711),
.B(n_1677),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1709),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1722),
.B(n_1632),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1726),
.B(n_1660),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1719),
.B(n_1700),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1699),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1671),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1699),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1711),
.B(n_1723),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1719),
.B(n_1700),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1719),
.B(n_1671),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1709),
.B(n_1627),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1700),
.B(n_1651),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1722),
.B(n_1690),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1722),
.B(n_1690),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1702),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1710),
.B(n_1697),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1702),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1707),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1721),
.A2(n_1668),
.B(n_1670),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1707),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1720),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1710),
.B(n_1692),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1710),
.B(n_1692),
.Y(n_1761)
);

NAND4xp25_ASAP7_75t_L g1762 ( 
.A(n_1723),
.B(n_1688),
.C(n_1686),
.D(n_1694),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1715),
.B(n_1651),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1726),
.Y(n_1764)
);

NOR2xp67_ASAP7_75t_SL g1765 ( 
.A(n_1721),
.B(n_1627),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1653),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1715),
.B(n_1653),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1712),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1726),
.B(n_1683),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1760),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1746),
.B(n_1738),
.Y(n_1773)
);

AND2x2_ASAP7_75t_SL g1774 ( 
.A(n_1727),
.B(n_1683),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1728),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1739),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1734),
.B(n_1712),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1760),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1761),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1728),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1733),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1746),
.B(n_1725),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1733),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1741),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1744),
.B(n_1748),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1738),
.B(n_1725),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1742),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1743),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1744),
.B(n_1748),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1741),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1734),
.Y(n_1791)
);

AOI32xp33_ASAP7_75t_L g1792 ( 
.A1(n_1729),
.A2(n_1672),
.A3(n_1726),
.B1(n_1685),
.B2(n_1664),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1769),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1757),
.A2(n_1676),
.B(n_1686),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1740),
.B(n_1646),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1749),
.B(n_1627),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1764),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1730),
.B(n_1705),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1745),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1753),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1770),
.B(n_1517),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1761),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1753),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1755),
.Y(n_1806)
);

NAND2x1_ASAP7_75t_SL g1807 ( 
.A(n_1742),
.B(n_1713),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1755),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1773),
.B(n_1737),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1793),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1775),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1776),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1791),
.B(n_1741),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1780),
.Y(n_1814)
);

INVx2_ASAP7_75t_SL g1815 ( 
.A(n_1777),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1773),
.B(n_1737),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1785),
.B(n_1732),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1777),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1777),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1781),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1772),
.B(n_1756),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1803),
.B(n_1741),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1785),
.B(n_1732),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1789),
.B(n_1747),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1798),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1789),
.B(n_1736),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1787),
.B(n_1736),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1783),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1772),
.B(n_1756),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1774),
.B(n_1731),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1787),
.B(n_1747),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1788),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1797),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1774),
.B(n_1735),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1798),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1807),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1825),
.B(n_1784),
.Y(n_1837)
);

AOI222xp33_ASAP7_75t_L g1838 ( 
.A1(n_1812),
.A2(n_1765),
.B1(n_1800),
.B2(n_1790),
.C1(n_1705),
.C2(n_1804),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1810),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1835),
.A2(n_1794),
.B1(n_1792),
.B2(n_1800),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1809),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1817),
.B(n_1778),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1815),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1815),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1818),
.B(n_1803),
.Y(n_1845)
);

OAI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1830),
.A2(n_1765),
.B1(n_1762),
.B2(n_1796),
.C(n_1804),
.Y(n_1846)
);

INVxp67_ASAP7_75t_SL g1847 ( 
.A(n_1809),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1834),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1822),
.A2(n_1796),
.B1(n_1779),
.B2(n_1778),
.C(n_1786),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1824),
.Y(n_1850)
);

NOR2x1_ASAP7_75t_L g1851 ( 
.A(n_1813),
.B(n_1819),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1824),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1816),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1824),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1836),
.A2(n_1568),
.B(n_1518),
.Y(n_1855)
);

NOR4xp25_ASAP7_75t_L g1856 ( 
.A(n_1811),
.B(n_1808),
.C(n_1806),
.D(n_1805),
.Y(n_1856)
);

OAI33xp33_ASAP7_75t_L g1857 ( 
.A1(n_1814),
.A2(n_1802),
.A3(n_1801),
.B1(n_1799),
.B2(n_1782),
.B3(n_1771),
.Y(n_1857)
);

NAND4xp75_ASAP7_75t_L g1858 ( 
.A(n_1817),
.B(n_1779),
.C(n_1701),
.D(n_1768),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1847),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1843),
.B(n_1823),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1841),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1851),
.B(n_1840),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1850),
.B(n_1823),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1852),
.B(n_1826),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1854),
.B(n_1826),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1845),
.B(n_1816),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1855),
.A2(n_1836),
.B(n_1831),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1853),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1852),
.Y(n_1869)
);

NOR2x1_ASAP7_75t_SL g1870 ( 
.A(n_1839),
.B(n_1827),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1842),
.B(n_1827),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1831),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1869),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1872),
.B(n_1844),
.Y(n_1874)
);

OAI21xp33_ASAP7_75t_L g1875 ( 
.A1(n_1862),
.A2(n_1837),
.B(n_1838),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1862),
.A2(n_1855),
.B(n_1846),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1867),
.A2(n_1848),
.B(n_1858),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1870),
.Y(n_1878)
);

NOR4xp25_ASAP7_75t_SL g1879 ( 
.A(n_1859),
.B(n_1849),
.C(n_1833),
.D(n_1828),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1866),
.B(n_1857),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1871),
.A2(n_1705),
.B1(n_1831),
.B2(n_1820),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1860),
.A2(n_1856),
.B(n_1832),
.Y(n_1882)
);

OAI21xp33_ASAP7_75t_L g1883 ( 
.A1(n_1863),
.A2(n_1865),
.B(n_1871),
.Y(n_1883)
);

OAI211xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1861),
.A2(n_1833),
.B(n_1828),
.C(n_1829),
.Y(n_1884)
);

OAI22xp33_ASAP7_75t_SL g1885 ( 
.A1(n_1878),
.A2(n_1868),
.B1(n_1821),
.B2(n_1829),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1873),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1880),
.A2(n_1864),
.B1(n_1872),
.B2(n_1705),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1875),
.B(n_1864),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1879),
.A2(n_1821),
.B(n_1782),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1874),
.Y(n_1890)
);

AOI211xp5_ASAP7_75t_L g1891 ( 
.A1(n_1877),
.A2(n_1786),
.B(n_1771),
.C(n_1768),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1883),
.B(n_1751),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1882),
.A2(n_1759),
.B(n_1758),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1887),
.B(n_1876),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1888),
.B(n_1892),
.Y(n_1895)
);

AND2x2_ASAP7_75t_SL g1896 ( 
.A(n_1890),
.B(n_1881),
.Y(n_1896)
);

AND3x1_ASAP7_75t_L g1897 ( 
.A(n_1891),
.B(n_1884),
.C(n_1759),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1885),
.A2(n_1750),
.B(n_1758),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1886),
.B(n_1795),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1889),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1893),
.B(n_1750),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1885),
.B(n_1750),
.Y(n_1902)
);

AOI222xp33_ASAP7_75t_L g1903 ( 
.A1(n_1900),
.A2(n_1705),
.B1(n_1706),
.B2(n_1693),
.C1(n_1763),
.C2(n_1754),
.Y(n_1903)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1904 ( 
.A1(n_1898),
.A2(n_1706),
.B(n_1714),
.C(n_1716),
.D(n_1717),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1901),
.B(n_1763),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1896),
.A2(n_1706),
.B1(n_1701),
.B2(n_1713),
.Y(n_1906)
);

NOR2xp67_ASAP7_75t_L g1907 ( 
.A(n_1902),
.B(n_1724),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1897),
.Y(n_1908)
);

AOI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1894),
.A2(n_1754),
.B1(n_1752),
.B2(n_1751),
.C(n_1766),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1908),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1905),
.A2(n_1895),
.B1(n_1899),
.B2(n_1906),
.C(n_1909),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1907),
.Y(n_1912)
);

NAND2xp33_ASAP7_75t_SL g1913 ( 
.A(n_1910),
.B(n_1904),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1913),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1914),
.Y(n_1915)
);

AOI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1914),
.A2(n_1912),
.B(n_1911),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1916),
.Y(n_1917)
);

OAI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1915),
.A2(n_1914),
.B(n_1903),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1917),
.B(n_1706),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1918),
.A2(n_1513),
.B1(n_1515),
.B2(n_1519),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1919),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1921),
.A2(n_1920),
.B1(n_1718),
.B2(n_1717),
.C(n_1708),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1922),
.B(n_1766),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_SL g1924 ( 
.A1(n_1923),
.A2(n_1541),
.B(n_1713),
.Y(n_1924)
);

OAI22x1_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1519),
.B1(n_1515),
.B2(n_1513),
.Y(n_1925)
);

AOI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1767),
.B(n_1752),
.C(n_1652),
.Y(n_1926)
);


endmodule