module fake_jpeg_3693_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_55),
.B1(n_40),
.B2(n_51),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_54),
.B1(n_56),
.B2(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_54),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_40),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_90),
.B1(n_47),
.B2(n_44),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_21),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_43),
.B1(n_47),
.B2(n_44),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_107),
.B1(n_92),
.B2(n_105),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_76),
.B1(n_82),
.B2(n_18),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_110),
.Y(n_135)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_116),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_14),
.B(n_38),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_2),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_39),
.C(n_33),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_26),
.C(n_25),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_3),
.B(n_4),
.Y(n_122)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_4),
.B(n_5),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_3),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_24),
.A3(n_23),
.B1(n_22),
.B2(n_9),
.C(n_10),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_113),
.A3(n_119),
.B1(n_122),
.B2(n_120),
.C1(n_11),
.C2(n_12),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.C(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_143),
.B1(n_128),
.B2(n_126),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_125),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_135),
.C(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_145),
.C(n_144),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_127),
.B(n_128),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_153),
.C(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_133),
.B1(n_139),
.B2(n_127),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_156),
.C(n_131),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_130),
.C(n_155),
.Y(n_159)
);

AO21x1_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_153),
.B(n_143),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_6),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_13),
.C(n_8),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_7),
.Y(n_164)
);


endmodule