module real_jpeg_22468_n_16 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_41),
.B1(n_49),
.B2(n_54),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_24),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_24),
.B1(n_44),
.B2(n_45),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_2),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_2),
.A2(n_14),
.B(n_45),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_41),
.B1(n_49),
.B2(n_117),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_92),
.B1(n_174),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_2),
.B(n_74),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_29),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_29),
.B(n_202),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_114),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_41),
.B1(n_49),
.B2(n_114),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_114),
.Y(n_252)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_5),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_112),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_112),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_5),
.A2(n_41),
.B1(n_49),
.B2(n_112),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_32),
.B1(n_41),
.B2(n_49),
.Y(n_101)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_7),
.A2(n_126),
.B(n_148),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_56),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_9),
.A2(n_41),
.B1(n_49),
.B2(n_56),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_290)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_11),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_41),
.B1(n_49),
.B2(n_119),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_119),
.Y(n_174)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_41),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_336),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_80),
.B(n_334),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_20),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_21),
.A2(n_52),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_22),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_336)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_27),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_27),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_23),
.B(n_117),
.CON(n_116),
.SN(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_31),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_33),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_27),
.B(n_29),
.Y(n_123)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_28),
.A2(n_34),
.B1(n_116),
.B2(n_123),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_28),
.A2(n_41),
.A3(n_64),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_29),
.A2(n_62),
.B(n_63),
.C(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_63),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_30),
.A2(n_53),
.B(n_57),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_33),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_36),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_72),
.C(n_76),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_37),
.A2(n_38),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_50),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_39),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_39),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_39),
.A2(n_58),
.B1(n_59),
.B2(n_310),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_47),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_40),
.A2(n_47),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_40),
.A2(n_43),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_40),
.A2(n_43),
.B1(n_170),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_40),
.A2(n_43),
.B1(n_191),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_40),
.A2(n_209),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_40),
.A2(n_43),
.B1(n_99),
.B2(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_40),
.A2(n_107),
.B(n_244),
.Y(n_278)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_43),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_43),
.B(n_117),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_44),
.B(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_93),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_46),
.A2(n_49),
.B(n_117),
.C(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_48),
.B(n_108),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g203 ( 
.A(n_49),
.B(n_63),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_50),
.A2(n_51),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_52),
.A2(n_57),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_52),
.A2(n_57),
.B1(n_132),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_52),
.A2(n_79),
.B(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_57),
.B(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_67),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_68),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_62),
.A2(n_68),
.B1(n_111),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_62),
.A2(n_68),
.B1(n_144),
.B2(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_62),
.B(n_71),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_62),
.A2(n_66),
.B(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_62),
.A2(n_68),
.B1(n_269),
.B2(n_290),
.Y(n_289)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_74),
.B(n_75),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_67),
.A2(n_75),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_67),
.A2(n_255),
.B(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_76),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_327),
.B(n_333),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_303),
.A3(n_322),
.B1(n_325),
.B2(n_326),
.C(n_339),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_282),
.B(n_302),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_260),
.B(n_281),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_149),
.B(n_234),
.C(n_259),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_137),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_86),
.B(n_137),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_120),
.B2(n_136),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_104),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_89),
.B(n_104),
.C(n_136),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_98),
.B2(n_103),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_90),
.B(n_103),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_94),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_92),
.A2(n_127),
.B1(n_159),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_92),
.A2(n_162),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_92),
.A2(n_93),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_96),
.A2(n_157),
.B(n_194),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_100),
.B(n_225),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_127),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_121),
.B(n_129),
.C(n_134),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_138),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_143),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_233),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_227),
.B(n_232),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_214),
.B(n_226),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_196),
.B(n_213),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_183),
.B(n_195),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_171),
.B(n_182),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_176),
.B(n_181),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_185),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_194),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_198),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_204),
.B1(n_211),
.B2(n_212),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_199),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_216),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_223),
.C(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_257),
.B2(n_258),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_246),
.C(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_256),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_254),
.C(n_256),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_280),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_274),
.C(n_280),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_270),
.C(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_276),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_293),
.B(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_278),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_284),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_300),
.B2(n_301),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_292),
.C(n_301),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B(n_291),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_290),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_305),
.C(n_314),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_291),
.B(n_305),
.CI(n_314),
.CON(n_324),
.SN(n_324)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_297),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_315),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_315),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_307),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_320),
.C(n_321),
.Y(n_328)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_330),
.Y(n_332)
);


endmodule