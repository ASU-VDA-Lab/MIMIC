module real_jpeg_6738_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_0),
.A2(n_43),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_0),
.A2(n_259),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_0),
.A2(n_126),
.B1(n_259),
.B2(n_351),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_0),
.A2(n_105),
.B1(n_259),
.B2(n_444),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_1),
.A2(n_96),
.B1(n_180),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_1),
.B(n_290),
.C(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_1),
.B(n_92),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_1),
.B(n_162),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_1),
.B(n_139),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_1),
.B(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_41),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_2),
.A2(n_127),
.B1(n_194),
.B2(n_286),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_2),
.A2(n_135),
.B1(n_163),
.B2(n_194),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_2),
.A2(n_194),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_3),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_3),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_3),
.Y(n_242)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_3),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_4),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_54),
.B1(n_56),
.B2(n_61),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_61),
.B1(n_90),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_5),
.A2(n_61),
.B1(n_120),
.B2(n_184),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_5),
.A2(n_61),
.B1(n_233),
.B2(n_237),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_6),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_7),
.A2(n_180),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_7),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_7),
.A2(n_310),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_7),
.A2(n_310),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_7),
.A2(n_40),
.B1(n_310),
.B2(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_8),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_40),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_9),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_9),
.A2(n_77),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_9),
.A2(n_77),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_9),
.A2(n_77),
.B1(n_297),
.B2(n_318),
.Y(n_429)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_42),
.B1(n_71),
.B2(n_74),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_11),
.A2(n_74),
.B1(n_106),
.B2(n_203),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_11),
.A2(n_74),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_11),
.A2(n_74),
.B1(n_168),
.B2(n_297),
.Y(n_406)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_12),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_42),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_13),
.A2(n_189),
.B1(n_251),
.B2(n_255),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_13),
.A2(n_189),
.B1(n_237),
.B2(n_373),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_13),
.A2(n_189),
.B1(n_448),
.B2(n_451),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_14),
.Y(n_171)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_14),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_15),
.Y(n_533)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_18),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_18),
.A2(n_50),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_18),
.A2(n_50),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_18),
.A2(n_50),
.B1(n_168),
.B2(n_172),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_528),
.B(n_531),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_64),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_51),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_46),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_24),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_24),
.B(n_193),
.Y(n_262)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_27),
.B(n_357),
.Y(n_420)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_30),
.Y(n_367)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_31),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_32),
.Y(n_358)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_34),
.Y(n_205)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_34),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_36),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_36),
.A2(n_436),
.B(n_440),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_51)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_49),
.B(n_283),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_51),
.B(n_66),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_62),
.B1(n_70),
.B2(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_52),
.A2(n_62),
.B1(n_70),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_52),
.A2(n_258),
.B(n_262),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_52),
.A2(n_62),
.B1(n_258),
.B2(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_55),
.Y(n_196)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_55),
.Y(n_473)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_59),
.Y(n_416)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_60),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_62),
.B(n_283),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_62),
.A2(n_192),
.B(n_471),
.Y(n_488)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_150),
.B(n_527),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_146),
.C(n_147),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_67),
.A2(n_68),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_78),
.C(n_114),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_69),
.B(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_78),
.A2(n_114),
.B1(n_115),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_78),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_79),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_79),
.A2(n_104),
.B1(n_107),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_79),
.A2(n_107),
.B1(n_202),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_79),
.A2(n_107),
.B1(n_398),
.B2(n_443),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_92),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_86),
.B2(n_90),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_85),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_85),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_85),
.Y(n_256)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_90),
.Y(n_400)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_92),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_92),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_92),
.A2(n_148),
.B1(n_201),
.B2(n_206),
.Y(n_200)
);

AOI22x1_ASAP7_75t_L g474 ( 
.A1(n_92),
.A2(n_148),
.B1(n_402),
.B2(n_475),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_95),
.Y(n_381)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_98),
.Y(n_248)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_98),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_98),
.Y(n_384)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_101),
.Y(n_453)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_107),
.B(n_365),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_107),
.A2(n_398),
.B(n_401),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_110),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_111),
.Y(n_399)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_114),
.A2(n_115),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_114),
.B(n_213),
.C(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_138),
.B(n_140),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_116),
.A2(n_282),
.B(n_284),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_116),
.A2(n_138),
.B1(n_307),
.B2(n_350),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_116),
.A2(n_284),
.B(n_350),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_116),
.A2(n_138),
.B1(n_447),
.B2(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_117),
.A2(n_139),
.B1(n_175),
.B2(n_183),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_117),
.A2(n_139),
.B1(n_183),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_117),
.A2(n_139),
.B1(n_175),
.B2(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_117),
.B(n_285),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_128),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_124),
.B2(n_126),
.Y(n_118)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_120),
.B(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_123),
.Y(n_290)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_128),
.A2(n_307),
.B(n_311),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_135),
.B2(n_137),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_134),
.Y(n_373)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_138),
.A2(n_311),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_139),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_146),
.B(n_147),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_148),
.A2(n_355),
.B(n_364),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_148),
.B(n_402),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_148),
.A2(n_364),
.B(n_491),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_521),
.B(n_526),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_274),
.B(n_518),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_263),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_220),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_154),
.B(n_220),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_154),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_197),
.CI(n_211),
.CON(n_154),
.SN(n_154)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_155),
.B(n_197),
.C(n_211),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B(n_186),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_174),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_157),
.A2(n_186),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_157),
.A2(n_174),
.B1(n_225),
.B2(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_166),
.B(n_167),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_158),
.A2(n_167),
.B1(n_232),
.B2(n_240),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_158),
.A2(n_295),
.B(n_300),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_158),
.A2(n_283),
.B(n_300),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_158),
.A2(n_424),
.B1(n_425),
.B2(n_428),
.Y(n_423)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_159),
.B(n_303),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_159),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_159),
.A2(n_161),
.B1(n_372),
.B2(n_406),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_159),
.A2(n_301),
.B1(n_429),
.B2(n_468),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_162),
.Y(n_302)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_170),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_171),
.Y(n_328)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_174),
.Y(n_462)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g374 ( 
.A1(n_177),
.A2(n_360),
.A3(n_375),
.B1(n_379),
.B2(n_382),
.Y(n_374)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_178),
.Y(n_309)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g415 ( 
.A1(n_203),
.A2(n_416),
.A3(n_417),
.B1(n_420),
.B2(n_421),
.Y(n_415)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_219),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_212),
.A2(n_213),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_212),
.B(n_265),
.C(n_269),
.Y(n_525)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.C(n_229),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_226),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_229),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_249),
.C(n_257),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_230),
.B(n_460),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_231),
.B(n_243),
.Y(n_485)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_232),
.Y(n_468)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_240),
.A2(n_323),
.B(n_329),
.Y(n_322)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_244),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_248),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_249),
.B(n_257),
.Y(n_460)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_250),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_256),
.Y(n_378)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_262),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_263),
.A2(n_519),
.B(n_520),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_273),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_264),
.B(n_273),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI311xp33_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_456),
.A3(n_494),
.B1(n_512),
.C1(n_513),
.Y(n_274)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_409),
.B(n_455),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_389),
.B(n_408),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_344),
.B(n_388),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_314),
.B(n_343),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_293),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_280),
.B(n_293),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_287),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_281),
.A2(n_287),
.B1(n_288),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_SL g355 ( 
.A1(n_283),
.A2(n_356),
.B(n_359),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_SL g436 ( 
.A1(n_283),
.A2(n_421),
.B(n_437),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_304),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_294),
.B(n_305),
.C(n_313),
.Y(n_345)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_302),
.A2(n_329),
.B(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_312),
.B2(n_313),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_332),
.B(n_342),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_321),
.B(n_331),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_330),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_330),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_340),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_340),
.Y(n_342)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_345),
.B(n_346),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_369),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_353),
.B2(n_354),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_353),
.C(n_369),
.Y(n_390)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_374),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_381),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_385),
.Y(n_382)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_390),
.B(n_391),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_396),
.B2(n_407),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_395),
.C(n_407),
.Y(n_410)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_396),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_403),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_404),
.C(n_405),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_410),
.B(n_411),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_433),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_412)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_422),
.B2(n_423),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_415),
.B(n_422),
.Y(n_489)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_430),
.B(n_431),
.C(n_433),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_441),
.B2(n_454),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_434),
.B(n_442),
.C(n_446),
.Y(n_503)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_446),
.Y(n_441)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_443),
.Y(n_491)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_479),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_SL g513 ( 
.A1(n_457),
.A2(n_479),
.B(n_514),
.C(n_517),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_476),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_458),
.B(n_476),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.C(n_463),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_461),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_469),
.C(n_474),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_467),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_469),
.A2(n_470),
.B1(n_474),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_474),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_492),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_492),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_485),
.C(n_486),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_481),
.A2(n_482),
.B1(n_485),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_485),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.C(n_490),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_487),
.A2(n_488),
.B1(n_490),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_507),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_515),
.B(n_516),
.Y(n_514)
);

NOR2x1_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_504),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_504),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_501),
.C(n_503),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_510),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_502),
.B1(n_503),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_503),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_509),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_525),
.Y(n_526)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

BUFx4f_ASAP7_75t_SL g532 ( 
.A(n_529),
.Y(n_532)
);

INVx13_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);


endmodule