module real_jpeg_25544_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_1),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_88),
.B1(n_112),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_88),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_3),
.A2(n_72),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_123),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_123),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_123),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_70),
.B1(n_73),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_79),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_79),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_79),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_77),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_8),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_41),
.B1(n_65),
.B2(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_51),
.B1(n_65),
.B2(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_11),
.B(n_125),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_113),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_11),
.A2(n_28),
.B(n_44),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_11),
.B(n_90),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_11),
.A2(n_25),
.B1(n_130),
.B2(n_225),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_65),
.B(n_239),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_15),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_151),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_150),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_127),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_20),
.B(n_127),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.C(n_104),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_21),
.A2(n_22),
.B1(n_93),
.B2(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_57),
.B1(n_58),
.B2(n_92),
.Y(n_22)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_24),
.B(n_42),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_25),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_97),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_25),
.A2(n_100),
.B1(n_216),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_25),
.A2(n_35),
.B(n_131),
.Y(n_248)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_26),
.B(n_40),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_26),
.A2(n_33),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_26),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_28),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_27),
.B(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_39),
.A2(n_96),
.B(n_118),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g218 ( 
.A(n_39),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B(n_52),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_43),
.A2(n_47),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_43),
.B(n_54),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_43),
.A2(n_102),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_43),
.B(n_113),
.Y(n_223)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_46),
.A2(n_49),
.B(n_113),
.C(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_49),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_48),
.B(n_85),
.Y(n_247)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_49),
.A2(n_65),
.A3(n_84),
.B1(n_240),
.B2(n_247),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_55),
.A2(n_135),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_55),
.A2(n_199),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_55),
.A2(n_207),
.B1(n_208),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_80),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_59),
.B(n_80),
.C(n_92),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_74),
.B2(n_78),
.Y(n_59)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_60),
.A2(n_78),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_69),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_61),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_63),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_66),
.A3(n_72),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_65),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_66),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_66),
.B(n_113),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_73),
.A2(n_111),
.B(n_113),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_74),
.Y(n_126)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_89),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_81),
.A2(n_83),
.B1(n_183),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_82),
.B(n_91),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_82),
.A2(n_90),
.B1(n_107),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_82),
.A2(n_90),
.B1(n_165),
.B2(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_87),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_103),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_102),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_104),
.A2(n_105),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_120),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_120),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_113),
.B(n_130),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_143),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_127),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_137),
.CI(n_149),
.CON(n_127),
.SN(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_136),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_129),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_148),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_188),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_170),
.B(n_187),
.Y(n_153)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_154),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_167),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_167),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_166),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_157),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_159),
.B(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_161),
.B(n_207),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_171),
.B(n_174),
.Y(n_275)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_175),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_177),
.Y(n_272)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.C(n_185),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_181),
.B(n_257),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_274),
.C(n_275),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_268),
.B(n_273),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_252),
.B(n_267),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_233),
.B(n_251),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_212),
.B(n_232),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_202),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_194),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_209),
.C(n_210),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_221),
.B(n_231),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_219),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_226),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_245),
.B1(n_249),
.B2(n_250),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_244),
.C(n_249),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_248),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_262),
.C(n_265),
.Y(n_269)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);


endmodule