module fake_jpeg_9145_n_175 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_38),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_44),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_16),
.B1(n_22),
.B2(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_34),
.Y(n_67)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_67),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_20),
.B1(n_24),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_72),
.B1(n_28),
.B2(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_27),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_63),
.B1(n_64),
.B2(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_27),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_35),
.B1(n_38),
.B2(n_14),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_45),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_87),
.C(n_72),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_1),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_90),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_72),
.B(n_62),
.C(n_51),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_35),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_84),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_74),
.B1(n_77),
.B2(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_85),
.Y(n_112)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_61),
.C(n_28),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_80),
.C(n_82),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_25),
.C(n_9),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_115),
.C(n_100),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_87),
.B(n_82),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_116),
.B(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_117),
.B1(n_91),
.B2(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_103),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_86),
.C(n_81),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_86),
.B1(n_23),
.B2(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_76),
.B1(n_23),
.B2(n_66),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_76),
.B(n_66),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_132),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_124),
.B(n_130),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_134),
.C(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_129),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_96),
.A3(n_91),
.B1(n_101),
.B2(n_11),
.C1(n_12),
.C2(n_8),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_111),
.B1(n_116),
.B2(n_93),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_122),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_145),
.B1(n_105),
.B2(n_4),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_115),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_2),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_114),
.C(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_93),
.C(n_102),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_105),
.B(n_3),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_152),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_8),
.C(n_9),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_5),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_11),
.Y(n_154)
);

AOI31xp67_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_2),
.A3(n_4),
.B(n_5),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_143),
.B1(n_141),
.B2(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_6),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_157),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_161),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_161),
.C(n_162),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.C(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_6),
.Y(n_175)
);


endmodule