module fake_jpeg_3619_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_62),
.Y(n_69)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_70),
.B1(n_64),
.B2(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_56),
.B1(n_61),
.B2(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_50),
.B1(n_63),
.B2(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_60),
.Y(n_91)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_63),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_52),
.B1(n_48),
.B2(n_49),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_92),
.B1(n_98),
.B2(n_99),
.Y(n_107)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_76),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_8),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_96),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_117)
);

FAx1_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_50),
.CI(n_2),
.CON(n_96),
.SN(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_50),
.B1(n_57),
.B2(n_5),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_83),
.B1(n_80),
.B2(n_23),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_4),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_7),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_117),
.B1(n_90),
.B2(n_13),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_11),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_124),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_15),
.B1(n_24),
.B2(n_25),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_13),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_29),
.B(n_41),
.C(n_17),
.D(n_20),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_136),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_31),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_138),
.C(n_34),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_139),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_27),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_14),
.B(n_15),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_117),
.B1(n_115),
.B2(n_14),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_123),
.B1(n_134),
.B2(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_45),
.B1(n_21),
.B2(n_22),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_149),
.B(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_145),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_39),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_32),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_138),
.B(n_121),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_161),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_159),
.B1(n_155),
.B2(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_160),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_36),
.A3(n_37),
.B1(n_154),
.B2(n_146),
.C1(n_141),
.C2(n_148),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_147),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_165),
.B(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_153),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_157),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_168),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_163),
.B(n_169),
.C(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_144),
.Y(n_176)
);


endmodule