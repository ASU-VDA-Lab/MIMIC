module fake_netlist_5_1435_n_120 (n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_120);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_120;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_29;
wire n_79;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_76;
wire n_36;
wire n_87;
wire n_77;
wire n_64;
wire n_106;
wire n_102;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_104;
wire n_41;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_6),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_1),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_11),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

CKINVDCx11_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_32),
.Y(n_66)
);

XNOR2x2_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_51),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_33),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_45),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_40),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_48),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

OAI21x1_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_70),
.B(n_75),
.Y(n_80)
);

NOR4xp25_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_31),
.C(n_29),
.D(n_43),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_35),
.B(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_61),
.Y(n_84)
);

AOI21x1_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_59),
.B(n_61),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_31),
.B1(n_62),
.B2(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_64),
.B1(n_59),
.B2(n_36),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_R g89 ( 
.A(n_83),
.B(n_63),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_2),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_86),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_87),
.B1(n_82),
.B2(n_81),
.C(n_84),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_93),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_90),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_91),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_98),
.B1(n_87),
.B2(n_81),
.C(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_80),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_80),
.B(n_92),
.C(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_102),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

OAI221xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_103),
.B1(n_105),
.B2(n_85),
.C(n_50),
.Y(n_109)
);

AOI211xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_41),
.B(n_64),
.C(n_92),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_64),
.B(n_65),
.C(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_111),
.B(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_109),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_117)
);

AOI31xp33_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_65),
.A3(n_56),
.B(n_54),
.Y(n_118)
);

OAI221xp5_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_115),
.B1(n_10),
.B2(n_15),
.C(n_19),
.Y(n_119)
);

OAI221xp5_ASAP7_75t_R g120 ( 
.A1(n_119),
.A2(n_118),
.B1(n_115),
.B2(n_26),
.C(n_21),
.Y(n_120)
);


endmodule