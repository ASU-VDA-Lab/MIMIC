module fake_jpeg_2333_n_124 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_13),
.C(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_35),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_61),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_49),
.B1(n_43),
.B2(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_69),
.B1(n_44),
.B2(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_0),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_53),
.B(n_51),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_59),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_47),
.C(n_42),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_38),
.B1(n_47),
.B2(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_15),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_59),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_79),
.Y(n_87)
);

AO21x2_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_59),
.B(n_58),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_81),
.C(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_12),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_1),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_20),
.B1(n_29),
.B2(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_1),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_94),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_93),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_17),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_95),
.C(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_11),
.B(n_32),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_103),
.B(n_9),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_7),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_9),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_111),
.C(n_112),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_96),
.B1(n_86),
.B2(n_10),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_R g115 ( 
.A(n_113),
.B(n_102),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_115),
.A2(n_112),
.B(n_110),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_107),
.C(n_99),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.C(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_116),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_98),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_10),
.Y(n_124)
);


endmodule