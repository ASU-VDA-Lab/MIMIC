module fake_ariane_2645_n_678 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_678);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_678;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_663;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_672;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_129;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_136;
wire n_334;
wire n_192;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_127;
wire n_531;
wire n_675;

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_66),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_44),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_35),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_59),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_22),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx8_ASAP7_75t_SL g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_65),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_29),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_70),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_31),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_33),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_30),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_42),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_32),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_16),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_10),
.B(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_6),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_61),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_27),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_26),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_28),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_103),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_50),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_0),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

OAI22x1_ASAP7_75t_R g191 ( 
.A1(n_179),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_1),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_2),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_138),
.B(n_4),
.Y(n_200)
);

BUFx8_ASAP7_75t_SL g201 ( 
.A(n_179),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_5),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_5),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_134),
.B(n_6),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_134),
.B(n_7),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_147),
.A2(n_7),
.B(n_8),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_8),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_156),
.B(n_9),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_127),
.B(n_9),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_10),
.B(n_11),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_166),
.A2(n_11),
.B(n_12),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_127),
.C(n_130),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

BUFx6f_ASAP7_75t_SL g235 ( 
.A(n_200),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_136),
.C(n_130),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

AO21x2_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_185),
.B(n_183),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_167),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_211),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_211),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_168),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_171),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_208),
.B(n_136),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_173),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_176),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_188),
.A2(n_180),
.B(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

NOR2x1p5_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_174),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_208),
.B(n_174),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_129),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_164),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_209),
.B(n_13),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_131),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_153),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_189),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_189),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_189),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_196),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_196),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_210),
.B1(n_213),
.B2(n_208),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_243),
.B(n_196),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_200),
.B1(n_205),
.B2(n_213),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_207),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_254),
.A2(n_210),
.B1(n_213),
.B2(n_149),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_212),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_212),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_222),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_219),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_210),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_215),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_229),
.B1(n_214),
.B2(n_226),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_235),
.A2(n_149),
.B1(n_218),
.B2(n_217),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_215),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_236),
.B(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_265),
.B(n_182),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_215),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_276),
.B(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_222),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_139),
.B1(n_182),
.B2(n_225),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_216),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_263),
.B(n_216),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_255),
.B(n_224),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_274),
.B(n_224),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_225),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_R g319 ( 
.A(n_266),
.B(n_133),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_232),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_229),
.B(n_226),
.C(n_214),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_262),
.A2(n_229),
.B1(n_226),
.B2(n_214),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_221),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g326 ( 
.A(n_270),
.B(n_214),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_268),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_234),
.A2(n_229),
.B(n_226),
.C(n_228),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_216),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_148),
.B1(n_150),
.B2(n_155),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_238),
.B(n_221),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_244),
.A2(n_221),
.B1(n_228),
.B2(n_204),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_216),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_304),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_244),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_282),
.A2(n_204),
.B(n_202),
.C(n_258),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_251),
.B(n_248),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_293),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_246),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_251),
.B(n_248),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_290),
.A2(n_157),
.B1(n_158),
.B2(n_240),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_292),
.B(n_202),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_281),
.A2(n_247),
.B(n_246),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_286),
.B(n_285),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_247),
.B(n_240),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_204),
.B(n_240),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_302),
.Y(n_348)
);

O2A1O1Ixp33_ASAP7_75t_SL g349 ( 
.A1(n_299),
.A2(n_191),
.B(n_14),
.C(n_15),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_201),
.C(n_145),
.Y(n_350)
);

AOI21x1_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_204),
.B(n_240),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_295),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_303),
.A2(n_204),
.B(n_69),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_307),
.A2(n_64),
.B(n_124),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_13),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_323),
.A2(n_63),
.B(n_123),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_14),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_325),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_71),
.B(n_122),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_288),
.B(n_15),
.Y(n_361)
);

NOR3xp33_ASAP7_75t_L g362 ( 
.A(n_296),
.B(n_327),
.C(n_284),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_288),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_298),
.B(n_201),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_330),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g366 ( 
.A1(n_314),
.A2(n_24),
.B(n_25),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_279),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_300),
.A2(n_34),
.B(n_36),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_SL g370 ( 
.A(n_311),
.B(n_37),
.C(n_38),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_280),
.A2(n_39),
.B(n_40),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_287),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_301),
.A2(n_41),
.B(n_43),
.Y(n_374)
);

OA22x2_ASAP7_75t_L g375 ( 
.A1(n_316),
.A2(n_305),
.B1(n_309),
.B2(n_313),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_45),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_320),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_315),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_318),
.B(n_120),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_322),
.A2(n_46),
.B(n_47),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_48),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_321),
.B(n_119),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_49),
.C(n_51),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_301),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_321),
.A2(n_57),
.B(n_58),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_118),
.Y(n_387)
);

NOR2x1_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_60),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_282),
.B(n_77),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_79),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_84),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_348),
.A2(n_85),
.B(n_87),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_347),
.A2(n_90),
.B(n_91),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_390),
.A2(n_96),
.B(n_97),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_334),
.B(n_101),
.Y(n_397)
);

NAND2x1p5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_102),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_345),
.B(n_358),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_364),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_374),
.A2(n_105),
.B(n_107),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_344),
.A2(n_108),
.B(n_110),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_111),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_373),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_113),
.C(n_114),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_336),
.A2(n_116),
.B(n_335),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_357),
.B(n_361),
.Y(n_409)
);

O2A1O1Ixp5_ASAP7_75t_L g410 ( 
.A1(n_376),
.A2(n_380),
.B(n_382),
.C(n_339),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_356),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_377),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_372),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_346),
.A2(n_369),
.B(n_354),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_385),
.A2(n_363),
.B(n_340),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_387),
.A2(n_365),
.B1(n_383),
.B2(n_384),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_360),
.A2(n_355),
.B(n_371),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_381),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_349),
.A2(n_345),
.B(n_347),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_345),
.A2(n_347),
.B(n_344),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_345),
.B(n_335),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_337),
.A2(n_341),
.B(n_351),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_390),
.B(n_338),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_390),
.B(n_338),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_411),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_410),
.A2(n_426),
.B(n_409),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_411),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_428),
.A2(n_416),
.B(n_422),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

AOI31xp67_ASAP7_75t_L g438 ( 
.A1(n_423),
.A2(n_409),
.A3(n_431),
.B(n_430),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_431),
.B(n_430),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_406),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_400),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

NAND2x1p5_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_429),
.Y(n_443)
);

OAI21x1_ASAP7_75t_SL g444 ( 
.A1(n_394),
.A2(n_417),
.B(n_420),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_408),
.B(n_404),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_432),
.Y(n_447)
);

O2A1O1Ixp5_ASAP7_75t_L g448 ( 
.A1(n_410),
.A2(n_421),
.B(n_424),
.C(n_392),
.Y(n_448)
);

AOI222xp33_ASAP7_75t_L g449 ( 
.A1(n_393),
.A2(n_405),
.B1(n_391),
.B2(n_415),
.C1(n_413),
.C2(n_412),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_396),
.B(n_407),
.Y(n_450)
);

NAND2x1_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_419),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_424),
.A2(n_418),
.B(n_429),
.C(n_395),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_393),
.Y(n_454)
);

OAI221xp5_ASAP7_75t_L g455 ( 
.A1(n_395),
.A2(n_348),
.B1(n_290),
.B2(n_292),
.C(n_197),
.Y(n_455)
);

AO21x2_ASAP7_75t_L g456 ( 
.A1(n_398),
.A2(n_409),
.B(n_427),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_409),
.A2(n_425),
.B(n_347),
.Y(n_457)
);

AO21x2_ASAP7_75t_L g458 ( 
.A1(n_409),
.A2(n_427),
.B(n_423),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_353),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_409),
.A2(n_338),
.B(n_431),
.C(n_430),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_410),
.A2(n_426),
.B(n_409),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

BUFx4f_ASAP7_75t_L g463 ( 
.A(n_393),
.Y(n_463)
);

INVx3_ASAP7_75t_SL g464 ( 
.A(n_406),
.Y(n_464)
);

AO31x2_ASAP7_75t_L g465 ( 
.A1(n_420),
.A2(n_427),
.A3(n_401),
.B(n_423),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_397),
.A2(n_288),
.B1(n_338),
.B2(n_361),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_463),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

CKINVDCx11_ASAP7_75t_R g470 ( 
.A(n_464),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_441),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_450),
.B(n_444),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_454),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_433),
.B(n_435),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_436),
.A2(n_453),
.B(n_448),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_433),
.B(n_435),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_460),
.Y(n_484)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_453),
.A2(n_448),
.B(n_446),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

BUFx12f_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_463),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_464),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_450),
.A2(n_457),
.B(n_461),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_465),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_456),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_437),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_456),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_457),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_468),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_492),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_468),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_472),
.B(n_434),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_472),
.B(n_434),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_477),
.B(n_465),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_477),
.B(n_482),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_437),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_494),
.B(n_465),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_477),
.B(n_465),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_458),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_486),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_489),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_466),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_476),
.B(n_455),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_499),
.A2(n_455),
.B1(n_487),
.B2(n_476),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_487),
.A2(n_476),
.B1(n_496),
.B2(n_481),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_483),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_474),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_495),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_495),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_515),
.B(n_490),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_507),
.B(n_491),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_531),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_527),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_503),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_491),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_521),
.B(n_475),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_511),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_513),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_519),
.B(n_471),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_527),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_532),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_532),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_518),
.B(n_485),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_518),
.B(n_485),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_512),
.B(n_471),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_485),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_505),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_525),
.B(n_474),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_521),
.B(n_478),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_517),
.B(n_526),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_526),
.B(n_478),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_525),
.B(n_478),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_522),
.B(n_535),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_542),
.B(n_516),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_553),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_516),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_553),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_522),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_504),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_545),
.B(n_508),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_565),
.B(n_524),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_541),
.B(n_520),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_550),
.B(n_520),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_554),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_541),
.B(n_520),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_506),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_554),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_544),
.B(n_528),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_548),
.B(n_506),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_546),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_549),
.B(n_528),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_555),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_533),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_543),
.B(n_528),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_568),
.B(n_505),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_556),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_566),
.B(n_561),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_556),
.B(n_533),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_557),
.B(n_533),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_557),
.B(n_470),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

OAI211xp5_ASAP7_75t_L g598 ( 
.A1(n_552),
.A2(n_529),
.B(n_530),
.C(n_467),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_549),
.B(n_558),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_574),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_566),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_570),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_596),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_572),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_559),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_579),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_537),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_575),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_586),
.B(n_559),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_586),
.A2(n_539),
.B1(n_537),
.B2(n_502),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_567),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_539),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_573),
.B(n_563),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_593),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_595),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_597),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_599),
.A2(n_590),
.B(n_586),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_604),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_611),
.A2(n_590),
.B(n_563),
.C(n_589),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_603),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_609),
.B(n_577),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_604),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_617),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_581),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_608),
.B(n_600),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_616),
.B(n_467),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_608),
.A2(n_609),
.B1(n_567),
.B2(n_583),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_619),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_621),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_623),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_618),
.Y(n_632)
);

OAI31xp33_ASAP7_75t_L g633 ( 
.A1(n_620),
.A2(n_609),
.A3(n_614),
.B(n_615),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_622),
.Y(n_634)
);

OAI222xp33_ASAP7_75t_L g635 ( 
.A1(n_632),
.A2(n_628),
.B1(n_626),
.B2(n_625),
.C1(n_627),
.C2(n_624),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_634),
.A2(n_630),
.B1(n_622),
.B2(n_601),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_629),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_634),
.B(n_613),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_631),
.A2(n_612),
.B1(n_578),
.B2(n_591),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_629),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_637),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_640),
.B(n_633),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_638),
.B(n_636),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_639),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_635),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_SL g646 ( 
.A(n_642),
.B(n_488),
.C(n_576),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_645),
.B(n_602),
.C(n_610),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_643),
.B(n_641),
.C(n_644),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_646),
.B(n_606),
.C(n_585),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_648),
.B(n_613),
.Y(n_650)
);

NOR3xp33_ASAP7_75t_L g651 ( 
.A(n_647),
.B(n_587),
.C(n_474),
.Y(n_651)
);

NAND4xp75_ASAP7_75t_L g652 ( 
.A(n_650),
.B(n_649),
.C(n_651),
.D(n_584),
.Y(n_652)
);

NOR2x1_ASAP7_75t_L g653 ( 
.A(n_650),
.B(n_617),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_650),
.B(n_534),
.Y(n_654)
);

OA22x2_ASAP7_75t_L g655 ( 
.A1(n_650),
.A2(n_591),
.B1(n_580),
.B2(n_605),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_650),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_656),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_655),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_654),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_653),
.Y(n_660)
);

OAI22x1_ASAP7_75t_L g661 ( 
.A1(n_652),
.A2(n_576),
.B1(n_551),
.B2(n_523),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_657),
.B(n_486),
.C(n_498),
.Y(n_662)
);

OR3x2_ASAP7_75t_L g663 ( 
.A(n_659),
.B(n_473),
.C(n_547),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_660),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_658),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_661),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_665),
.B(n_486),
.C(n_513),
.Y(n_667)
);

OAI22x1_ASAP7_75t_L g668 ( 
.A1(n_664),
.A2(n_551),
.B1(n_523),
.B2(n_509),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_666),
.A2(n_509),
.B1(n_551),
.B2(n_560),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_662),
.A2(n_584),
.B(n_581),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_667),
.A2(n_663),
.B1(n_571),
.B2(n_569),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_670),
.B(n_571),
.Y(n_672)
);

OAI211xp5_ASAP7_75t_SL g673 ( 
.A1(n_668),
.A2(n_562),
.B(n_547),
.C(n_536),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_669),
.B(n_538),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_674),
.A2(n_473),
.B1(n_538),
.B2(n_540),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_675),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_672),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_677),
.A2(n_673),
.B1(n_671),
.B2(n_473),
.Y(n_678)
);


endmodule