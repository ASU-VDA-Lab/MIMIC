module real_aes_6762_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_0), .A2(n_200), .B(n_203), .C(n_284), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_1), .A2(n_233), .B(n_311), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g153 ( .A1(n_2), .A2(n_10), .B1(n_154), .B2(n_157), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_3), .B(n_300), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_4), .A2(n_81), .B1(n_82), .B2(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_4), .Y(n_526) );
INVx1_ASAP7_75t_L g186 ( .A(n_5), .Y(n_186) );
AND2x6_ASAP7_75t_L g200 ( .A(n_5), .B(n_184), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_5), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g274 ( .A(n_6), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_7), .B(n_211), .Y(n_286) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_8), .A2(n_26), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g219 ( .A(n_9), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_11), .A2(n_209), .B(n_296), .C(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_12), .B(n_300), .Y(n_299) );
AOI22xp33_ASAP7_75t_SL g135 ( .A1(n_13), .A2(n_51), .B1(n_136), .B2(n_139), .Y(n_135) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_14), .A2(n_28), .B1(n_90), .B2(n_94), .Y(n_93) );
AOI22xp33_ASAP7_75t_SL g144 ( .A1(n_15), .A2(n_32), .B1(n_145), .B2(n_148), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_16), .B(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_17), .A2(n_314), .B(n_329), .C(n_331), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_18), .B(n_211), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_19), .B(n_211), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_20), .Y(n_250) );
INVx1_ASAP7_75t_L g207 ( .A(n_21), .Y(n_207) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_22), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_23), .Y(n_282) );
AOI22xp5_ASAP7_75t_SL g517 ( .A1(n_23), .A2(n_81), .B1(n_82), .B2(n_282), .Y(n_517) );
INVx1_ASAP7_75t_L g239 ( .A(n_24), .Y(n_239) );
INVx2_ASAP7_75t_L g198 ( .A(n_25), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_27), .Y(n_288) );
OAI221xp5_ASAP7_75t_L g177 ( .A1(n_28), .A2(n_42), .B1(n_50), .B2(n_178), .C(n_179), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_28), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g125 ( .A1(n_29), .A2(n_72), .B1(n_126), .B2(n_130), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g313 ( .A1(n_30), .A2(n_314), .B(n_315), .C(n_317), .Y(n_313) );
INVxp67_ASAP7_75t_L g240 ( .A(n_31), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_33), .A2(n_166), .B1(n_167), .B2(n_173), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_33), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_34), .A2(n_203), .B(n_206), .C(n_214), .Y(n_202) );
CKINVDCx14_ASAP7_75t_R g312 ( .A(n_35), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_36), .A2(n_258), .B(n_272), .C(n_273), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_37), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_38), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_39), .B(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_40), .A2(n_76), .B1(n_171), .B2(n_172), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_40), .Y(n_171) );
INVx1_ASAP7_75t_L g327 ( .A(n_41), .Y(n_327) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_42), .A2(n_63), .B1(n_90), .B2(n_94), .Y(n_97) );
INVxp67_ASAP7_75t_L g181 ( .A(n_42), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g270 ( .A(n_43), .Y(n_270) );
INVx1_ASAP7_75t_L g184 ( .A(n_44), .Y(n_184) );
INVx1_ASAP7_75t_L g218 ( .A(n_45), .Y(n_218) );
INVx1_ASAP7_75t_SL g316 ( .A(n_46), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_47), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_48), .B(n_300), .Y(n_333) );
INVx1_ASAP7_75t_L g253 ( .A(n_49), .Y(n_253) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_50), .A2(n_69), .B1(n_90), .B2(n_91), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_52), .A2(n_233), .B(n_269), .Y(n_268) );
AOI22xp33_ASAP7_75t_SL g159 ( .A1(n_53), .A2(n_67), .B1(n_160), .B2(n_162), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_54), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_55), .A2(n_233), .B(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_56), .A2(n_232), .B(n_234), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_57), .Y(n_201) );
INVx1_ASAP7_75t_L g294 ( .A(n_58), .Y(n_294) );
AOI22xp33_ASAP7_75t_SL g101 ( .A1(n_59), .A2(n_71), .B1(n_102), .B2(n_107), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_60), .B(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_61), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_61), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_61), .A2(n_233), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g297 ( .A(n_62), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_64), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_64), .Y(n_80) );
INVx2_ASAP7_75t_L g216 ( .A(n_65), .Y(n_216) );
INVx1_ASAP7_75t_L g285 ( .A(n_66), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_68), .A2(n_203), .B(n_252), .C(n_260), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_70), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_73), .B(n_223), .Y(n_275) );
INVx1_ASAP7_75t_L g90 ( .A(n_74), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_74), .Y(n_92) );
INVx2_ASAP7_75t_L g330 ( .A(n_75), .Y(n_330) );
INVx1_ASAP7_75t_L g172 ( .A(n_76), .Y(n_172) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_174), .B1(n_187), .B2(n_512), .C(n_516), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_165), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND3x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_134), .C(n_152), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_111), .Y(n_84) );
OAI21xp5_ASAP7_75t_SL g85 ( .A1(n_86), .A2(n_100), .B(n_101), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x6_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x4_ASAP7_75t_L g108 ( .A(n_88), .B(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_93), .Y(n_88) );
AND2x2_ASAP7_75t_L g106 ( .A(n_89), .B(n_97), .Y(n_106) );
INVx2_ASAP7_75t_L g116 ( .A(n_89), .Y(n_116) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
AND2x2_ASAP7_75t_L g115 ( .A(n_93), .B(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g124 ( .A(n_93), .B(n_116), .Y(n_124) );
INVx2_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
AND2x4_ASAP7_75t_L g138 ( .A(n_95), .B(n_115), .Y(n_138) );
AND2x6_ASAP7_75t_L g156 ( .A(n_95), .B(n_123), .Y(n_156) );
AND2x2_ASAP7_75t_L g161 ( .A(n_95), .B(n_147), .Y(n_161) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g117 ( .A(n_96), .B(n_99), .Y(n_117) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g143 ( .A(n_97), .B(n_110), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_97), .B(n_99), .Y(n_151) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g105 ( .A(n_99), .Y(n_105) );
INVx1_ASAP7_75t_L g110 ( .A(n_99), .Y(n_110) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g128 ( .A(n_105), .B(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g127 ( .A(n_106), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g131 ( .A(n_106), .B(n_132), .Y(n_131) );
BUFx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_118), .C(n_125), .Y(n_111) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND2x2_ASAP7_75t_L g142 ( .A(n_115), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g147 ( .A(n_116), .B(n_129), .Y(n_147) );
AND2x4_ASAP7_75t_L g122 ( .A(n_117), .B(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g146 ( .A(n_117), .B(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx5_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x6_ASAP7_75t_L g150 ( .A(n_133), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_144), .Y(n_134) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx6_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx8_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g158 ( .A(n_143), .B(n_147), .Y(n_158) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g163 ( .A(n_147), .B(n_164), .Y(n_163) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx6_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_159), .Y(n_152) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx11_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx2_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
BUFx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_167), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
AND3x1_ASAP7_75t_SL g176 ( .A(n_177), .B(n_182), .C(n_185), .Y(n_176) );
INVxp67_ASAP7_75t_L g521 ( .A(n_177), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_182), .A2(n_514), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g528 ( .A(n_182), .Y(n_528) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OAI322xp33_ASAP7_75t_L g516 ( .A1(n_183), .A2(n_285), .A3(n_517), .B1(n_518), .B2(n_522), .C1(n_525), .C2(n_527), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_183), .B(n_186), .Y(n_524) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_SL g527 ( .A(n_185), .B(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR4x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_402), .C(n_449), .D(n_489), .Y(n_188) );
NAND3xp33_ASAP7_75t_SL g189 ( .A(n_190), .B(n_348), .C(n_377), .Y(n_189) );
AOI211xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_263), .B(n_301), .C(n_341), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_191), .A2(n_361), .B(n_378), .C(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_225), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_193), .B(n_340), .Y(n_339) );
INVx3_ASAP7_75t_SL g344 ( .A(n_193), .Y(n_344) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_193), .Y(n_356) );
AND2x4_ASAP7_75t_L g360 ( .A(n_193), .B(n_308), .Y(n_360) );
AND2x2_ASAP7_75t_L g371 ( .A(n_193), .B(n_248), .Y(n_371) );
OR2x2_ASAP7_75t_L g395 ( .A(n_193), .B(n_304), .Y(n_395) );
AND2x2_ASAP7_75t_L g408 ( .A(n_193), .B(n_309), .Y(n_408) );
AND2x2_ASAP7_75t_L g448 ( .A(n_193), .B(n_434), .Y(n_448) );
AND2x2_ASAP7_75t_L g455 ( .A(n_193), .B(n_418), .Y(n_455) );
AND2x2_ASAP7_75t_L g485 ( .A(n_193), .B(n_226), .Y(n_485) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_220), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_201), .B(n_202), .C(n_215), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_195), .A2(n_250), .B(n_251), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_195), .A2(n_282), .B(n_283), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_196), .B(n_200), .Y(n_195) );
AND2x4_ASAP7_75t_L g233 ( .A(n_196), .B(n_200), .Y(n_233) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
INVx1_ASAP7_75t_L g213 ( .A(n_197), .Y(n_213) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g204 ( .A(n_198), .Y(n_204) );
INVx1_ASAP7_75t_L g332 ( .A(n_198), .Y(n_332) );
INVx1_ASAP7_75t_L g205 ( .A(n_199), .Y(n_205) );
INVx3_ASAP7_75t_L g209 ( .A(n_199), .Y(n_209) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_199), .Y(n_211) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_199), .Y(n_242) );
BUFx3_ASAP7_75t_L g214 ( .A(n_200), .Y(n_214) );
INVx4_ASAP7_75t_SL g243 ( .A(n_200), .Y(n_243) );
INVx5_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
AND2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
BUFx3_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_204), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_210), .C(n_212), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_208), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_238) );
INVx5_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_209), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
INVx4_ASAP7_75t_L g314 ( .A(n_211), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_212), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_213), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_214), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_215), .A2(n_268), .B(n_275), .Y(n_267) );
INVx1_ASAP7_75t_L g280 ( .A(n_215), .Y(n_280) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g224 ( .A(n_216), .B(n_217), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_249), .B(n_261), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_222), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
INVx4_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_223), .Y(n_291) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g230 ( .A(n_224), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_225), .B(n_412), .Y(n_424) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_247), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_226), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g362 ( .A(n_226), .B(n_247), .Y(n_362) );
BUFx3_ASAP7_75t_L g370 ( .A(n_226), .Y(n_370) );
OR2x2_ASAP7_75t_L g391 ( .A(n_226), .B(n_266), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_226), .B(n_412), .Y(n_502) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_231), .B(n_244), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_228), .A2(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g305 ( .A(n_231), .Y(n_305) );
BUFx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_236), .B(n_237), .C(n_243), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_236), .A2(n_243), .B(n_270), .C(n_271), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_SL g293 ( .A1(n_236), .A2(n_243), .B(n_294), .C(n_295), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_236), .A2(n_243), .B(n_312), .C(n_313), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_236), .A2(n_243), .B(n_327), .C(n_328), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_241), .B(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_241), .B(n_330), .Y(n_329) );
INVx4_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g255 ( .A(n_242), .Y(n_255) );
INVx1_ASAP7_75t_L g260 ( .A(n_243), .Y(n_260) );
INVx1_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_246), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g307 ( .A(n_247), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g355 ( .A(n_247), .Y(n_355) );
AND2x2_ASAP7_75t_L g418 ( .A(n_247), .B(n_309), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_247), .A2(n_421), .B1(n_423), .B2(n_425), .C(n_426), .Y(n_420) );
AND2x2_ASAP7_75t_L g434 ( .A(n_247), .B(n_304), .Y(n_434) );
AND2x2_ASAP7_75t_L g460 ( .A(n_247), .B(n_344), .Y(n_460) );
INVx2_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g340 ( .A(n_248), .B(n_309), .Y(n_340) );
BUFx2_ASAP7_75t_L g474 ( .A(n_248), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_256), .C(n_257), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g284 ( .A1(n_254), .A2(n_257), .B(n_285), .C(n_286), .Y(n_284) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_254), .Y(n_515) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g298 ( .A(n_259), .Y(n_298) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI32xp33_ASAP7_75t_L g440 ( .A1(n_264), .A2(n_401), .A3(n_415), .B1(n_441), .B2(n_442), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_276), .Y(n_264) );
AND2x2_ASAP7_75t_L g381 ( .A(n_265), .B(n_323), .Y(n_381) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g363 ( .A(n_266), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_266), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g435 ( .A(n_266), .B(n_323), .Y(n_435) );
AND2x2_ASAP7_75t_L g446 ( .A(n_266), .B(n_338), .Y(n_446) );
BUFx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g347 ( .A(n_267), .B(n_324), .Y(n_347) );
AND2x2_ASAP7_75t_L g351 ( .A(n_267), .B(n_324), .Y(n_351) );
AND2x2_ASAP7_75t_L g386 ( .A(n_267), .B(n_337), .Y(n_386) );
AND2x2_ASAP7_75t_L g393 ( .A(n_267), .B(n_289), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_267), .A2(n_344), .B(n_355), .C(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g452 ( .A(n_267), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_267), .B(n_278), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_276), .B(n_335), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_276), .B(n_351), .Y(n_441) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g346 ( .A(n_277), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_289), .Y(n_277) );
AND2x2_ASAP7_75t_L g338 ( .A(n_278), .B(n_290), .Y(n_338) );
OR2x2_ASAP7_75t_L g353 ( .A(n_278), .B(n_290), .Y(n_353) );
AND2x2_ASAP7_75t_L g376 ( .A(n_278), .B(n_337), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_278), .Y(n_380) );
AND2x2_ASAP7_75t_L g399 ( .A(n_278), .B(n_336), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_278), .A2(n_364), .B1(n_410), .B2(n_411), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_278), .B(n_452), .Y(n_476) );
AND2x2_ASAP7_75t_L g491 ( .A(n_278), .B(n_351), .Y(n_491) );
INVx4_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx3_ASAP7_75t_L g321 ( .A(n_279), .Y(n_321) );
AND2x2_ASAP7_75t_L g365 ( .A(n_279), .B(n_290), .Y(n_365) );
AND2x2_ASAP7_75t_L g367 ( .A(n_279), .B(n_323), .Y(n_367) );
AND3x2_ASAP7_75t_L g429 ( .A(n_279), .B(n_393), .C(n_430), .Y(n_429) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_287), .Y(n_279) );
AND2x2_ASAP7_75t_L g464 ( .A(n_289), .B(n_336), .Y(n_464) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g323 ( .A(n_290), .B(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_290), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_290), .B(n_335), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_290), .B(n_376), .C(n_452), .Y(n_504) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_299), .Y(n_290) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_291), .A2(n_310), .B(n_319), .Y(n_309) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_291), .A2(n_325), .B(n_333), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_320), .B1(n_334), .B2(n_339), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_304), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g416 ( .A(n_304), .Y(n_416) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_307), .A2(n_433), .A3(n_434), .B(n_435), .Y(n_432) );
AND2x2_ASAP7_75t_L g457 ( .A(n_307), .B(n_344), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_307), .B(n_370), .Y(n_503) );
AND2x2_ASAP7_75t_L g412 ( .A(n_308), .B(n_344), .Y(n_412) );
AND2x2_ASAP7_75t_L g473 ( .A(n_308), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g343 ( .A(n_309), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g401 ( .A(n_309), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_314), .B(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_321), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_322), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AOI221x1_ASAP7_75t_SL g389 ( .A1(n_323), .A2(n_390), .B1(n_392), .B2(n_394), .C(n_396), .Y(n_389) );
INVx2_ASAP7_75t_L g337 ( .A(n_324), .Y(n_337) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_324), .Y(n_431) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g419 ( .A(n_334), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_335), .B(n_352), .Y(n_444) );
INVx1_ASAP7_75t_SL g507 ( .A(n_335), .Y(n_507) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g425 ( .A(n_338), .B(n_351), .Y(n_425) );
INVx1_ASAP7_75t_L g493 ( .A(n_339), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_339), .B(n_422), .Y(n_506) );
INVx2_ASAP7_75t_SL g345 ( .A(n_340), .Y(n_345) );
AND2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_344), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_340), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_340), .B(n_415), .Y(n_442) );
AOI21xp33_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_345), .B(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_343), .B(n_415), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_343), .B(n_370), .Y(n_511) );
OR2x2_ASAP7_75t_L g383 ( .A(n_344), .B(n_362), .Y(n_383) );
AND2x2_ASAP7_75t_L g482 ( .A(n_344), .B(n_473), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g357 ( .A1(n_345), .A2(n_358), .B1(n_363), .B2(n_366), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_345), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g405 ( .A(n_347), .B(n_353), .Y(n_405) );
INVx1_ASAP7_75t_L g469 ( .A(n_347), .Y(n_469) );
AOI311xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_354), .A3(n_356), .B(n_357), .C(n_368), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_352), .A2(n_484), .B1(n_496), .B2(n_499), .C(n_501), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_352), .B(n_507), .Y(n_509) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_397), .B(n_398), .C(n_400), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_359), .A2(n_361), .B(n_466), .C(n_467), .Y(n_465) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_360), .B(n_434), .Y(n_500) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_363), .A2(n_383), .B1(n_384), .B2(n_387), .C(n_389), .Y(n_382) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g385 ( .A(n_365), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g468 ( .A(n_365), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_369), .A2(n_427), .B(n_428), .C(n_432), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_370), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_370), .B(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g392 ( .A(n_376), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_380), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g494 ( .A(n_383), .Y(n_494) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_386), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g421 ( .A(n_386), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g498 ( .A(n_386), .Y(n_498) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g439 ( .A(n_388), .B(n_415), .Y(n_439) );
INVx1_ASAP7_75t_SL g433 ( .A(n_395), .Y(n_433) );
INVx1_ASAP7_75t_L g410 ( .A(n_401), .Y(n_410) );
NAND3xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_420), .C(n_436), .Y(n_402) );
AOI322xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .A3(n_407), .B1(n_409), .B2(n_413), .C1(n_417), .C2(n_419), .Y(n_403) );
AOI211xp5_ASAP7_75t_L g456 ( .A1(n_404), .A2(n_457), .B(n_458), .C(n_465), .Y(n_456) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_407), .A2(n_428), .B1(n_459), .B2(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g417 ( .A(n_415), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g454 ( .A(n_415), .B(n_455), .Y(n_454) );
AOI32xp33_ASAP7_75t_L g505 ( .A1(n_415), .A2(n_506), .A3(n_507), .B1(n_508), .B2(n_510), .Y(n_505) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g427 ( .A(n_418), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_418), .A2(n_471), .B1(n_475), .B2(n_477), .C(n_480), .Y(n_470) );
AND2x2_ASAP7_75t_L g484 ( .A(n_418), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g487 ( .A(n_422), .B(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g497 ( .A(n_422), .B(n_498), .Y(n_497) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_452), .Y(n_488) );
AOI211xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B(n_440), .C(n_443), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B(n_447), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_453), .B(n_456), .C(n_470), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_464), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g479 ( .A(n_476), .Y(n_479) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B(n_486), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI211xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_492), .B(n_495), .C(n_505), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx14_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
endmodule