module fake_jpeg_10012_n_233 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_25),
.Y(n_44)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_26),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_30),
.A2(n_28),
.B1(n_20),
.B2(n_14),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_34),
.B1(n_37),
.B2(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_62),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_67),
.B(n_71),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_28),
.B1(n_27),
.B2(n_22),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_17),
.B(n_23),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_36),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_37),
.B1(n_38),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_74),
.B1(n_76),
.B2(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_34),
.B1(n_22),
.B2(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_55),
.B1(n_50),
.B2(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_57),
.B1(n_32),
.B2(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_32),
.B1(n_27),
.B2(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_83),
.B1(n_90),
.B2(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_49),
.B1(n_52),
.B2(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_14),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_91),
.CI(n_94),
.CON(n_112),
.SN(n_112)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_40),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_95),
.B(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_102),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_16),
.B(n_23),
.C(n_21),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_20),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_97),
.B(n_80),
.C(n_89),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_40),
.CI(n_58),
.CON(n_94),
.SN(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_20),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_99),
.C(n_101),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_58),
.C(n_51),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_116),
.B1(n_110),
.B2(n_94),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_73),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_110),
.B(n_113),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_123),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_59),
.B(n_69),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_58),
.C(n_75),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_115),
.C(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_70),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_63),
.C(n_78),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_2),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_119),
.B(n_82),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_63),
.C(n_78),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_19),
.B(n_17),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_2),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_93),
.B(n_94),
.C(n_95),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_134),
.B(n_123),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_118),
.C(n_112),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_112),
.C(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_88),
.B1(n_70),
.B2(n_78),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_106),
.B1(n_112),
.B2(n_117),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_88),
.B1(n_84),
.B2(n_70),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_102),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_90),
.B1(n_63),
.B2(n_20),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_161),
.B1(n_162),
.B2(n_126),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_119),
.C(n_109),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_157),
.Y(n_175)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_155),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_124),
.B(n_18),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_98),
.C(n_122),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_122),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_51),
.B1(n_18),
.B2(n_13),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_51),
.B1(n_18),
.B2(n_13),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_168),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_138),
.B1(n_161),
.B2(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_157),
.B1(n_146),
.B2(n_152),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_139),
.B1(n_131),
.B2(n_126),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_124),
.B1(n_127),
.B2(n_131),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_124),
.B1(n_128),
.B2(n_134),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_176),
.B1(n_124),
.B2(n_18),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_160),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_18),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_177),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_148),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_185),
.C(n_189),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_156),
.C(n_150),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_176),
.B1(n_164),
.B2(n_5),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_191),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_18),
.C(n_12),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_2),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_166),
.B1(n_169),
.B2(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_188),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_3),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_184),
.B(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_3),
.B(n_4),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_196),
.B1(n_6),
.B2(n_7),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_195),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_218),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_192),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_6),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_210),
.B1(n_209),
.B2(n_211),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_193),
.C(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_220),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_11),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_214),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_7),
.Y(n_225)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_227),
.Y(n_229)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_221),
.B(n_213),
.Y(n_228)
);

A2O1A1O1Ixp25_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_225),
.B(n_215),
.C(n_226),
.D(n_9),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_10),
.B(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_231),
.B(n_10),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_10),
.Y(n_233)
);


endmodule