module fake_jpeg_16901_n_63 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_13),
.B1(n_9),
.B2(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_35),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_20),
.B1(n_21),
.B2(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_18),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_11),
.B(n_15),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_34),
.C(n_35),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_10),
.C(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_30),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_16),
.B1(n_10),
.B2(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_18),
.C(n_17),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_12),
.B1(n_16),
.B2(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_31),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.C(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_39),
.C(n_48),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_45),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_56),
.B(n_44),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_5),
.B(n_7),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_51),
.B(n_1),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_5),
.B1(n_7),
.B2(n_3),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_3),
.B2(n_1),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_0),
.B(n_1),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_2),
.Y(n_63)
);


endmodule