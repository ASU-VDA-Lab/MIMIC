module fake_jpeg_7809_n_325 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_24),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_29),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_48),
.B(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_26),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_31),
.B1(n_28),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_31),
.B1(n_28),
.B2(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_31),
.B1(n_28),
.B2(n_33),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_60),
.B1(n_70),
.B2(n_33),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_35),
.B1(n_21),
.B2(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_67),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_18),
.B1(n_17),
.B2(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_17),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_56),
.B(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_78),
.Y(n_123)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_83),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_34),
.B1(n_19),
.B2(n_23),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_94),
.B(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_40),
.Y(n_134)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_88),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_105),
.C(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_102),
.Y(n_114)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_30),
.B1(n_19),
.B2(n_34),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_107),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_55),
.B(n_32),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_38),
.C(n_39),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_40),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_126),
.C(n_130),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_93),
.B1(n_104),
.B2(n_72),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_43),
.B1(n_50),
.B2(n_64),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_108),
.B1(n_80),
.B2(n_75),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_14),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_137),
.B(n_128),
.C(n_123),
.D(n_127),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_105),
.B1(n_79),
.B2(n_84),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_131),
.B1(n_117),
.B2(n_92),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_54),
.B1(n_69),
.B2(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_66),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_12),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_73),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_148),
.C(n_169),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_156),
.B1(n_116),
.B2(n_129),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_140),
.A2(n_165),
.B(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_91),
.B1(n_98),
.B2(n_76),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_143),
.B1(n_20),
.B2(n_27),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_111),
.B1(n_113),
.B2(n_135),
.Y(n_143)
);

AOI222xp33_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_127),
.B1(n_137),
.B2(n_134),
.C1(n_117),
.C2(n_81),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_122),
.B(n_121),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_151),
.B1(n_152),
.B2(n_115),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_96),
.B1(n_106),
.B2(n_69),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_106),
.B1(n_96),
.B2(n_75),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_45),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_8),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_86),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_164),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_0),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_45),
.B(n_62),
.Y(n_179)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

AOI22x1_ASAP7_75t_SL g162 ( 
.A1(n_118),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_162)
);

FAx1_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_20),
.CI(n_22),
.CON(n_174),
.SN(n_174)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_78),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_90),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_45),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_22),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_129),
.C(n_121),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_159),
.B1(n_139),
.B2(n_142),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_168),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_180),
.A2(n_160),
.B(n_154),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_62),
.C(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_198),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_192),
.B(n_176),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_133),
.B1(n_136),
.B2(n_109),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_194),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_136),
.B1(n_109),
.B2(n_103),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_41),
.B1(n_109),
.B2(n_45),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_199),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_45),
.C(n_41),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_202),
.C(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_164),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_45),
.C(n_41),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_203),
.B(n_212),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_221),
.B(n_229),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_222),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_217),
.C(n_225),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_158),
.C(n_153),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g220 ( 
.A(n_176),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_161),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_171),
.B(n_41),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_200),
.Y(n_225)
);

NOR4xp25_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_185),
.C(n_183),
.D(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_247),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_199),
.B1(n_196),
.B2(n_175),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_175),
.B1(n_190),
.B2(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_237),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_177),
.B(n_194),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_242),
.B(n_10),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_179),
.B(n_190),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_208),
.B1(n_204),
.B2(n_206),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_252),
.B1(n_205),
.B2(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_191),
.C(n_182),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_246),
.C(n_217),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_182),
.C(n_174),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_223),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_193),
.B1(n_174),
.B2(n_184),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_228),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_193),
.B1(n_184),
.B2(n_150),
.Y(n_252)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_228),
.B(n_209),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_269),
.Y(n_286)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_221),
.B(n_216),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_264),
.B1(n_254),
.B2(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_267),
.C(n_268),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_207),
.B1(n_222),
.B2(n_150),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_239),
.B1(n_249),
.B2(n_232),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_270),
.Y(n_274)
);

OAI322xp33_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_95),
.A3(n_77),
.B1(n_41),
.B2(n_11),
.C1(n_5),
.C2(n_6),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_16),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_41),
.C(n_2),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_1),
.C(n_2),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_1),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_9),
.B(n_15),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_277),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_248),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_280),
.C(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_278),
.B1(n_270),
.B2(n_242),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_284),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_248),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_245),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_246),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_247),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_254),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_294),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_295),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_283),
.A2(n_253),
.B1(n_266),
.B2(n_258),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_266),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_236),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_236),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_271),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_260),
.B(n_256),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_301),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_297),
.A2(n_243),
.B1(n_238),
.B2(n_247),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_306),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_256),
.B(n_238),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_307),
.B(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_280),
.C(n_2),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_289),
.B1(n_4),
.B2(n_3),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_297),
.B(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_296),
.B(n_292),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_316),
.A3(n_311),
.B1(n_315),
.B2(n_301),
.C1(n_307),
.C2(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_289),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_6),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_12),
.A3(n_15),
.B1(n_6),
.B2(n_7),
.C1(n_16),
.C2(n_13),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_15),
.B(n_3),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_318),
.B(n_320),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_3),
.Y(n_325)
);


endmodule