module fake_jpeg_5967_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_31),
.Y(n_53)
);

BUFx2_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_23),
.B1(n_38),
.B2(n_19),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_17),
.B1(n_20),
.B2(n_19),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_34),
.B1(n_29),
.B2(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_23),
.B1(n_33),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_23),
.B1(n_33),
.B2(n_25),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_33),
.B1(n_17),
.B2(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_28),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_84),
.B1(n_34),
.B2(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_70),
.B(n_78),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_72),
.Y(n_111)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_76),
.Y(n_118)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_28),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_48),
.B1(n_22),
.B2(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_34),
.B1(n_22),
.B2(n_28),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_44),
.B1(n_22),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_99),
.B1(n_108),
.B2(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_103),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_102),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_58),
.B(n_48),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_30),
.B(n_35),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_47),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_106),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_45),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_58),
.B1(n_46),
.B2(n_59),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_116),
.B1(n_74),
.B2(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_113),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_115),
.B1(n_76),
.B2(n_81),
.Y(n_128)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_74),
.B1(n_49),
.B2(n_39),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_126),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_128),
.B1(n_21),
.B2(n_109),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_131),
.B1(n_141),
.B2(n_144),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_124),
.B(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_133),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_47),
.B(n_65),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_113),
.B(n_105),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_132),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_63),
.B1(n_79),
.B2(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_32),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_42),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_142),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_42),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_36),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_79),
.B1(n_83),
.B2(n_52),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_42),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_83),
.B1(n_52),
.B2(n_65),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_115),
.B1(n_110),
.B2(n_102),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_21),
.B1(n_36),
.B2(n_42),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_154),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_155),
.B(n_167),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_164),
.B1(n_172),
.B2(n_31),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_98),
.B(n_117),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_98),
.C(n_117),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_160),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_104),
.C(n_42),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_109),
.B1(n_36),
.B2(n_21),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_120),
.B1(n_123),
.B2(n_134),
.Y(n_176)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_31),
.B(n_32),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_122),
.B(n_126),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_26),
.Y(n_191)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_144),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_122),
.B(n_36),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_189),
.B1(n_0),
.B2(n_1),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_126),
.B(n_138),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_178),
.A2(n_181),
.B(n_174),
.Y(n_215)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_145),
.A2(n_141),
.B1(n_112),
.B2(n_129),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_26),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_171),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_195),
.C(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_156),
.B1(n_163),
.B2(n_145),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_16),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_26),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_150),
.B(n_15),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_169),
.B(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_211),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_204),
.C(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_159),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_165),
.C(n_148),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_214),
.C(n_215),
.Y(n_220)
);

AOI221x1_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_160),
.B1(n_26),
.B2(n_15),
.C(n_31),
.Y(n_210)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_173),
.A2(n_26),
.B1(n_1),
.B2(n_3),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_212),
.B(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_13),
.C(n_4),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_3),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_223),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_195),
.C(n_175),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_191),
.C(n_190),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_183),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_5),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_179),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_231),
.B(n_188),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_176),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_189),
.C(n_192),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_6),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_215),
.B(n_198),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_243),
.B1(n_220),
.B2(n_222),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_213),
.B1(n_197),
.B2(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_221),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_208),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_224),
.A2(n_211),
.B1(n_202),
.B2(n_188),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_234),
.B1(n_232),
.B2(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_223),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_253),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_254),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_224),
.Y(n_253)
);

NAND2xp67_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_220),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_239),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_259),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_218),
.B1(n_244),
.B2(n_8),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_9),
.Y(n_267)
);

AOI21x1_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_6),
.B(n_7),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_9),
.B(n_10),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_7),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_7),
.B(n_9),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_248),
.B1(n_255),
.B2(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_268),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_10),
.B(n_12),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_257),
.A3(n_256),
.B1(n_261),
.B2(n_259),
.C1(n_10),
.C2(n_11),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_12),
.C(n_272),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_270),
.C(n_274),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_276),
.Y(n_277)
);


endmodule