module real_aes_10938_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1382;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_1893;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_1945;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_1404;
wire n_602;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1580;
wire n_1000;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1691;
wire n_1176;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_0), .A2(n_575), .B1(n_578), .B2(n_587), .C(n_590), .Y(n_574) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_0), .A2(n_646), .B(n_648), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_1), .A2(n_357), .B1(n_413), .B2(n_640), .Y(n_1307) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1), .Y(n_1334) );
INVx1_ASAP7_75t_L g1345 ( .A(n_2), .Y(n_1345) );
OAI221xp5_ASAP7_75t_L g1374 ( .A1(n_2), .A2(n_193), .B1(n_1375), .B2(n_1376), .C(n_1377), .Y(n_1374) );
INVxp67_ASAP7_75t_L g1899 ( .A(n_3), .Y(n_1899) );
AOI221xp5_ASAP7_75t_L g1924 ( .A1(n_3), .A2(n_205), .B1(n_1916), .B2(n_1925), .C(n_1927), .Y(n_1924) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_4), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g962 ( .A1(n_5), .A2(n_541), .B1(n_895), .B2(n_963), .C(n_969), .Y(n_962) );
INVx1_ASAP7_75t_L g985 ( .A(n_5), .Y(n_985) );
INVx1_ASAP7_75t_L g511 ( .A(n_6), .Y(n_511) );
XNOR2x2_ASAP7_75t_L g1128 ( .A(n_7), .B(n_1129), .Y(n_1128) );
INVxp33_ASAP7_75t_L g1196 ( .A(n_8), .Y(n_1196) );
AOI221xp5_ASAP7_75t_L g1227 ( .A1(n_8), .A2(n_111), .B1(n_1228), .B2(n_1229), .C(n_1230), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_9), .A2(n_82), .B1(n_1091), .B2(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1268 ( .A(n_9), .Y(n_1268) );
CKINVDCx5p33_ASAP7_75t_R g1613 ( .A(n_10), .Y(n_1613) );
OAI221xp5_ASAP7_75t_L g1884 ( .A1(n_11), .A2(n_256), .B1(n_1885), .B2(n_1886), .C(n_1887), .Y(n_1884) );
INVx1_ASAP7_75t_L g1920 ( .A(n_11), .Y(n_1920) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_12), .A2(n_123), .B1(n_516), .B2(n_601), .C(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g990 ( .A(n_12), .Y(n_990) );
INVx1_ASAP7_75t_L g1210 ( .A(n_13), .Y(n_1210) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_14), .A2(n_188), .B1(n_596), .B2(n_599), .C(n_600), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_14), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_15), .A2(n_334), .B1(n_691), .B2(n_692), .C(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g704 ( .A(n_15), .Y(n_704) );
AO22x1_ASAP7_75t_L g947 ( .A1(n_16), .A2(n_948), .B1(n_992), .B2(n_993), .Y(n_947) );
INVx1_ASAP7_75t_L g993 ( .A(n_16), .Y(n_993) );
INVx1_ASAP7_75t_L g1514 ( .A(n_17), .Y(n_1514) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_18), .A2(n_320), .B1(n_761), .B2(n_762), .Y(n_841) );
INVxp33_ASAP7_75t_SL g868 ( .A(n_18), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g1907 ( .A(n_19), .Y(n_1907) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_20), .A2(n_325), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
INVx1_ASAP7_75t_L g1117 ( .A(n_20), .Y(n_1117) );
INVx1_ASAP7_75t_L g1264 ( .A(n_21), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_21), .A2(n_102), .B1(n_557), .B2(n_565), .Y(n_1283) );
INVx1_ASAP7_75t_L g670 ( .A(n_22), .Y(n_670) );
INVxp33_ASAP7_75t_SL g832 ( .A(n_23), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_23), .A2(n_172), .B1(n_405), .B2(n_425), .C(n_852), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_24), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_25), .A2(n_160), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_25), .A2(n_253), .B1(n_425), .B2(n_796), .C(n_799), .Y(n_795) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_26), .A2(n_86), .B1(n_1042), .B2(n_1043), .C(n_1045), .Y(n_1041) );
INVx1_ASAP7_75t_L g1048 ( .A(n_26), .Y(n_1048) );
INVx1_ASAP7_75t_L g1253 ( .A(n_27), .Y(n_1253) );
OAI221xp5_ASAP7_75t_L g1270 ( .A1(n_27), .A2(n_541), .B1(n_1104), .B2(n_1271), .C(n_1274), .Y(n_1270) );
OAI221xp5_ASAP7_75t_L g1891 ( .A1(n_28), .A2(n_127), .B1(n_600), .B2(n_1892), .C(n_1893), .Y(n_1891) );
OAI22xp5_ASAP7_75t_L g1914 ( .A1(n_28), .A2(n_127), .B1(n_1043), .B2(n_1618), .Y(n_1914) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_29), .A2(n_32), .B1(n_692), .B2(n_1134), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_29), .A2(n_285), .B1(n_565), .B2(n_1173), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_30), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_31), .A2(n_207), .B1(n_406), .B2(n_1086), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_31), .A2(n_207), .B1(n_878), .B2(n_879), .Y(n_1093) );
INVxp67_ASAP7_75t_SL g1170 ( .A(n_32), .Y(n_1170) );
AO221x2_ASAP7_75t_L g1696 ( .A1(n_33), .A2(n_270), .B1(n_1653), .B2(n_1674), .C(n_1697), .Y(n_1696) );
CKINVDCx16_ASAP7_75t_R g1705 ( .A(n_34), .Y(n_1705) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_35), .A2(n_226), .B1(n_1075), .B2(n_1077), .Y(n_1074) );
INVxp67_ASAP7_75t_SL g1099 ( .A(n_35), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_36), .A2(n_336), .B1(n_878), .B2(n_879), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_36), .A2(n_336), .B1(n_937), .B2(n_938), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_37), .A2(n_56), .B1(n_504), .B2(n_676), .C(n_677), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_37), .A2(n_295), .B1(n_715), .B2(n_716), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_38), .Y(n_584) );
INVx1_ASAP7_75t_L g679 ( .A(n_39), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_39), .A2(n_56), .B1(n_709), .B2(n_710), .C(n_712), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_40), .A2(n_352), .B1(n_723), .B2(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1486 ( .A(n_40), .Y(n_1486) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_41), .A2(n_83), .B1(n_604), .B2(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g642 ( .A(n_41), .Y(n_642) );
INVx1_ASAP7_75t_L g1152 ( .A(n_42), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_42), .A2(n_182), .B1(n_930), .B2(n_1158), .C(n_1160), .Y(n_1157) );
INVx1_ASAP7_75t_L g696 ( .A(n_43), .Y(n_696) );
INVxp33_ASAP7_75t_L g1594 ( .A(n_44), .Y(n_1594) );
AOI221xp5_ASAP7_75t_L g1619 ( .A1(n_44), .A2(n_110), .B1(n_1248), .B2(n_1620), .C(n_1621), .Y(n_1619) );
AOI22xp33_ASAP7_75t_SL g1603 ( .A1(n_45), .A2(n_176), .B1(n_1604), .B2(n_1605), .Y(n_1603) );
AOI22xp33_ASAP7_75t_L g1629 ( .A1(n_45), .A2(n_176), .B1(n_1630), .B2(n_1631), .Y(n_1629) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_46), .A2(n_142), .B1(n_758), .B2(n_1110), .C(n_1112), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_46), .A2(n_166), .B1(n_1121), .B2(n_1123), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_47), .A2(n_53), .B1(n_691), .B2(n_956), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_47), .A2(n_123), .B1(n_557), .B2(n_565), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_48), .A2(n_307), .B1(n_757), .B2(n_843), .Y(n_842) );
INVxp33_ASAP7_75t_L g867 ( .A(n_48), .Y(n_867) );
INVx1_ASAP7_75t_L g366 ( .A(n_49), .Y(n_366) );
INVx1_ASAP7_75t_L g1182 ( .A(n_50), .Y(n_1182) );
INVx1_ASAP7_75t_L g1442 ( .A(n_51), .Y(n_1442) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_52), .Y(n_1235) );
INVx1_ASAP7_75t_L g989 ( .A(n_53), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_54), .A2(n_192), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
INVx1_ASAP7_75t_L g1278 ( .A(n_54), .Y(n_1278) );
INVx1_ASAP7_75t_L g1155 ( .A(n_55), .Y(n_1155) );
INVx1_ASAP7_75t_L g829 ( .A(n_57), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g1363 ( .A(n_58), .Y(n_1363) );
AOI22xp33_ASAP7_75t_SL g1607 ( .A1(n_59), .A2(n_314), .B1(n_761), .B2(n_1608), .Y(n_1607) );
AOI221xp5_ASAP7_75t_L g1625 ( .A1(n_59), .A2(n_314), .B1(n_1305), .B2(n_1626), .C(n_1627), .Y(n_1625) );
CKINVDCx5p33_ASAP7_75t_R g1418 ( .A(n_60), .Y(n_1418) );
INVx1_ASAP7_75t_L g1084 ( .A(n_61), .Y(n_1084) );
OAI211xp5_ASAP7_75t_SL g1105 ( .A1(n_61), .A2(n_471), .B(n_1106), .C(n_1113), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_62), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g1904 ( .A(n_63), .Y(n_1904) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_64), .A2(n_119), .B1(n_913), .B2(n_960), .Y(n_959) );
OAI22xp5_ASAP7_75t_SL g976 ( .A1(n_64), .A2(n_119), .B1(n_437), .B2(n_449), .Y(n_976) );
XOR2x2_ASAP7_75t_L g732 ( .A(n_65), .B(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_66), .A2(n_356), .B1(n_412), .B2(n_418), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_66), .A2(n_340), .B1(n_541), .B2(n_544), .Y(n_540) );
INVx1_ASAP7_75t_L g1532 ( .A(n_67), .Y(n_1532) );
OAI221xp5_ASAP7_75t_L g1537 ( .A1(n_67), .A2(n_290), .B1(n_1538), .B2(n_1539), .C(n_1540), .Y(n_1537) );
AOI22xp33_ASAP7_75t_SL g1609 ( .A1(n_68), .A2(n_144), .B1(n_761), .B2(n_1605), .Y(n_1609) );
INVxp67_ASAP7_75t_SL g1616 ( .A(n_68), .Y(n_1616) );
INVxp33_ASAP7_75t_L g1180 ( .A(n_69), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_69), .A2(n_133), .B1(n_1220), .B2(n_1222), .C(n_1224), .Y(n_1219) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_70), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g1710 ( .A1(n_71), .A2(n_333), .B1(n_1653), .B2(n_1674), .Y(n_1710) );
INVx1_ASAP7_75t_L g666 ( .A(n_72), .Y(n_666) );
INVxp33_ASAP7_75t_SL g750 ( .A(n_73), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_73), .A2(n_249), .B1(n_784), .B2(n_786), .C(n_788), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g1909 ( .A(n_74), .Y(n_1909) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_75), .A2(n_181), .B1(n_528), .B2(n_586), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_75), .A2(n_181), .B1(n_624), .B2(n_626), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g1549 ( .A1(n_76), .A2(n_339), .B1(n_1043), .B2(n_1550), .Y(n_1549) );
OAI221xp5_ASAP7_75t_L g1570 ( .A1(n_76), .A2(n_339), .B1(n_1187), .B2(n_1189), .C(n_1571), .Y(n_1570) );
INVxp33_ASAP7_75t_L g1195 ( .A(n_77), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_77), .A2(n_283), .B1(n_1024), .B2(n_1232), .Y(n_1231) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_78), .A2(n_238), .B1(n_1187), .B2(n_1189), .C(n_1190), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_78), .A2(n_238), .B1(n_1043), .B2(n_1218), .Y(n_1217) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_79), .A2(n_541), .B1(n_1104), .B2(n_1146), .C(n_1151), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_79), .A2(n_244), .B1(n_412), .B2(n_796), .C(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g974 ( .A(n_80), .Y(n_974) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_81), .A2(n_253), .B1(n_761), .B2(n_762), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_81), .A2(n_160), .B1(n_723), .B2(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g1269 ( .A(n_82), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_83), .A2(n_136), .B1(n_402), .B2(n_640), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_84), .A2(n_322), .B1(n_611), .B2(n_614), .Y(n_1020) );
INVx1_ASAP7_75t_L g1046 ( .A(n_84), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g740 ( .A(n_85), .Y(n_740) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_85), .A2(n_296), .B1(n_779), .B2(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g1049 ( .A(n_86), .Y(n_1049) );
XOR2xp5_ASAP7_75t_L g387 ( .A(n_87), .B(n_388), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g1310 ( .A(n_88), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1454 ( .A(n_89), .Y(n_1454) );
INVx1_ASAP7_75t_L g745 ( .A(n_90), .Y(n_745) );
INVx1_ASAP7_75t_L g507 ( .A(n_91), .Y(n_507) );
INVx1_ASAP7_75t_L g1559 ( .A(n_92), .Y(n_1559) );
AOI22xp33_ASAP7_75t_SL g1610 ( .A1(n_93), .A2(n_130), .B1(n_1604), .B2(n_1608), .Y(n_1610) );
INVxp67_ASAP7_75t_L g1624 ( .A(n_93), .Y(n_1624) );
INVx1_ASAP7_75t_L g1366 ( .A(n_94), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_94), .A2(n_315), .B1(n_402), .B2(n_428), .Y(n_1378) );
INVx1_ASAP7_75t_L g886 ( .A(n_95), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_95), .A2(n_113), .B1(n_400), .B2(n_928), .Y(n_927) );
CKINVDCx5p33_ASAP7_75t_R g1905 ( .A(n_96), .Y(n_1905) );
AOI22xp33_ASAP7_75t_SL g1348 ( .A1(n_97), .A2(n_189), .B1(n_843), .B2(n_1349), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_97), .A2(n_190), .B1(n_1387), .B2(n_1388), .Y(n_1386) );
INVx1_ASAP7_75t_L g1457 ( .A(n_98), .Y(n_1457) );
OAI221xp5_ASAP7_75t_L g1474 ( .A1(n_98), .A2(n_148), .B1(n_599), .B2(n_1187), .C(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1467 ( .A(n_99), .Y(n_1467) );
CKINVDCx5p33_ASAP7_75t_R g1463 ( .A(n_100), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_101), .A2(n_313), .B1(n_400), .B2(n_405), .Y(n_399) );
INVx1_ASAP7_75t_L g478 ( .A(n_101), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_102), .A2(n_349), .B1(n_958), .B2(n_1112), .C(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1254 ( .A(n_103), .Y(n_1254) );
OAI211xp5_ASAP7_75t_L g1260 ( .A1(n_103), .A2(n_471), .B(n_1261), .C(n_1267), .Y(n_1260) );
INVx1_ASAP7_75t_L g1420 ( .A(n_104), .Y(n_1420) );
OAI222xp33_ASAP7_75t_L g1499 ( .A1(n_105), .A2(n_155), .B1(n_308), .B2(n_614), .C1(n_1189), .C2(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1522 ( .A(n_105), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g1464 ( .A1(n_106), .A2(n_224), .B1(n_721), .B2(n_1036), .C(n_1404), .Y(n_1464) );
INVx1_ASAP7_75t_L g1473 ( .A(n_106), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_107), .A2(n_233), .B1(n_406), .B2(n_1086), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_107), .A2(n_233), .B1(n_878), .B2(n_879), .Y(n_1279) );
INVx1_ASAP7_75t_L g1300 ( .A(n_108), .Y(n_1300) );
OAI221xp5_ASAP7_75t_L g1323 ( .A1(n_108), .A2(n_126), .B1(n_1190), .B2(n_1324), .C(n_1325), .Y(n_1323) );
AO22x2_ASAP7_75t_L g994 ( .A1(n_109), .A2(n_995), .B1(n_1050), .B2(n_1051), .Y(n_994) );
CKINVDCx14_ASAP7_75t_R g1050 ( .A(n_109), .Y(n_1050) );
INVxp33_ASAP7_75t_SL g1600 ( .A(n_110), .Y(n_1600) );
INVxp67_ASAP7_75t_L g1199 ( .A(n_111), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g1403 ( .A1(n_112), .A2(n_247), .B1(n_1036), .B2(n_1385), .C(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1427 ( .A(n_112), .Y(n_1427) );
INVx1_ASAP7_75t_L g884 ( .A(n_113), .Y(n_884) );
BUFx2_ASAP7_75t_L g398 ( .A(n_114), .Y(n_398) );
BUFx2_ASAP7_75t_L g432 ( .A(n_114), .Y(n_432) );
INVx1_ASAP7_75t_L g446 ( .A(n_114), .Y(n_446) );
OR2x2_ASAP7_75t_L g598 ( .A(n_114), .B(n_527), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_115), .A2(n_152), .B1(n_528), .B2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g636 ( .A(n_115), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g1309 ( .A(n_116), .Y(n_1309) );
INVx1_ASAP7_75t_L g968 ( .A(n_117), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_117), .A2(n_228), .B1(n_401), .B2(n_787), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_118), .A2(n_122), .B1(n_1357), .B2(n_1359), .Y(n_1356) );
INVx1_ASAP7_75t_L g1391 ( .A(n_118), .Y(n_1391) );
CKINVDCx5p33_ASAP7_75t_R g1548 ( .A(n_120), .Y(n_1548) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_121), .A2(n_212), .B1(n_761), .B2(n_762), .Y(n_764) );
INVxp33_ASAP7_75t_SL g808 ( .A(n_121), .Y(n_808) );
INVx1_ASAP7_75t_L g1383 ( .A(n_122), .Y(n_1383) );
INVx1_ASAP7_75t_L g953 ( .A(n_124), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_124), .A2(n_266), .B1(n_777), .B2(n_787), .Y(n_987) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_125), .Y(n_909) );
INVx1_ASAP7_75t_L g1301 ( .A(n_126), .Y(n_1301) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_128), .A2(n_262), .B1(n_757), .B2(n_758), .Y(n_765) );
INVxp33_ASAP7_75t_L g806 ( .A(n_128), .Y(n_806) );
CKINVDCx16_ASAP7_75t_R g1707 ( .A(n_129), .Y(n_1707) );
INVxp33_ASAP7_75t_L g1633 ( .A(n_130), .Y(n_1633) );
INVx1_ASAP7_75t_L g1081 ( .A(n_131), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_131), .A2(n_541), .B1(n_1095), .B2(n_1097), .C(n_1104), .Y(n_1094) );
INVx1_ASAP7_75t_L g695 ( .A(n_132), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_132), .A2(n_334), .B1(n_700), .B2(n_702), .C(n_703), .Y(n_699) );
INVxp33_ASAP7_75t_L g1185 ( .A(n_133), .Y(n_1185) );
NAND2xp33_ASAP7_75t_SL g1296 ( .A(n_134), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1319 ( .A(n_134), .Y(n_1319) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_135), .A2(n_471), .B1(n_898), .B2(n_903), .C(n_908), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g932 ( .A1(n_135), .A2(n_221), .B1(n_933), .B2(n_935), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_136), .A2(n_149), .B1(n_611), .B2(n_614), .Y(n_610) );
INVx1_ASAP7_75t_L g1598 ( .A(n_137), .Y(n_1598) );
INVx1_ASAP7_75t_L g831 ( .A(n_138), .Y(n_831) );
INVx1_ASAP7_75t_L g1888 ( .A(n_139), .Y(n_1888) );
INVx1_ASAP7_75t_L g1238 ( .A(n_140), .Y(n_1238) );
INVx1_ASAP7_75t_L g893 ( .A(n_141), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_141), .A2(n_146), .B1(n_930), .B2(n_931), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_142), .A2(n_210), .B1(n_557), .B2(n_565), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_143), .Y(n_1419) );
INVxp33_ASAP7_75t_L g1634 ( .A(n_144), .Y(n_1634) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_145), .A2(n_329), .B1(n_1653), .B2(n_1674), .Y(n_1695) );
INVx1_ASAP7_75t_L g890 ( .A(n_146), .Y(n_890) );
INVx1_ASAP7_75t_L g1395 ( .A(n_147), .Y(n_1395) );
INVx1_ASAP7_75t_L g1456 ( .A(n_148), .Y(n_1456) );
INVx1_ASAP7_75t_L g650 ( .A(n_149), .Y(n_650) );
INVxp67_ASAP7_75t_SL g1591 ( .A(n_150), .Y(n_1591) );
OAI22xp33_ASAP7_75t_L g1617 ( .A1(n_150), .A2(n_178), .B1(n_1043), .B2(n_1618), .Y(n_1617) );
AOI22xp5_ASAP7_75t_L g1684 ( .A1(n_151), .A2(n_156), .B1(n_1685), .B2(n_1688), .Y(n_1684) );
INVx1_ASAP7_75t_L g631 ( .A(n_152), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_153), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_154), .A2(n_248), .B1(n_1164), .B2(n_1413), .C(n_1415), .Y(n_1412) );
INVx1_ASAP7_75t_L g1437 ( .A(n_154), .Y(n_1437) );
INVx1_ASAP7_75t_L g1530 ( .A(n_155), .Y(n_1530) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_157), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g1690 ( .A1(n_158), .A2(n_343), .B1(n_1645), .B2(n_1691), .Y(n_1690) );
AO221x2_ASAP7_75t_L g1718 ( .A1(n_159), .A2(n_219), .B1(n_1645), .B2(n_1653), .C(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1149 ( .A(n_161), .Y(n_1149) );
INVx1_ASAP7_75t_L g1650 ( .A(n_162), .Y(n_1650) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_163), .A2(n_285), .B1(n_516), .B2(n_1137), .C(n_1139), .Y(n_1136) );
INVxp67_ASAP7_75t_SL g1171 ( .A(n_163), .Y(n_1171) );
INVx1_ASAP7_75t_L g1651 ( .A(n_164), .Y(n_1651) );
INVx1_ASAP7_75t_L g1003 ( .A(n_165), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1039 ( .A1(n_165), .A2(n_317), .B1(n_787), .B2(n_864), .Y(n_1039) );
INVx1_ASAP7_75t_L g1107 ( .A(n_166), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_167), .Y(n_1402) );
INVx1_ASAP7_75t_L g1184 ( .A(n_168), .Y(n_1184) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_169), .A2(n_209), .B1(n_761), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_169), .A2(n_264), .B1(n_786), .B2(n_863), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g1709 ( .A1(n_170), .A2(n_348), .B1(n_1685), .B2(n_1688), .Y(n_1709) );
INVx1_ASAP7_75t_L g1365 ( .A(n_171), .Y(n_1365) );
AOI21xp33_ASAP7_75t_L g1379 ( .A1(n_171), .A2(n_648), .B(n_1380), .Y(n_1379) );
INVxp33_ASAP7_75t_SL g827 ( .A(n_172), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g1295 ( .A1(n_173), .A2(n_306), .B1(n_406), .B2(n_1087), .Y(n_1295) );
INVx1_ASAP7_75t_L g1318 ( .A(n_173), .Y(n_1318) );
INVx1_ASAP7_75t_L g1648 ( .A(n_174), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1666 ( .A(n_174), .B(n_1660), .Y(n_1666) );
INVx1_ASAP7_75t_L g1508 ( .A(n_175), .Y(n_1508) );
INVx2_ASAP7_75t_L g378 ( .A(n_177), .Y(n_378) );
INVxp67_ASAP7_75t_SL g1592 ( .A(n_178), .Y(n_1592) );
INVxp67_ASAP7_75t_L g1510 ( .A(n_179), .Y(n_1510) );
OAI222xp33_ASAP7_75t_L g1524 ( .A1(n_179), .A2(n_186), .B1(n_278), .B2(n_427), .C1(n_700), .C2(n_1124), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g1557 ( .A(n_180), .Y(n_1557) );
AOI21xp33_ASAP7_75t_L g1153 ( .A1(n_182), .A2(n_588), .B(n_1137), .Y(n_1153) );
BUFx3_ASAP7_75t_L g404 ( .A(n_183), .Y(n_404) );
INVx1_ASAP7_75t_L g410 ( .A(n_183), .Y(n_410) );
INVx1_ASAP7_75t_L g1720 ( .A(n_184), .Y(n_1720) );
XNOR2x2_ASAP7_75t_L g1881 ( .A(n_184), .B(n_1882), .Y(n_1881) );
AOI22xp33_ASAP7_75t_L g1940 ( .A1(n_184), .A2(n_1941), .B1(n_1945), .B2(n_1947), .Y(n_1940) );
INVx1_ASAP7_75t_L g502 ( .A(n_185), .Y(n_502) );
INVxp67_ASAP7_75t_L g1513 ( .A(n_186), .Y(n_1513) );
INVxp67_ASAP7_75t_L g1902 ( .A(n_187), .Y(n_1902) );
AOI22xp33_ASAP7_75t_L g1928 ( .A1(n_187), .A2(n_261), .B1(n_412), .B2(n_1929), .Y(n_1928) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_188), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g1384 ( .A1(n_189), .A2(n_286), .B1(n_633), .B2(n_712), .C(n_1385), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_190), .A2(n_286), .B1(n_1351), .B2(n_1353), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_191), .A2(n_264), .B1(n_757), .B2(n_836), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g858 ( .A1(n_191), .A2(n_209), .B1(n_709), .B2(n_859), .C(n_861), .Y(n_858) );
INVx1_ASAP7_75t_L g1277 ( .A(n_192), .Y(n_1277) );
INVx1_ASAP7_75t_L g1344 ( .A(n_193), .Y(n_1344) );
AOI221xp5_ASAP7_75t_L g1546 ( .A1(n_194), .A2(n_298), .B1(n_648), .B2(n_935), .C(n_1232), .Y(n_1546) );
INVx1_ASAP7_75t_L g1566 ( .A(n_194), .Y(n_1566) );
INVx1_ASAP7_75t_L g998 ( .A(n_195), .Y(n_998) );
AOI21xp33_ASAP7_75t_L g1040 ( .A1(n_195), .A2(n_777), .B(n_861), .Y(n_1040) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_196), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g1304 ( .A1(n_197), .A2(n_269), .B1(n_633), .B2(n_1026), .C(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1329 ( .A(n_197), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_198), .A2(n_287), .B1(n_1407), .B2(n_1408), .Y(n_1406) );
OAI221xp5_ASAP7_75t_L g1429 ( .A1(n_198), .A2(n_287), .B1(n_600), .B2(n_1324), .C(n_1325), .Y(n_1429) );
INVx1_ASAP7_75t_L g1205 ( .A(n_199), .Y(n_1205) );
INVx1_ASAP7_75t_L g1643 ( .A(n_200), .Y(n_1643) );
INVx1_ASAP7_75t_L g680 ( .A(n_201), .Y(n_680) );
INVx1_ASAP7_75t_L g1150 ( .A(n_202), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_203), .A2(n_340), .B1(n_425), .B2(n_426), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_203), .A2(n_356), .B1(n_461), .B2(n_471), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_204), .Y(n_454) );
INVxp67_ASAP7_75t_L g1901 ( .A(n_205), .Y(n_1901) );
INVx1_ASAP7_75t_L g1721 ( .A(n_206), .Y(n_1721) );
INVx1_ASAP7_75t_L g395 ( .A(n_208), .Y(n_395) );
INVx1_ASAP7_75t_L g444 ( .A(n_208), .Y(n_444) );
INVx1_ASAP7_75t_L g1108 ( .A(n_210), .Y(n_1108) );
INVx1_ASAP7_75t_L g1595 ( .A(n_211), .Y(n_1595) );
INVxp67_ASAP7_75t_SL g775 ( .A(n_212), .Y(n_775) );
XNOR2xp5_ASAP7_75t_L g1496 ( .A(n_213), .B(n_1497), .Y(n_1496) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_214), .A2(n_817), .B1(n_818), .B2(n_872), .Y(n_816) );
INVx1_ASAP7_75t_L g872 ( .A(n_214), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g1290 ( .A(n_215), .Y(n_1290) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_216), .A2(n_662), .B(n_697), .Y(n_661) );
INVx1_ASAP7_75t_L g731 ( .A(n_216), .Y(n_731) );
INVx1_ASAP7_75t_L g1679 ( .A(n_216), .Y(n_1679) );
INVxp67_ASAP7_75t_L g1503 ( .A(n_217), .Y(n_1503) );
AOI221xp5_ASAP7_75t_L g1526 ( .A1(n_217), .A2(n_324), .B1(n_633), .B2(n_1026), .C(n_1415), .Y(n_1526) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_218), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_220), .Y(n_1008) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_221), .A2(n_541), .B1(n_881), .B2(n_887), .C(n_895), .Y(n_880) );
XOR2xp5_ASAP7_75t_L g571 ( .A(n_222), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g1175 ( .A(n_223), .Y(n_1175) );
INVx1_ASAP7_75t_L g1471 ( .A(n_224), .Y(n_1471) );
AOI22xp5_ASAP7_75t_L g1694 ( .A1(n_225), .A2(n_292), .B1(n_1685), .B2(n_1688), .Y(n_1694) );
INVxp67_ASAP7_75t_SL g1103 ( .A(n_226), .Y(n_1103) );
INVx1_ASAP7_75t_L g689 ( .A(n_227), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_227), .A2(n_297), .B1(n_648), .B2(n_720), .C(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g966 ( .A(n_228), .Y(n_966) );
INVx1_ASAP7_75t_L g1263 ( .A(n_229), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_229), .A2(n_349), .B1(n_1121), .B2(n_1123), .Y(n_1284) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_230), .Y(n_1448) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_231), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_232), .Y(n_915) );
AOI221xp5_ASAP7_75t_L g1552 ( .A1(n_234), .A2(n_275), .B1(n_931), .B2(n_1220), .C(n_1415), .Y(n_1552) );
INVx1_ASAP7_75t_L g1578 ( .A(n_234), .Y(n_1578) );
INVx1_ASAP7_75t_L g1211 ( .A(n_235), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_236), .A2(n_240), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
INVx1_ASAP7_75t_L g1030 ( .A(n_236), .Y(n_1030) );
OA332x1_ASAP7_75t_L g996 ( .A1(n_237), .A2(n_575), .A3(n_587), .B1(n_997), .B2(n_1002), .B3(n_1006), .C1(n_1010), .C2(n_1015), .Y(n_996) );
AOI21xp5_ASAP7_75t_L g1034 ( .A1(n_237), .A2(n_1035), .B(n_1036), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_239), .A2(n_318), .B1(n_913), .B2(n_960), .Y(n_1141) );
OAI221xp5_ASAP7_75t_L g1168 ( .A1(n_239), .A2(n_318), .B1(n_943), .B2(n_1090), .C(n_1091), .Y(n_1168) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_240), .A2(n_322), .B1(n_777), .B2(n_787), .Y(n_1033) );
CKINVDCx16_ASAP7_75t_R g1675 ( .A(n_241), .Y(n_1675) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_242), .A2(n_251), .B1(n_412), .B2(n_418), .Y(n_411) );
INVx1_ASAP7_75t_L g496 ( .A(n_242), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_243), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1131 ( .A1(n_244), .A2(n_471), .B(n_1132), .C(n_1142), .Y(n_1131) );
INVx1_ASAP7_75t_L g1143 ( .A(n_245), .Y(n_1143) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_246), .Y(n_1453) );
INVx1_ASAP7_75t_L g1425 ( .A(n_247), .Y(n_1425) );
INVx1_ASAP7_75t_L g1434 ( .A(n_248), .Y(n_1434) );
INVxp33_ASAP7_75t_SL g742 ( .A(n_249), .Y(n_742) );
INVx1_ASAP7_75t_L g1521 ( .A(n_250), .Y(n_1521) );
INVx1_ASAP7_75t_L g492 ( .A(n_251), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_252), .Y(n_971) );
INVx1_ASAP7_75t_L g1585 ( .A(n_254), .Y(n_1585) );
INVx1_ASAP7_75t_L g1144 ( .A(n_255), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g1915 ( .A1(n_256), .A2(n_354), .B1(n_1916), .B2(n_1917), .C(n_1918), .Y(n_1915) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_257), .A2(n_288), .B1(n_640), .B2(n_1387), .Y(n_1416) );
INVx1_ASAP7_75t_L g1438 ( .A(n_257), .Y(n_1438) );
INVx1_ASAP7_75t_L g1073 ( .A(n_258), .Y(n_1073) );
CKINVDCx20_ASAP7_75t_R g1635 ( .A(n_259), .Y(n_1635) );
INVx1_ASAP7_75t_L g403 ( .A(n_260), .Y(n_403) );
BUFx3_ASAP7_75t_L g409 ( .A(n_260), .Y(n_409) );
INVxp67_ASAP7_75t_L g1897 ( .A(n_261), .Y(n_1897) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_262), .Y(n_794) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_263), .Y(n_374) );
AND2x2_ASAP7_75t_L g465 ( .A(n_263), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g520 ( .A(n_263), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_263), .B(n_341), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g1449 ( .A1(n_265), .A2(n_321), .B1(n_401), .B2(n_721), .C(n_1305), .Y(n_1449) );
INVx1_ASAP7_75t_L g1480 ( .A(n_265), .Y(n_1480) );
INVx1_ASAP7_75t_L g952 ( .A(n_266), .Y(n_952) );
INVx1_ASAP7_75t_L g1661 ( .A(n_267), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_268), .Y(n_907) );
INVx1_ASAP7_75t_L g1335 ( .A(n_269), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_271), .Y(n_970) );
INVx1_ASAP7_75t_L g1680 ( .A(n_272), .Y(n_1680) );
INVx2_ASAP7_75t_L g396 ( .A(n_273), .Y(n_396) );
OR2x2_ASAP7_75t_L g555 ( .A(n_273), .B(n_444), .Y(n_555) );
INVx1_ASAP7_75t_L g1491 ( .A(n_274), .Y(n_1491) );
INVx1_ASAP7_75t_L g1576 ( .A(n_275), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_276), .A2(n_294), .B1(n_546), .B2(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_276), .A2(n_294), .B1(n_617), .B2(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g1505 ( .A(n_277), .Y(n_1505) );
INVxp67_ASAP7_75t_L g1511 ( .A(n_278), .Y(n_1511) );
CKINVDCx16_ASAP7_75t_R g1677 ( .A(n_279), .Y(n_1677) );
INVx1_ASAP7_75t_L g581 ( .A(n_280), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_280), .A2(n_633), .B(n_634), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_281), .Y(n_1461) );
AO22x2_ASAP7_75t_L g873 ( .A1(n_282), .A2(n_874), .B1(n_875), .B2(n_944), .Y(n_873) );
INVx1_ASAP7_75t_L g944 ( .A(n_282), .Y(n_944) );
INVxp67_ASAP7_75t_L g1201 ( .A(n_283), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_284), .A2(n_332), .B1(n_425), .B2(n_426), .Y(n_1547) );
INVx1_ASAP7_75t_L g1564 ( .A(n_284), .Y(n_1564) );
INVx1_ASAP7_75t_L g1432 ( .A(n_288), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_289), .Y(n_900) );
AOI221xp5_ASAP7_75t_L g1533 ( .A1(n_290), .A2(n_316), .B1(n_1534), .B2(n_1535), .C(n_1536), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_291), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g1555 ( .A(n_293), .Y(n_1555) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_295), .Y(n_678) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_296), .Y(n_737) );
INVx1_ASAP7_75t_L g687 ( .A(n_297), .Y(n_687) );
INVx1_ASAP7_75t_L g1568 ( .A(n_298), .Y(n_1568) );
CKINVDCx5p33_ASAP7_75t_R g1312 ( .A(n_299), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g1933 ( .A(n_300), .Y(n_1933) );
INVx1_ASAP7_75t_L g1313 ( .A(n_301), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_302), .A2(n_335), .B1(n_1134), .B2(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1392 ( .A(n_302), .Y(n_1392) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_303), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_303), .A2(n_359), .B1(n_779), .B2(n_781), .Y(n_850) );
OAI221xp5_ASAP7_75t_SL g683 ( .A1(n_304), .A2(n_347), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_304), .A2(n_347), .B1(n_401), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_305), .A2(n_338), .B1(n_1228), .B2(n_1388), .Y(n_1405) );
INVx1_ASAP7_75t_L g1424 ( .A(n_305), .Y(n_1424) );
INVx1_ASAP7_75t_L g1322 ( .A(n_306), .Y(n_1322) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_307), .Y(n_865) );
INVx1_ASAP7_75t_L g1519 ( .A(n_308), .Y(n_1519) );
CKINVDCx5p33_ASAP7_75t_R g1466 ( .A(n_309), .Y(n_1466) );
INVx1_ASAP7_75t_L g1698 ( .A(n_310), .Y(n_1698) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_311), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g1303 ( .A(n_312), .Y(n_1303) );
INVx1_ASAP7_75t_L g484 ( .A(n_313), .Y(n_484) );
INVx1_ASAP7_75t_L g1361 ( .A(n_315), .Y(n_1361) );
OAI332xp33_ASAP7_75t_L g1501 ( .A1(n_316), .A2(n_587), .A3(n_1019), .B1(n_1502), .B2(n_1506), .B3(n_1509), .C1(n_1512), .C2(n_1515), .Y(n_1501) );
INVx1_ASAP7_75t_L g999 ( .A(n_317), .Y(n_999) );
CKINVDCx5p33_ASAP7_75t_R g1411 ( .A(n_319), .Y(n_1411) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_320), .Y(n_849) );
INVx1_ASAP7_75t_L g1482 ( .A(n_321), .Y(n_1482) );
XNOR2xp5_ASAP7_75t_L g1946 ( .A(n_323), .B(n_1882), .Y(n_1946) );
INVx1_ASAP7_75t_L g1507 ( .A(n_324), .Y(n_1507) );
INVx1_ASAP7_75t_L g1116 ( .A(n_325), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_326), .Y(n_368) );
AND3x2_ASAP7_75t_L g1649 ( .A(n_326), .B(n_366), .C(n_1650), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_326), .B(n_366), .Y(n_1658) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_327), .Y(n_1241) );
INVx2_ASAP7_75t_L g379 ( .A(n_328), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_330), .A2(n_471), .B(n_951), .C(n_954), .Y(n_950) );
INVx1_ASAP7_75t_L g986 ( .A(n_330), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1553 ( .A1(n_331), .A2(n_345), .B1(n_1024), .B2(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1574 ( .A(n_331), .Y(n_1574) );
INVx1_ASAP7_75t_L g1569 ( .A(n_332), .Y(n_1569) );
INVx1_ASAP7_75t_L g1373 ( .A(n_335), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_337), .Y(n_1246) );
INVx1_ASAP7_75t_L g1428 ( .A(n_338), .Y(n_1428) );
INVx1_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
INVx2_ASAP7_75t_L g466 ( .A(n_341), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g1245 ( .A(n_342), .Y(n_1245) );
INVx1_ASAP7_75t_L g531 ( .A(n_344), .Y(n_531) );
INVx1_ASAP7_75t_L g1579 ( .A(n_345), .Y(n_1579) );
INVx1_ASAP7_75t_L g1703 ( .A(n_346), .Y(n_1703) );
INVx1_ASAP7_75t_L g1059 ( .A(n_348), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g1558 ( .A(n_350), .Y(n_1558) );
AOI21xp33_ASAP7_75t_L g1299 ( .A1(n_351), .A2(n_413), .B(n_648), .Y(n_1299) );
INVx1_ASAP7_75t_L g1321 ( .A(n_351), .Y(n_1321) );
INVx1_ASAP7_75t_L g1478 ( .A(n_352), .Y(n_1478) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_353), .Y(n_1004) );
INVxp33_ASAP7_75t_SL g1889 ( .A(n_354), .Y(n_1889) );
INVx1_ASAP7_75t_L g1069 ( .A(n_355), .Y(n_1069) );
INVx1_ASAP7_75t_L g1331 ( .A(n_357), .Y(n_1331) );
INVx1_ASAP7_75t_L g1206 ( .A(n_358), .Y(n_1206) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_359), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_382), .B(n_1637), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_369), .Y(n_363) );
AND2x4_ASAP7_75t_L g1939 ( .A(n_364), .B(n_370), .Y(n_1939) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_SL g1944 ( .A(n_365), .Y(n_1944) );
NAND2xp5_ASAP7_75t_L g1949 ( .A(n_365), .B(n_367), .Y(n_1949) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g1943 ( .A(n_367), .B(n_1944), .Y(n_1943) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g499 ( .A(n_373), .B(n_381), .Y(n_499) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g588 ( .A(n_374), .B(n_589), .Y(n_588) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
BUFx2_ASAP7_75t_L g495 ( .A(n_376), .Y(n_495) );
INVx1_ASAP7_75t_L g513 ( .A(n_376), .Y(n_513) );
OR2x2_ASAP7_75t_L g614 ( .A(n_376), .B(n_598), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_376), .A2(n_509), .B1(n_678), .B2(n_679), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_376), .A2(n_509), .B1(n_695), .B2(n_696), .Y(n_694) );
INVx2_ASAP7_75t_SL g892 ( .A(n_376), .Y(n_892) );
BUFx6f_ASAP7_75t_L g1007 ( .A(n_376), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x4_ASAP7_75t_L g469 ( .A(n_378), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g475 ( .A(n_378), .Y(n_475) );
INVx2_ASAP7_75t_L g483 ( .A(n_378), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_378), .Y(n_491) );
AND2x2_ASAP7_75t_L g530 ( .A(n_378), .B(n_379), .Y(n_530) );
INVx2_ASAP7_75t_L g470 ( .A(n_379), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_379), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g490 ( .A(n_379), .Y(n_490) );
INVx1_ASAP7_75t_L g537 ( .A(n_379), .Y(n_537) );
INVx1_ASAP7_75t_L g548 ( .A(n_379), .Y(n_548) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_1054), .B2(n_1055), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
XNOR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_814), .Y(n_384) );
AO22x2_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_732), .B1(n_812), .B2(n_813), .Y(n_385) );
INVx1_ASAP7_75t_L g812 ( .A(n_386), .Y(n_812) );
XNOR2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_570), .Y(n_386) );
NAND4xp75_ASAP7_75t_L g388 ( .A(n_389), .B(n_459), .C(n_551), .D(n_560), .Y(n_388) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_390), .B(n_435), .Y(n_389) );
AOI33xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_399), .A3(n_411), .B1(n_423), .B2(n_424), .B3(n_429), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_392), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_392), .Y(n_926) );
INVx2_ASAP7_75t_L g1066 ( .A(n_392), .Y(n_1066) );
OR2x6_ASAP7_75t_L g392 ( .A(n_393), .B(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g1306 ( .A(n_393), .Y(n_1306) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g634 ( .A(n_394), .Y(n_634) );
BUFx3_ASAP7_75t_L g713 ( .A(n_394), .Y(n_713) );
INVx1_ASAP7_75t_L g861 ( .A(n_394), .Y(n_861) );
INVx1_ASAP7_75t_L g979 ( .A(n_394), .Y(n_979) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x4_ASAP7_75t_L g433 ( .A(n_395), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
AND2x2_ASAP7_75t_L g594 ( .A(n_397), .B(n_517), .Y(n_594) );
AND2x4_ASAP7_75t_L g674 ( .A(n_397), .B(n_499), .Y(n_674) );
INVx2_ASAP7_75t_L g727 ( .A(n_397), .Y(n_727) );
AND2x4_ASAP7_75t_L g755 ( .A(n_397), .B(n_499), .Y(n_755) );
BUFx2_ASAP7_75t_L g871 ( .A(n_397), .Y(n_871) );
OR2x2_ASAP7_75t_L g978 ( .A(n_397), .B(n_979), .Y(n_978) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g550 ( .A(n_398), .Y(n_550) );
OR2x6_ASAP7_75t_L g587 ( .A(n_398), .B(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx3_ASAP7_75t_L g425 ( .A(n_401), .Y(n_425) );
INVx1_ASAP7_75t_L g785 ( .A(n_401), .Y(n_785) );
INVx2_ASAP7_75t_L g1221 ( .A(n_401), .Y(n_1221) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g563 ( .A(n_402), .Y(n_563) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_402), .Y(n_619) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_402), .Y(n_633) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_402), .Y(n_777) );
BUFx3_ASAP7_75t_L g1087 ( .A(n_402), .Y(n_1087) );
BUFx2_ASAP7_75t_L g1228 ( .A(n_402), .Y(n_1228) );
BUFx2_ASAP7_75t_L g1626 ( .A(n_402), .Y(n_1626) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g569 ( .A(n_403), .Y(n_569) );
INVx2_ASAP7_75t_L g416 ( .A(n_404), .Y(n_416) );
AND2x2_ASAP7_75t_L g422 ( .A(n_404), .B(n_409), .Y(n_422) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x6_ASAP7_75t_L g557 ( .A(n_407), .B(n_554), .Y(n_557) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_407), .B(n_554), .Y(n_1173) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
INVx2_ASAP7_75t_L g622 ( .A(n_408), .Y(n_622) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_408), .Y(n_787) );
INVx1_ASAP7_75t_L g1223 ( .A(n_408), .Y(n_1223) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx2_ASAP7_75t_L g417 ( .A(n_409), .Y(n_417) );
INVx1_ASAP7_75t_L g568 ( .A(n_410), .Y(n_568) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g552 ( .A(n_413), .B(n_553), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_413), .A2(n_650), .B(n_651), .C(n_657), .Y(n_649) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g802 ( .A(n_414), .Y(n_802) );
INVx1_ASAP7_75t_L g1035 ( .A(n_414), .Y(n_1035) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g559 ( .A(n_415), .B(n_442), .Y(n_559) );
INVx6_ASAP7_75t_L g647 ( .A(n_415), .Y(n_647) );
BUFx2_ASAP7_75t_L g1387 ( .A(n_415), .Y(n_1387) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
INVx1_ASAP7_75t_L g452 ( .A(n_417), .Y(n_452) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g803 ( .A(n_420), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g1159 ( .A(n_420), .Y(n_1159) );
BUFx6f_ASAP7_75t_L g1229 ( .A(n_420), .Y(n_1229) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_421), .Y(n_721) );
INVx2_ASAP7_75t_L g1298 ( .A(n_421), .Y(n_1298) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_422), .Y(n_628) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g702 ( .A(n_428), .Y(n_702) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_428), .Y(n_723) );
BUFx6f_ASAP7_75t_L g1024 ( .A(n_428), .Y(n_1024) );
INVx1_ASAP7_75t_L g1167 ( .A(n_428), .Y(n_1167) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g977 ( .A1(n_430), .A2(n_978), .B1(n_980), .B2(n_984), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g1064 ( .A1(n_430), .A2(n_1065), .B1(n_1067), .B2(n_1079), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_430), .A2(n_1065), .B1(n_1244), .B2(n_1252), .Y(n_1243) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx4f_ASAP7_75t_L g940 ( .A(n_431), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_431), .A2(n_1066), .B1(n_1157), .B2(n_1161), .C(n_1168), .Y(n_1156) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AND2x4_ASAP7_75t_L g558 ( .A(n_432), .B(n_559), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_433), .Y(n_648) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_433), .Y(n_791) );
INVx2_ASAP7_75t_L g856 ( .A(n_433), .Y(n_856) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_433), .Y(n_1036) );
INVx1_ASAP7_75t_L g1536 ( .A(n_433), .Y(n_1536) );
OAI221xp5_ASAP7_75t_L g1918 ( .A1(n_433), .A2(n_1080), .B1(n_1888), .B2(n_1919), .C(n_1920), .Y(n_1918) );
AND2x4_ASAP7_75t_L g442 ( .A(n_434), .B(n_443), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_447), .B1(n_448), .B2(n_454), .C(n_455), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_436), .A2(n_909), .B1(n_911), .B2(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
OR2x2_ASAP7_75t_L g781 ( .A(n_438), .B(n_782), .Y(n_781) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_438), .B(n_441), .Y(n_1091) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_439), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
AND2x4_ASAP7_75t_L g706 ( .A(n_439), .B(n_442), .Y(n_706) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_439), .B(n_442), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_439), .B(n_442), .Y(n_1458) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g453 ( .A(n_441), .Y(n_453) );
INVx1_ASAP7_75t_L g458 ( .A(n_441), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .Y(n_441) );
BUFx2_ASAP7_75t_L g658 ( .A(n_442), .Y(n_658) );
AND2x4_ASAP7_75t_L g705 ( .A(n_442), .B(n_654), .Y(n_705) );
AND2x4_ASAP7_75t_L g780 ( .A(n_442), .B(n_654), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_442), .Y(n_782) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x6_ASAP7_75t_L g767 ( .A(n_445), .B(n_518), .Y(n_767) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g554 ( .A(n_446), .B(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g577 ( .A(n_446), .B(n_465), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_447), .A2(n_454), .B1(n_535), .B2(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g924 ( .A(n_449), .Y(n_924) );
INVx2_ASAP7_75t_L g1258 ( .A(n_449), .Y(n_1258) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g654 ( .A(n_451), .Y(n_654) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g975 ( .A(n_455), .B(n_976), .C(n_977), .Y(n_975) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_455), .Y(n_1088) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_458), .B(n_798), .Y(n_943) );
OAI31xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_476), .A3(n_540), .B(n_549), .Y(n_459) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g879 ( .A(n_462), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_462), .A2(n_545), .B1(n_952), .B2(n_953), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_462), .A2(n_545), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
AND2x4_ASAP7_75t_L g472 ( .A(n_463), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g542 ( .A(n_465), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g545 ( .A(n_465), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g519 ( .A(n_466), .Y(n_519) );
INVx1_ASAP7_75t_L g589 ( .A(n_466), .Y(n_589) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g592 ( .A(n_468), .Y(n_592) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_469), .Y(n_486) );
INVx3_ASAP7_75t_L g506 ( .A(n_469), .Y(n_506) );
AND2x4_ASAP7_75t_L g474 ( .A(n_470), .B(n_475), .Y(n_474) );
INVx8_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_473), .Y(n_837) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_474), .Y(n_586) );
BUFx3_ASAP7_75t_L g601 ( .A(n_474), .Y(n_601) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_474), .Y(n_609) );
BUFx2_ASAP7_75t_L g672 ( .A(n_474), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_487), .B1(n_500), .B2(n_508), .C(n_521), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_484), .B2(n_485), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g501 ( .A(n_480), .Y(n_501) );
INVx2_ASAP7_75t_L g1504 ( .A(n_480), .Y(n_1504) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g684 ( .A(n_481), .Y(n_684) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g580 ( .A(n_482), .Y(n_580) );
BUFx2_ASAP7_75t_L g965 ( .A(n_482), .Y(n_965) );
INVx1_ASAP7_75t_L g539 ( .A(n_483), .Y(n_539) );
AND2x4_ASAP7_75t_L g546 ( .A(n_483), .B(n_547), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_485), .A2(n_1011), .B1(n_1012), .B2(n_1014), .Y(n_1010) );
OAI221xp5_ASAP7_75t_L g1106 ( .A1(n_485), .A2(n_882), .B1(n_1107), .B2(n_1108), .C(n_1109), .Y(n_1106) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g763 ( .A(n_486), .Y(n_763) );
INVx4_ASAP7_75t_L g840 ( .A(n_486), .Y(n_840) );
INVx2_ASAP7_75t_SL g885 ( .A(n_486), .Y(n_885) );
BUFx3_ASAP7_75t_L g1581 ( .A(n_486), .Y(n_1581) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_492), .B1(n_493), .B2(n_496), .C(n_497), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g1151 ( .A1(n_488), .A2(n_1152), .B(n_1153), .Y(n_1151) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g533 ( .A(n_489), .Y(n_533) );
BUFx2_ASAP7_75t_L g889 ( .A(n_489), .Y(n_889) );
INVx2_ASAP7_75t_L g896 ( .A(n_489), .Y(n_896) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_490), .B(n_491), .Y(n_510) );
INVx1_ASAP7_75t_L g669 ( .A(n_491), .Y(n_669) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g1333 ( .A(n_494), .Y(n_1333) );
INVx2_ASAP7_75t_SL g1337 ( .A(n_494), .Y(n_1337) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g1095 ( .A1(n_497), .A2(n_891), .B1(n_1069), .B2(n_1073), .C(n_1096), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_497), .A2(n_891), .B1(n_1245), .B2(n_1246), .C(n_1272), .Y(n_1271) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_SL g894 ( .A(n_499), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_503), .B2(n_507), .Y(n_500) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_501), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_511), .B1(n_561), .B2(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g956 ( .A(n_505), .Y(n_956) );
INVx3_ASAP7_75t_L g1203 ( .A(n_505), .Y(n_1203) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g583 ( .A(n_506), .Y(n_583) );
INVx3_ASAP7_75t_L g613 ( .A(n_506), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g551 ( .A1(n_507), .A2(n_514), .B1(n_531), .B2(n_552), .C1(n_556), .C2(n_558), .Y(n_551) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_511), .B1(n_512), .B2(n_514), .C(n_515), .Y(n_508) );
BUFx3_ASAP7_75t_L g1005 ( .A(n_509), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_509), .A2(n_1007), .B1(n_1008), .B2(n_1009), .Y(n_1006) );
BUFx3_ASAP7_75t_L g1197 ( .A(n_509), .Y(n_1197) );
INVx2_ASAP7_75t_L g1273 ( .A(n_509), .Y(n_1273) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g1512 ( .A1(n_512), .A2(n_1433), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g901 ( .A(n_513), .Y(n_901) );
INVx1_ASAP7_75t_L g1575 ( .A(n_513), .Y(n_1575) );
INVx1_ASAP7_75t_L g1898 ( .A(n_513), .Y(n_1898) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_515), .A2(n_899), .B1(n_900), .B2(n_901), .C(n_902), .Y(n_898) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g1112 ( .A(n_517), .Y(n_1112) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_531), .B(n_532), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp67_ASAP7_75t_L g917 ( .A(n_523), .B(n_727), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
AND2x2_ASAP7_75t_L g910 ( .A(n_524), .B(n_665), .Y(n_910) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_524), .B(n_665), .Y(n_1115) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI21xp33_ASAP7_75t_L g532 ( .A1(n_525), .A2(n_533), .B(n_534), .Y(n_532) );
OR2x6_ASAP7_75t_L g895 ( .A(n_525), .B(n_896), .Y(n_895) );
OR2x6_ASAP7_75t_L g913 ( .A(n_525), .B(n_539), .Y(n_913) );
INVx1_ASAP7_75t_L g961 ( .A(n_525), .Y(n_961) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_525), .B(n_896), .Y(n_1104) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g576 ( .A(n_528), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g688 ( .A(n_529), .Y(n_688) );
INVx2_ASAP7_75t_L g1349 ( .A(n_529), .Y(n_1349) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_530), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_533), .A2(n_891), .B1(n_894), .B2(n_970), .C(n_971), .Y(n_969) );
BUFx2_ASAP7_75t_L g1096 ( .A(n_533), .Y(n_1096) );
NAND2x1_ASAP7_75t_SL g596 ( .A(n_535), .B(n_597), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g960 ( .A(n_535), .B(n_961), .Y(n_960) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_538), .B(n_597), .Y(n_599) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
CKINVDCx6p67_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g958 ( .A(n_543), .Y(n_958) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g878 ( .A(n_545), .Y(n_878) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_546), .Y(n_606) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_546), .Y(n_676) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_546), .Y(n_691) );
INVx1_ASAP7_75t_L g1135 ( .A(n_546), .Y(n_1135) );
INVx1_ASAP7_75t_L g1352 ( .A(n_546), .Y(n_1352) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g659 ( .A(n_549), .Y(n_659) );
BUFx8_ASAP7_75t_SL g972 ( .A(n_549), .Y(n_972) );
AOI31xp33_ASAP7_75t_L g1614 ( .A1(n_549), .A2(n_1615), .A3(n_1623), .B(n_1632), .Y(n_1614) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g811 ( .A(n_550), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_552), .A2(n_561), .B1(n_902), .B2(n_906), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_552), .A2(n_561), .B1(n_989), .B2(n_990), .C(n_991), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_552), .A2(n_561), .B1(n_1170), .B2(n_1171), .C(n_1172), .Y(n_1169) );
AND2x2_ASAP7_75t_L g561 ( .A(n_553), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x6_ASAP7_75t_L g565 ( .A(n_554), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_554), .B(n_1122), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_554), .B(n_1124), .Y(n_1123) );
INVx2_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_555), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g624 ( .A(n_555), .B(n_625), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g1022 ( .A1(n_555), .A2(n_1023), .B(n_1025), .C(n_1027), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_556), .A2(n_564), .B1(n_900), .B2(n_907), .Y(n_920) );
CKINVDCx6p67_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g771 ( .A(n_558), .Y(n_771) );
OR2x6_ASAP7_75t_L g916 ( .A(n_558), .B(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g725 ( .A(n_559), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_559), .B(n_1046), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_562), .A2(n_1009), .B1(n_1011), .B2(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g709 ( .A(n_563), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_563), .A2(n_702), .B1(n_1149), .B2(n_1150), .Y(n_1160) );
INVx2_ASAP7_75t_SL g1248 ( .A(n_563), .Y(n_1248) );
CKINVDCx6p67_ASAP7_75t_R g564 ( .A(n_565), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_566), .A2(n_631), .B(n_632), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_566), .A2(n_745), .B1(n_748), .B2(n_789), .C(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g1083 ( .A(n_566), .Y(n_1083) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g643 ( .A(n_567), .Y(n_643) );
INVx1_ASAP7_75t_L g652 ( .A(n_567), .Y(n_652) );
BUFx2_ASAP7_75t_L g854 ( .A(n_567), .Y(n_854) );
BUFx4f_ASAP7_75t_L g982 ( .A(n_567), .Y(n_982) );
INVx1_ASAP7_75t_L g1072 ( .A(n_567), .Y(n_1072) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OR2x2_ASAP7_75t_L g625 ( .A(n_568), .B(n_569), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_660), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_602), .C(n_615), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_595), .Y(n_573) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g605 ( .A(n_577), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_577), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g612 ( .A(n_577), .B(n_613), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_577), .A2(n_594), .B1(n_683), .B2(n_690), .Y(n_682) );
AND2x4_ASAP7_75t_L g744 ( .A(n_577), .B(n_583), .Y(n_744) );
AND2x6_ASAP7_75t_L g746 ( .A(n_577), .B(n_601), .Y(n_746) );
AND2x4_ASAP7_75t_L g749 ( .A(n_577), .B(n_688), .Y(n_749) );
AND2x2_ASAP7_75t_L g751 ( .A(n_577), .B(n_606), .Y(n_751) );
AND2x2_ASAP7_75t_L g833 ( .A(n_577), .B(n_606), .Y(n_833) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_577), .B(n_606), .Y(n_1367) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B1(n_582), .B2(n_584), .C(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g905 ( .A(n_579), .Y(n_905) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g1013 ( .A(n_580), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_580), .Y(n_1148) );
INVx2_ASAP7_75t_L g1262 ( .A(n_580), .Y(n_1262) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g685 ( .A(n_583), .Y(n_685) );
INVx1_ASAP7_75t_L g967 ( .A(n_583), .Y(n_967) );
BUFx3_ASAP7_75t_L g1208 ( .A(n_583), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_584), .A2(n_636), .B1(n_637), .B2(n_639), .Y(n_635) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_586), .Y(n_1140) );
BUFx2_ASAP7_75t_L g1359 ( .A(n_586), .Y(n_1359) );
INVx1_ASAP7_75t_L g1193 ( .A(n_587), .Y(n_1193) );
OAI33xp33_ASAP7_75t_L g1326 ( .A1(n_587), .A2(n_1212), .A3(n_1327), .B1(n_1332), .B2(n_1336), .B3(n_1338), .Y(n_1326) );
OAI33xp33_ASAP7_75t_L g1430 ( .A1(n_587), .A2(n_767), .A3(n_1431), .B1(n_1435), .B2(n_1439), .B3(n_1441), .Y(n_1430) );
OAI33xp33_ASAP7_75t_L g1476 ( .A1(n_587), .A2(n_1212), .A3(n_1477), .B1(n_1481), .B2(n_1487), .B3(n_1488), .Y(n_1476) );
OAI33xp33_ASAP7_75t_L g1572 ( .A1(n_587), .A2(n_1515), .A3(n_1573), .B1(n_1577), .B2(n_1582), .B3(n_1583), .Y(n_1572) );
HB1xp67_ASAP7_75t_L g1895 ( .A(n_587), .Y(n_1895) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .C(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g1330 ( .A(n_592), .Y(n_1330) );
HB1xp67_ASAP7_75t_L g1353 ( .A(n_592), .Y(n_1353) );
INVx2_ASAP7_75t_L g1188 ( .A(n_596), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1324 ( .A(n_596), .Y(n_1324) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_597), .B(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g664 ( .A(n_597), .B(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g667 ( .A(n_597), .B(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g671 ( .A(n_597), .B(n_672), .Y(n_671) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx4f_ASAP7_75t_L g1189 ( .A(n_599), .Y(n_1189) );
BUFx4f_ASAP7_75t_L g1325 ( .A(n_599), .Y(n_1325) );
BUFx3_ASAP7_75t_L g1190 ( .A(n_600), .Y(n_1190) );
BUFx2_ASAP7_75t_L g1475 ( .A(n_600), .Y(n_1475) );
BUFx2_ASAP7_75t_L g1571 ( .A(n_600), .Y(n_1571) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_601), .Y(n_1266) );
NOR2xp33_ASAP7_75t_SL g602 ( .A(n_603), .B(n_610), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g1018 ( .A(n_605), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_605), .A2(n_749), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1500 ( .A(n_605), .Y(n_1500) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g1019 ( .A(n_608), .Y(n_1019) );
INVx2_ASAP7_75t_SL g759 ( .A(n_609), .Y(n_759) );
BUFx6f_ASAP7_75t_L g843 ( .A(n_609), .Y(n_843) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g693 ( .A(n_613), .Y(n_693) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_613), .Y(n_1001) );
INVx1_ASAP7_75t_L g1102 ( .A(n_613), .Y(n_1102) );
INVx2_ASAP7_75t_L g1485 ( .A(n_613), .Y(n_1485) );
INVx2_ASAP7_75t_L g681 ( .A(n_614), .Y(n_681) );
AND2x4_ASAP7_75t_L g770 ( .A(n_614), .B(n_771), .Y(n_770) );
OAI31xp33_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_623), .A3(n_629), .B(n_659), .Y(n_615) );
INVx1_ASAP7_75t_L g1372 ( .A(n_617), .Y(n_1372) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_619), .A2(n_628), .B1(n_696), .B2(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g1124 ( .A(n_619), .Y(n_1124) );
BUFx4f_ASAP7_75t_L g1164 ( .A(n_619), .Y(n_1164) );
AND2x4_ASAP7_75t_L g627 ( .A(n_620), .B(n_628), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_620), .A2(n_666), .B1(n_670), .B2(n_699), .C1(n_705), .C2(n_706), .Y(n_698) );
AND2x4_ASAP7_75t_L g776 ( .A(n_620), .B(n_777), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_620), .A2(n_627), .B1(n_717), .B2(n_1514), .C(n_1524), .Y(n_1523) );
INVx4_ASAP7_75t_L g809 ( .A(n_621), .Y(n_809) );
INVx1_ASAP7_75t_L g640 ( .A(n_622), .Y(n_640) );
INVx2_ASAP7_75t_L g1251 ( .A(n_622), .Y(n_1251) );
INVx6_ASAP7_75t_L g807 ( .A(n_624), .Y(n_807) );
INVx1_ASAP7_75t_L g638 ( .A(n_625), .Y(n_638) );
INVx1_ASAP7_75t_L g701 ( .A(n_625), .Y(n_701) );
INVx2_ASAP7_75t_L g790 ( .A(n_625), .Y(n_790) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_625), .Y(n_1068) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_627), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g1302 ( .A1(n_627), .A2(n_717), .B1(n_1303), .B2(n_1304), .C(n_1307), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_627), .Y(n_1382) );
HB1xp67_ASAP7_75t_L g1410 ( .A(n_627), .Y(n_1410) );
AOI221xp5_ASAP7_75t_L g1447 ( .A1(n_627), .A2(n_717), .B1(n_1448), .B2(n_1449), .C(n_1450), .Y(n_1447) );
INVx2_ASAP7_75t_SL g711 ( .A(n_628), .Y(n_711) );
AND2x4_ASAP7_75t_L g717 ( .A(n_628), .B(n_658), .Y(n_717) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_628), .Y(n_798) );
INVx1_ASAP7_75t_L g860 ( .A(n_628), .Y(n_860) );
BUFx3_ASAP7_75t_L g935 ( .A(n_628), .Y(n_935) );
BUFx4f_ASAP7_75t_L g1026 ( .A(n_628), .Y(n_1026) );
INVx1_ASAP7_75t_L g1414 ( .A(n_628), .Y(n_1414) );
OAI211xp5_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_635), .B(n_641), .C(n_649), .Y(n_629) );
BUFx3_ASAP7_75t_L g1529 ( .A(n_633), .Y(n_1529) );
INVx1_ASAP7_75t_L g800 ( .A(n_634), .Y(n_800) );
BUFx2_ASAP7_75t_L g1927 ( .A(n_634), .Y(n_1927) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_637), .A2(n_829), .B1(n_831), .B2(n_853), .C(n_855), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g984 ( .A1(n_637), .A2(n_981), .B1(n_985), .B2(n_986), .C(n_987), .Y(n_984) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B(n_644), .C(n_645), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g1224 ( .A1(n_643), .A2(n_789), .B1(n_1182), .B2(n_1184), .C(n_1225), .Y(n_1224) );
OAI211xp5_ASAP7_75t_L g1377 ( .A1(n_643), .A2(n_1363), .B(n_1378), .C(n_1379), .Y(n_1377) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_646), .Y(n_715) );
INVx1_ASAP7_75t_L g934 ( .A(n_646), .Y(n_934) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g720 ( .A(n_647), .Y(n_720) );
INVx1_ASAP7_75t_L g864 ( .A(n_647), .Y(n_864) );
BUFx6f_ASAP7_75t_L g1233 ( .A(n_647), .Y(n_1233) );
INVx2_ASAP7_75t_SL g1380 ( .A(n_647), .Y(n_1380) );
INVx1_ASAP7_75t_L g1535 ( .A(n_647), .Y(n_1535) );
NAND2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g1032 ( .A(n_652), .Y(n_1032) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g1543 ( .A1(n_659), .A2(n_1544), .B1(n_1559), .B2(n_1560), .Y(n_1543) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_661), .B(n_728), .Y(n_660) );
INVx1_ASAP7_75t_L g730 ( .A(n_662), .Y(n_730) );
NAND3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_673), .C(n_682), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B1(n_667), .B2(n_670), .C(n_671), .Y(n_663) );
INVx1_ASAP7_75t_L g739 ( .A(n_664), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_664), .A2(n_821), .B1(n_823), .B2(n_824), .C(n_825), .Y(n_820) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_664), .A2(n_667), .B1(n_671), .B2(n_1048), .C(n_1049), .Y(n_1047) );
AOI221xp5_ASAP7_75t_L g1343 ( .A1(n_664), .A2(n_667), .B1(n_671), .B2(n_1344), .C(n_1345), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g1540 ( .A1(n_664), .A2(n_671), .B(n_1521), .Y(n_1540) );
AOI221xp5_ASAP7_75t_L g1590 ( .A1(n_664), .A2(n_667), .B1(n_671), .B2(n_1591), .C(n_1592), .Y(n_1590) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_667), .Y(n_736) );
INVx1_ASAP7_75t_L g822 ( .A(n_667), .Y(n_822) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_671), .A2(n_736), .B1(n_737), .B2(n_738), .C(n_740), .Y(n_735) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_671), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_672), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
HB1xp67_ASAP7_75t_L g1608 ( .A(n_672), .Y(n_1608) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_680), .B2(n_681), .Y(n_673) );
BUFx2_ASAP7_75t_L g1347 ( .A(n_674), .Y(n_1347) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_680), .A2(n_719), .B1(n_722), .B2(n_724), .Y(n_718) );
INVx2_ASAP7_75t_L g883 ( .A(n_684), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_685), .A2(n_1147), .B1(n_1149), .B2(n_1150), .Y(n_1146) );
INVx1_ASAP7_75t_L g1355 ( .A(n_685), .Y(n_1355) );
BUFx3_ASAP7_75t_L g757 ( .A(n_688), .Y(n_757) );
INVx1_ASAP7_75t_L g1138 ( .A(n_688), .Y(n_1138) );
INVx1_ASAP7_75t_L g1358 ( .A(n_688), .Y(n_1358) );
BUFx3_ASAP7_75t_L g761 ( .A(n_691), .Y(n_761) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g729 ( .A(n_697), .Y(n_729) );
AOI31xp33_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_707), .A3(n_718), .B(n_726), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g1525 ( .A1(n_700), .A2(n_1167), .B1(n_1505), .B2(n_1508), .C(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g716 ( .A(n_702), .Y(n_716) );
INVx4_ASAP7_75t_L g1375 ( .A(n_705), .Y(n_1375) );
INVx2_ASAP7_75t_L g1408 ( .A(n_705), .Y(n_1408) );
AOI322xp5_ASAP7_75t_L g1294 ( .A1(n_706), .A2(n_780), .A3(n_1295), .B1(n_1296), .B2(n_1299), .C1(n_1300), .C2(n_1301), .Y(n_1294) );
INVx2_ASAP7_75t_SL g1376 ( .A(n_706), .Y(n_1376) );
INVx2_ASAP7_75t_L g1407 ( .A(n_706), .Y(n_1407) );
AOI222xp33_ASAP7_75t_SL g1518 ( .A1(n_706), .A2(n_724), .B1(n_1519), .B2(n_1520), .C1(n_1521), .C2(n_1522), .Y(n_1518) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_714), .B(n_717), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g931 ( .A(n_711), .Y(n_931) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g1230 ( .A(n_713), .Y(n_1230) );
INVx3_ASAP7_75t_L g1415 ( .A(n_713), .Y(n_1415) );
INVx1_ASAP7_75t_L g1027 ( .A(n_717), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_717), .A2(n_1382), .B1(n_1383), .B2(n_1384), .C(n_1386), .Y(n_1381) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_717), .A2(n_1410), .B1(n_1411), .B2(n_1412), .C(n_1416), .Y(n_1409) );
AOI221xp5_ASAP7_75t_L g1551 ( .A1(n_717), .A2(n_793), .B1(n_1552), .B2(n_1553), .C(n_1555), .Y(n_1551) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_720), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_720), .A2(n_1008), .B1(n_1014), .B2(n_1024), .Y(n_1023) );
BUFx3_ASAP7_75t_L g1554 ( .A(n_720), .Y(n_1554) );
INVx1_ASAP7_75t_L g1078 ( .A(n_723), .Y(n_1078) );
INVx1_ASAP7_75t_L g1462 ( .A(n_723), .Y(n_1462) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI31xp33_ASAP7_75t_SL g1092 ( .A1(n_726), .A2(n_1093), .A3(n_1094), .B(n_1105), .Y(n_1092) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_731), .Y(n_728) );
INVx2_ASAP7_75t_L g813 ( .A(n_732), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_768), .Y(n_733) );
AND4x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_741), .C(n_747), .D(n_752), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_745), .B2(n_746), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_743), .A2(n_746), .B1(n_1463), .B2(n_1471), .Y(n_1470) );
BUFx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
BUFx2_ASAP7_75t_L g828 ( .A(n_744), .Y(n_828) );
BUFx2_ASAP7_75t_L g1181 ( .A(n_744), .Y(n_1181) );
BUFx2_ASAP7_75t_L g1362 ( .A(n_744), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_744), .A2(n_746), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
BUFx2_ASAP7_75t_L g1565 ( .A(n_744), .Y(n_1565) );
BUFx2_ASAP7_75t_L g1601 ( .A(n_744), .Y(n_1601) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_746), .A2(n_827), .B1(n_828), .B2(n_829), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_746), .A2(n_1180), .B1(n_1181), .B2(n_1182), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_746), .A2(n_1181), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_746), .A2(n_1361), .B1(n_1362), .B2(n_1363), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_746), .A2(n_1564), .B1(n_1565), .B2(n_1566), .Y(n_1563) );
BUFx2_ASAP7_75t_L g1596 ( .A(n_746), .Y(n_1596) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_749), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_749), .A2(n_833), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_749), .A2(n_1365), .B1(n_1366), .B2(n_1367), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_749), .A2(n_751), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_749), .A2(n_833), .B1(n_1461), .B2(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1538 ( .A(n_749), .Y(n_1538) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_749), .A2(n_1367), .B1(n_1568), .B2(n_1569), .Y(n_1567) );
BUFx2_ASAP7_75t_L g1599 ( .A(n_749), .Y(n_1599) );
AOI33xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .A3(n_760), .B1(n_764), .B2(n_765), .B3(n_766), .Y(n_752) );
AOI33xp33_ASAP7_75t_L g834 ( .A1(n_753), .A2(n_766), .A3(n_835), .B1(n_838), .B2(n_841), .B3(n_842), .Y(n_834) );
AOI33xp33_ASAP7_75t_L g1602 ( .A1(n_753), .A2(n_1603), .A3(n_1607), .B1(n_1609), .B2(n_1610), .B3(n_1611), .Y(n_1602) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_763), .A2(n_904), .B1(n_906), .B2(n_907), .Y(n_903) );
INVx1_ASAP7_75t_L g1015 ( .A(n_766), .Y(n_1015) );
AOI33xp33_ASAP7_75t_L g1346 ( .A1(n_766), .A2(n_1347), .A3(n_1348), .B1(n_1350), .B2(n_1354), .B3(n_1356), .Y(n_1346) );
INVx2_ASAP7_75t_L g1515 ( .A(n_766), .Y(n_1515) );
INVx6_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx5_ASAP7_75t_L g1213 ( .A(n_767), .Y(n_1213) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_772), .B(n_773), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_769), .A2(n_811), .B1(n_1215), .B2(n_1235), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_769), .A2(n_1369), .B1(n_1446), .B2(n_1467), .Y(n_1445) );
INVx1_ASAP7_75t_L g1935 ( .A(n_769), .Y(n_1935) );
INVx5_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g845 ( .A(n_770), .Y(n_845) );
INVx2_ASAP7_75t_SL g1314 ( .A(n_770), .Y(n_1314) );
INVx2_ASAP7_75t_L g1394 ( .A(n_770), .Y(n_1394) );
INVx1_ASAP7_75t_L g1560 ( .A(n_770), .Y(n_1560) );
AOI31xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_792), .A3(n_805), .B(n_810), .Y(n_773) );
AOI211xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_778), .C(n_783), .Y(n_774) );
AOI211xp5_ASAP7_75t_L g848 ( .A1(n_776), .A2(n_849), .B(n_850), .C(n_851), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_776), .A2(n_807), .B1(n_1205), .B2(n_1210), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_776), .B(n_1312), .Y(n_1311) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_776), .A2(n_1402), .B1(n_1403), .B2(n_1405), .C(n_1406), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_776), .B(n_1466), .Y(n_1465) );
AOI221xp5_ASAP7_75t_L g1545 ( .A1(n_776), .A2(n_1546), .B1(n_1547), .B2(n_1548), .C(n_1549), .Y(n_1545) );
AOI211xp5_ASAP7_75t_L g1615 ( .A1(n_776), .A2(n_1616), .B(n_1617), .C(n_1619), .Y(n_1615) );
HB1xp67_ASAP7_75t_L g1913 ( .A(n_776), .Y(n_1913) );
BUFx3_ASAP7_75t_L g937 ( .A(n_777), .Y(n_937) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_777), .Y(n_1076) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_SL g1042 ( .A(n_780), .Y(n_1042) );
INVx1_ASAP7_75t_L g1218 ( .A(n_780), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_780), .A2(n_1456), .B1(n_1457), .B2(n_1458), .Y(n_1455) );
INVx1_ASAP7_75t_L g1550 ( .A(n_780), .Y(n_1550) );
INVx2_ASAP7_75t_SL g1618 ( .A(n_780), .Y(n_1618) );
INVx1_ASAP7_75t_SL g804 ( .A(n_782), .Y(n_804) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_787), .Y(n_928) );
INVx1_ASAP7_75t_L g939 ( .A(n_787), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_789), .A2(n_970), .B1(n_971), .B2(n_981), .C(n_983), .Y(n_980) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g1080 ( .A(n_790), .Y(n_1080) );
INVx1_ASAP7_75t_L g1122 ( .A(n_790), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_801), .C(n_803), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_793), .A2(n_803), .B1(n_858), .B2(n_862), .C(n_865), .Y(n_857) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_793), .A2(n_803), .B1(n_1211), .B2(n_1227), .C(n_1231), .Y(n_1226) );
INVx1_ASAP7_75t_L g1923 ( .A(n_793), .Y(n_1923) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g1623 ( .A1(n_803), .A2(n_1410), .B1(n_1624), .B2(n_1625), .C(n_1629), .Y(n_1623) );
INVx1_ASAP7_75t_L g1931 ( .A(n_803), .Y(n_1931) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_807), .A2(n_809), .B1(n_867), .B2(n_868), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_807), .A2(n_809), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_807), .A2(n_809), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_807), .A2(n_809), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_807), .A2(n_809), .B1(n_1453), .B2(n_1454), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_807), .A2(n_809), .B1(n_1557), .B2(n_1558), .Y(n_1556) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_807), .A2(n_809), .B1(n_1633), .B2(n_1634), .Y(n_1632) );
AOI22xp33_ASAP7_75t_L g1932 ( .A1(n_807), .A2(n_809), .B1(n_1904), .B2(n_1907), .Y(n_1932) );
AOI211xp5_ASAP7_75t_L g1216 ( .A1(n_809), .A2(n_1206), .B(n_1217), .C(n_1219), .Y(n_1216) );
INVx1_ASAP7_75t_L g1369 ( .A(n_810), .Y(n_1369) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI31xp33_ASAP7_75t_L g1021 ( .A1(n_811), .A2(n_1022), .A3(n_1028), .B(n_1041), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_945), .B1(n_1052), .B2(n_1053), .Y(n_814) );
INVx1_ASAP7_75t_L g1052 ( .A(n_815), .Y(n_1052) );
XNOR2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_873), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_844), .Y(n_818) );
AND4x1_ASAP7_75t_L g819 ( .A(n_820), .B(n_826), .C(n_830), .D(n_834), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_840), .A2(n_1262), .B1(n_1263), .B2(n_1264), .C(n_1265), .Y(n_1261) );
OAI22xp33_ASAP7_75t_L g1502 ( .A1(n_840), .A2(n_1503), .B1(n_1504), .B2(n_1505), .Y(n_1502) );
AOI21xp33_ASAP7_75t_SL g844 ( .A1(n_845), .A2(n_846), .B(n_847), .Y(n_844) );
AOI31xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_857), .A3(n_866), .B(n_869), .Y(n_847) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_SL g1919 ( .A(n_854), .Y(n_1919) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g1534 ( .A(n_860), .Y(n_1534) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g1292 ( .A1(n_870), .A2(n_1293), .B1(n_1313), .B2(n_1314), .Y(n_1292) );
CKINVDCx8_ASAP7_75t_R g870 ( .A(n_871), .Y(n_870) );
OAI31xp33_ASAP7_75t_L g876 ( .A1(n_871), .A2(n_877), .A3(n_880), .B(n_897), .Y(n_876) );
OAI21xp5_ASAP7_75t_SL g1130 ( .A1(n_871), .A2(n_1131), .B(n_1145), .Y(n_1130) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND3xp33_ASAP7_75t_SL g875 ( .A(n_876), .B(n_914), .C(n_918), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_881) );
OAI22xp5_ASAP7_75t_SL g1577 ( .A1(n_882), .A2(n_1578), .B1(n_1579), .B2(n_1580), .Y(n_1577) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g1200 ( .A(n_883), .Y(n_1200) );
INVx2_ASAP7_75t_L g1436 ( .A(n_883), .Y(n_1436) );
INVx1_ASAP7_75t_L g1440 ( .A(n_883), .Y(n_1440) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_890), .B1(n_891), .B2(n_893), .C(n_894), .Y(n_887) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_888), .A2(n_1303), .B1(n_1309), .B2(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g899 ( .A(n_889), .Y(n_899) );
INVx1_ASAP7_75t_L g1479 ( .A(n_889), .Y(n_1479) );
OAI22xp33_ASAP7_75t_L g1002 ( .A1(n_891), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_891), .A2(n_1195), .B1(n_1196), .B2(n_1197), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g1209 ( .A1(n_891), .A2(n_1197), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
OAI22xp33_ASAP7_75t_L g1506 ( .A1(n_891), .A2(n_896), .B1(n_1507), .B2(n_1508), .Y(n_1506) );
INVx3_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
OAI22xp33_ASAP7_75t_L g1441 ( .A1(n_896), .A2(n_1337), .B1(n_1411), .B2(n_1418), .Y(n_1441) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_904), .A2(n_1205), .B1(n_1206), .B2(n_1207), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1582 ( .A1(n_904), .A2(n_1202), .B1(n_1548), .B2(n_1558), .Y(n_1582) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B1(n_911), .B2(n_912), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_912), .A2(n_1114), .B1(n_1116), .B2(n_1117), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_912), .A2(n_1114), .B1(n_1268), .B2(n_1269), .Y(n_1267) );
CKINVDCx11_ASAP7_75t_R g912 ( .A(n_913), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_916), .B(n_974), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_916), .B(n_1062), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_916), .B(n_1155), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_916), .B(n_1241), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_922), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
NAND3xp33_ASAP7_75t_SL g922 ( .A(n_923), .B(n_925), .C(n_941), .Y(n_922) );
INVx1_ASAP7_75t_L g1090 ( .A(n_924), .Y(n_1090) );
AOI33xp33_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .A3(n_929), .B1(n_932), .B2(n_936), .B3(n_940), .Y(n_925) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g1702 ( .A1(n_944), .A2(n_1656), .B1(n_1663), .B2(n_1703), .Y(n_1702) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_946), .Y(n_1053) );
XNOR2x1_ASAP7_75t_L g946 ( .A(n_947), .B(n_994), .Y(n_946) );
INVx1_ASAP7_75t_L g992 ( .A(n_948), .Y(n_992) );
NAND4xp25_ASAP7_75t_L g948 ( .A(n_949), .B(n_973), .C(n_975), .D(n_988), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_962), .B(n_972), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_957), .B(n_959), .Y(n_954) );
INVx1_ASAP7_75t_L g1111 ( .A(n_958), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_964), .A2(n_998), .B1(n_999), .B2(n_1000), .Y(n_997) );
BUFx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g1276 ( .A(n_965), .Y(n_1276) );
INVx5_ASAP7_75t_L g1281 ( .A(n_972), .Y(n_1281) );
INVx2_ASAP7_75t_SL g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1038 ( .A(n_982), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1697 ( .A1(n_993), .A2(n_1657), .B1(n_1665), .B2(n_1698), .Y(n_1697) );
INVx1_ASAP7_75t_SL g1051 ( .A(n_995), .Y(n_1051) );
NAND4xp75_ASAP7_75t_L g995 ( .A(n_996), .B(n_1016), .C(n_1021), .D(n_1047), .Y(n_995) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI211xp5_ASAP7_75t_L g1037 ( .A1(n_1004), .A2(n_1038), .B(n_1039), .C(n_1040), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1332 ( .A1(n_1005), .A2(n_1333), .B1(n_1334), .B2(n_1335), .Y(n_1332) );
BUFx3_ASAP7_75t_L g1908 ( .A(n_1005), .Y(n_1908) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1007), .Y(n_1490) );
BUFx2_ASAP7_75t_L g1584 ( .A(n_1007), .Y(n_1584) );
BUFx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1328 ( .A(n_1013), .Y(n_1328) );
NOR2x1_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1020), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1037), .Y(n_1028) );
OAI211xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1031), .B(n_1033), .C(n_1034), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1621 ( .A1(n_1031), .A2(n_1068), .B1(n_1595), .B2(n_1598), .C(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1036), .Y(n_1225) );
INVx3_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1285), .Y(n_1055) );
XNOR2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1125), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
XNOR2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
AND4x1_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1063), .C(n_1092), .D(n_1118), .Y(n_1060) );
NOR3xp33_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1088), .C(n_1089), .Y(n_1063) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1069), .B1(n_1070), .B2(n_1073), .C(n_1074), .Y(n_1067) );
OAI221xp5_ASAP7_75t_L g1252 ( .A1(n_1068), .A2(n_1082), .B1(n_1253), .B2(n_1254), .C(n_1255), .Y(n_1252) );
OAI221xp5_ASAP7_75t_L g1244 ( .A1(n_1070), .A2(n_1080), .B1(n_1245), .B2(n_1246), .C(n_1247), .Y(n_1244) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1082), .B2(n_1084), .C(n_1085), .Y(n_1079) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1916 ( .A(n_1086), .Y(n_1916) );
BUFx3_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NOR3xp33_ASAP7_75t_SL g1242 ( .A(n_1088), .B(n_1243), .C(n_1256), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1099), .B1(n_1100), .B2(n_1103), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1900 ( .A1(n_1098), .A2(n_1207), .B1(n_1901), .B2(n_1902), .Y(n_1900) );
OAI22xp33_ASAP7_75t_L g1903 ( .A1(n_1098), .A2(n_1898), .B1(n_1904), .B2(n_1905), .Y(n_1903) );
OAI22xp5_ASAP7_75t_L g1274 ( .A1(n_1100), .A2(n_1275), .B1(n_1277), .B2(n_1278), .Y(n_1274) );
INVx2_ASAP7_75t_SL g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_1102), .A2(n_1275), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1120), .Y(n_1118) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
XOR2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1236), .Y(n_1126) );
XNOR2xp5_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1174), .Y(n_1127) );
NAND4xp25_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1154), .C(n_1156), .D(n_1169), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1136), .B(n_1141), .Y(n_1132) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g1162 ( .A1(n_1143), .A2(n_1144), .B1(n_1163), .B2(n_1165), .Y(n_1162) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1929 ( .A(n_1167), .Y(n_1929) );
XNOR2x1_ASAP7_75t_SL g1174 ( .A(n_1175), .B(n_1176), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1214), .Y(n_1176) );
NOR3xp33_ASAP7_75t_SL g1177 ( .A(n_1178), .B(n_1186), .C(n_1191), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1183), .Y(n_1178) );
HB1xp67_ASAP7_75t_L g1890 ( .A(n_1181), .Y(n_1890) );
INVx2_ASAP7_75t_SL g1187 ( .A(n_1188), .Y(n_1187) );
INVx2_ASAP7_75t_L g1892 ( .A(n_1188), .Y(n_1892) );
OAI33xp33_ASAP7_75t_L g1191 ( .A1(n_1192), .A2(n_1194), .A3(n_1198), .B1(n_1204), .B2(n_1209), .B3(n_1212), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g1573 ( .A1(n_1197), .A2(n_1574), .B1(n_1575), .B2(n_1576), .Y(n_1573) );
OAI22xp33_ASAP7_75t_L g1583 ( .A1(n_1197), .A2(n_1555), .B1(n_1557), .B2(n_1584), .Y(n_1583) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1200), .B1(n_1201), .B2(n_1202), .Y(n_1198) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1906 ( .A1(n_1207), .A2(n_1907), .B1(n_1908), .B2(n_1909), .Y(n_1906) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1208), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g1606 ( .A(n_1208), .Y(n_1606) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1212), .Y(n_1611) );
OAI33xp33_ASAP7_75t_L g1894 ( .A1(n_1212), .A2(n_1895), .A3(n_1896), .B1(n_1900), .B2(n_1903), .B3(n_1906), .Y(n_1894) );
CKINVDCx8_ASAP7_75t_R g1212 ( .A(n_1213), .Y(n_1212) );
NAND3xp33_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1226), .C(n_1234), .Y(n_1215) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1223), .Y(n_1620) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1223), .Y(n_1631) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1228), .Y(n_1460) );
INVx4_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1233), .Y(n_1404) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1233), .Y(n_1451) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
XNOR2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
AND4x1_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1242), .C(n_1259), .D(n_1282), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1251), .Y(n_1389) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
OAI31xp33_ASAP7_75t_L g1259 ( .A1(n_1260), .A2(n_1270), .A3(n_1279), .B(n_1280), .Y(n_1259) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1273), .Y(n_1433) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_SL g1280 ( .A(n_1281), .Y(n_1280) );
AOI22xp33_ASAP7_75t_SL g1910 ( .A1(n_1281), .A2(n_1911), .B1(n_1933), .B2(n_1934), .Y(n_1910) );
NOR2xp33_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1287), .B1(n_1492), .B2(n_1636), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
XNOR2x2_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1396), .Y(n_1287) );
XNOR2xp5_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1340), .Y(n_1288) );
XNOR2xp5_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1291), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1315), .Y(n_1291) );
NAND4xp25_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1302), .C(n_1308), .D(n_1311), .Y(n_1293) );
INVx1_ASAP7_75t_L g1926 ( .A(n_1297), .Y(n_1926) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx3_ASAP7_75t_L g1385 ( .A(n_1298), .Y(n_1385) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_1310), .A2(n_1312), .B1(n_1328), .B2(n_1339), .Y(n_1338) );
NOR3xp33_ASAP7_75t_SL g1315 ( .A(n_1316), .B(n_1323), .C(n_1326), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1320), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g1893 ( .A(n_1325), .Y(n_1893) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1329), .B1(n_1330), .B2(n_1331), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_1330), .A2(n_1436), .B1(n_1437), .B2(n_1438), .Y(n_1435) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_1337), .A2(n_1432), .B1(n_1433), .B2(n_1434), .Y(n_1431) );
OAI22xp33_ASAP7_75t_L g1477 ( .A1(n_1337), .A2(n_1478), .B1(n_1479), .B2(n_1480), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g1439 ( .A1(n_1339), .A2(n_1402), .B1(n_1419), .B2(n_1440), .Y(n_1439) );
XNOR2x1_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1395), .Y(n_1340) );
NAND2x1_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1368), .Y(n_1341) );
AND4x1_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1346), .C(n_1360), .D(n_1364), .Y(n_1342) );
BUFx3_ASAP7_75t_L g1604 ( .A(n_1349), .Y(n_1604) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1362), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_1367), .A2(n_1594), .B1(n_1595), .B2(n_1596), .Y(n_1593) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1367), .Y(n_1885) );
AOI22xp5_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1370), .B1(n_1393), .B2(n_1394), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_1369), .A2(n_1394), .B1(n_1400), .B2(n_1420), .Y(n_1399) );
AOI21xp5_ASAP7_75t_SL g1516 ( .A1(n_1369), .A2(n_1517), .B(n_1537), .Y(n_1516) );
NAND3xp33_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1381), .C(n_1390), .Y(n_1370) );
AOI21xp5_ASAP7_75t_SL g1371 ( .A1(n_1372), .A2(n_1373), .B(n_1374), .Y(n_1371) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1375), .Y(n_1520) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1385), .Y(n_1628) );
HB1xp67_ASAP7_75t_L g1630 ( .A(n_1387), .Y(n_1630) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1388), .Y(n_1531) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx2_ASAP7_75t_SL g1917 ( .A(n_1389), .Y(n_1917) );
AOI21xp5_ASAP7_75t_L g1612 ( .A1(n_1394), .A2(n_1613), .B(n_1614), .Y(n_1612) );
XNOR2xp5_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1443), .Y(n_1396) );
XOR2x2_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1442), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1421), .Y(n_1398) );
NAND3xp33_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1409), .C(n_1417), .Y(n_1400) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
NOR3xp33_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1429), .C(n_1430), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1426), .Y(n_1422) );
OAI22xp33_ASAP7_75t_L g1488 ( .A1(n_1433), .A2(n_1448), .B1(n_1453), .B2(n_1489), .Y(n_1488) );
OAI22xp5_ASAP7_75t_SL g1896 ( .A1(n_1433), .A2(n_1897), .B1(n_1898), .B2(n_1899), .Y(n_1896) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_1436), .A2(n_1482), .B1(n_1483), .B2(n_1486), .Y(n_1481) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_1440), .A2(n_1454), .B1(n_1466), .B2(n_1485), .Y(n_1487) );
XNOR2x1_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1491), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1468), .Y(n_1444) );
NAND5xp2_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1452), .C(n_1455), .D(n_1459), .E(n_1465), .Y(n_1446) );
OAI221xp5_ASAP7_75t_SL g1459 ( .A1(n_1460), .A2(n_1461), .B1(n_1462), .B2(n_1463), .C(n_1464), .Y(n_1459) );
NOR3xp33_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1474), .C(n_1476), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1472), .Y(n_1469) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx2_ASAP7_75t_SL g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1654 ( .A1(n_1491), .A2(n_1655), .B1(n_1661), .B2(n_1662), .Y(n_1654) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1492), .Y(n_1636) );
AO22x2_ASAP7_75t_L g1492 ( .A1(n_1493), .A2(n_1494), .B1(n_1586), .B2(n_1587), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
XNOR2xp5_ASAP7_75t_L g1494 ( .A(n_1495), .B(n_1541), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1516), .Y(n_1497) );
NOR2xp33_ASAP7_75t_L g1498 ( .A(n_1499), .B(n_1501), .Y(n_1498) );
NAND4xp25_ASAP7_75t_SL g1517 ( .A(n_1518), .B(n_1523), .C(n_1525), .D(n_1527), .Y(n_1517) );
OAI221xp5_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1530), .B1(n_1531), .B2(n_1532), .C(n_1533), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1536), .Y(n_1622) );
XNOR2x1_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1585), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1561), .Y(n_1542) );
NAND3xp33_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1551), .C(n_1556), .Y(n_1544) );
NOR3xp33_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1570), .C(n_1572), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1567), .Y(n_1562) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
INVx2_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
XOR2x2_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1635), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1612), .Y(n_1588) );
AND4x1_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1593), .C(n_1597), .D(n_1602), .Y(n_1589) );
INVxp67_ASAP7_75t_SL g1886 ( .A(n_1596), .Y(n_1886) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_1598), .A2(n_1599), .B1(n_1600), .B2(n_1601), .Y(n_1597) );
AOI22xp33_ASAP7_75t_L g1887 ( .A1(n_1599), .A2(n_1888), .B1(n_1889), .B2(n_1890), .Y(n_1887) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
OAI221xp5_ASAP7_75t_L g1637 ( .A1(n_1638), .A2(n_1879), .B1(n_1881), .B2(n_1936), .C(n_1940), .Y(n_1637) );
AND4x1_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1806), .C(n_1820), .D(n_1852), .Y(n_1638) );
AOI211xp5_ASAP7_75t_L g1639 ( .A1(n_1640), .A2(n_1667), .B(n_1768), .C(n_1782), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1783 ( .A(n_1640), .B(n_1784), .Y(n_1783) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1640), .B(n_1741), .Y(n_1829) );
AOI221xp5_ASAP7_75t_L g1847 ( .A1(n_1640), .A2(n_1717), .B1(n_1745), .B2(n_1848), .C(n_1849), .Y(n_1847) );
OAI333xp33_ASAP7_75t_L g1871 ( .A1(n_1640), .A2(n_1715), .A3(n_1773), .B1(n_1808), .B2(n_1872), .B3(n_1874), .C1(n_1875), .C2(n_1877), .C3(n_1878), .Y(n_1871) );
CKINVDCx5p33_ASAP7_75t_R g1640 ( .A(n_1641), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1641), .B(n_1775), .Y(n_1808) );
OAI32xp33_ASAP7_75t_L g1828 ( .A1(n_1641), .A2(n_1681), .A3(n_1741), .B1(n_1800), .B2(n_1829), .Y(n_1828) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1641), .Y(n_1862) );
NAND2xp5_ASAP7_75t_L g1877 ( .A(n_1641), .B(n_1700), .Y(n_1877) );
OR2x6_ASAP7_75t_SL g1641 ( .A(n_1642), .B(n_1654), .Y(n_1641) );
OAI22xp5_ASAP7_75t_L g1642 ( .A1(n_1643), .A2(n_1644), .B1(n_1651), .B2(n_1652), .Y(n_1642) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1645), .Y(n_1706) );
AND2x4_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1649), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1646), .B(n_1649), .Y(n_1674) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
AND2x4_ASAP7_75t_L g1653 ( .A(n_1647), .B(n_1649), .Y(n_1653) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1659 ( .A(n_1648), .B(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1650), .Y(n_1660) );
INVx2_ASAP7_75t_L g1691 ( .A(n_1652), .Y(n_1691) );
INVx2_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_SL g1676 ( .A(n_1653), .Y(n_1676) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1655), .Y(n_1880) );
BUFx3_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OAI22xp5_ASAP7_75t_L g1678 ( .A1(n_1656), .A2(n_1665), .B1(n_1679), .B2(n_1680), .Y(n_1678) );
OAI22xp33_ASAP7_75t_L g1719 ( .A1(n_1656), .A2(n_1665), .B1(n_1720), .B2(n_1721), .Y(n_1719) );
BUFx6f_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1659), .Y(n_1657) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1658), .B(n_1666), .Y(n_1665) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1658), .Y(n_1687) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1659), .Y(n_1686) );
HB1xp67_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1666), .Y(n_1689) );
NAND5xp2_ASAP7_75t_L g1667 ( .A(n_1668), .B(n_1736), .C(n_1749), .D(n_1757), .E(n_1761), .Y(n_1667) );
AOI211xp5_ASAP7_75t_SL g1668 ( .A1(n_1669), .A2(n_1699), .B(n_1711), .C(n_1732), .Y(n_1668) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1669), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1681), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1670), .B(n_1714), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1670), .B(n_1715), .Y(n_1731) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1670), .B(n_1683), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1760 ( .A(n_1670), .B(n_1683), .Y(n_1760) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1670), .B(n_1792), .Y(n_1791) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_1670), .B(n_1726), .Y(n_1803) );
OR2x2_ASAP7_75t_L g1805 ( .A(n_1670), .B(n_1726), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1827 ( .A(n_1670), .B(n_1725), .Y(n_1827) );
AND2x2_ASAP7_75t_L g1832 ( .A(n_1670), .B(n_1692), .Y(n_1832) );
NOR2xp33_ASAP7_75t_L g1843 ( .A(n_1670), .B(n_1743), .Y(n_1843) );
NOR2xp33_ASAP7_75t_L g1873 ( .A(n_1670), .B(n_1696), .Y(n_1873) );
CKINVDCx6p67_ASAP7_75t_R g1670 ( .A(n_1671), .Y(n_1670) );
OR2x2_ASAP7_75t_L g1763 ( .A(n_1671), .B(n_1715), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1671), .B(n_1750), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1671), .B(n_1715), .Y(n_1798) );
AND2x2_ASAP7_75t_L g1800 ( .A(n_1671), .B(n_1692), .Y(n_1800) );
NAND2xp5_ASAP7_75t_L g1812 ( .A(n_1671), .B(n_1813), .Y(n_1812) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1671), .B(n_1714), .Y(n_1816) );
AND2x2_ASAP7_75t_L g1846 ( .A(n_1671), .B(n_1725), .Y(n_1846) );
OR2x2_ASAP7_75t_L g1855 ( .A(n_1671), .B(n_1751), .Y(n_1855) );
OR2x6_ASAP7_75t_SL g1671 ( .A(n_1672), .B(n_1678), .Y(n_1671) );
OAI22xp5_ASAP7_75t_L g1672 ( .A1(n_1673), .A2(n_1675), .B1(n_1676), .B2(n_1677), .Y(n_1672) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
OAI22xp5_ASAP7_75t_L g1704 ( .A1(n_1676), .A2(n_1705), .B1(n_1706), .B2(n_1707), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1682), .B(n_1692), .Y(n_1681) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1682), .B(n_1713), .Y(n_1712) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1682), .Y(n_1724) );
NOR2xp33_ASAP7_75t_L g1776 ( .A(n_1682), .B(n_1777), .Y(n_1776) );
NOR2xp33_ASAP7_75t_L g1813 ( .A(n_1682), .B(n_1751), .Y(n_1813) );
INVx4_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1683), .B(n_1731), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1743 ( .A(n_1683), .B(n_1692), .Y(n_1743) );
INVx2_ASAP7_75t_L g1755 ( .A(n_1683), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1683), .B(n_1701), .Y(n_1792) );
OR2x2_ASAP7_75t_L g1839 ( .A(n_1683), .B(n_1766), .Y(n_1839) );
NAND2xp5_ASAP7_75t_L g1845 ( .A(n_1683), .B(n_1846), .Y(n_1845) );
OR2x2_ASAP7_75t_L g1850 ( .A(n_1683), .B(n_1751), .Y(n_1850) );
OR2x2_ASAP7_75t_L g1854 ( .A(n_1683), .B(n_1855), .Y(n_1854) );
NAND2xp5_ASAP7_75t_L g1874 ( .A(n_1683), .B(n_1767), .Y(n_1874) );
AND2x2_ASAP7_75t_L g1876 ( .A(n_1683), .B(n_1745), .Y(n_1876) );
AND2x6_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1690), .Y(n_1683) );
AND2x4_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1687), .Y(n_1685) );
OAI21xp33_ASAP7_75t_SL g1948 ( .A1(n_1686), .A2(n_1944), .B(n_1949), .Y(n_1948) );
AND2x4_ASAP7_75t_L g1688 ( .A(n_1687), .B(n_1689), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1696), .Y(n_1692) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1693), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1693), .B(n_1726), .Y(n_1725) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1693), .B(n_1696), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1695), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1696), .B(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1696), .Y(n_1726) );
NAND2xp5_ASAP7_75t_L g1780 ( .A(n_1699), .B(n_1781), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1859 ( .A(n_1699), .B(n_1848), .Y(n_1859) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1700), .B(n_1708), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1700), .B(n_1717), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1700), .B(n_1729), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1700), .B(n_1741), .Y(n_1740) );
OR2x2_ASAP7_75t_L g1773 ( .A(n_1700), .B(n_1708), .Y(n_1773) );
INVx3_ASAP7_75t_L g1775 ( .A(n_1700), .Y(n_1775) );
AOI21xp5_ASAP7_75t_L g1867 ( .A1(n_1700), .A2(n_1868), .B(n_1871), .Y(n_1867) );
INVx3_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1734 ( .A(n_1701), .B(n_1735), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1866 ( .A(n_1701), .B(n_1708), .Y(n_1866) );
OR2x2_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1704), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1708), .B(n_1718), .Y(n_1717) );
OR2x2_ASAP7_75t_L g1735 ( .A(n_1708), .B(n_1718), .Y(n_1735) );
INVx2_ASAP7_75t_L g1741 ( .A(n_1708), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1708), .B(n_1729), .Y(n_1745) );
OR2x2_ASAP7_75t_L g1756 ( .A(n_1708), .B(n_1729), .Y(n_1756) );
AOI22xp5_ASAP7_75t_L g1809 ( .A1(n_1708), .A2(n_1777), .B1(n_1810), .B2(n_1814), .Y(n_1809) );
OAI221xp5_ASAP7_75t_L g1836 ( .A1(n_1708), .A2(n_1835), .B1(n_1837), .B2(n_1845), .C(n_1847), .Y(n_1836) );
AND2x4_ASAP7_75t_L g1708 ( .A(n_1709), .B(n_1710), .Y(n_1708) );
OAI21xp5_ASAP7_75t_SL g1711 ( .A1(n_1712), .A2(n_1716), .B(n_1722), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1713), .B(n_1775), .Y(n_1774) );
A2O1A1Ixp33_ASAP7_75t_SL g1806 ( .A1(n_1713), .A2(n_1807), .B(n_1809), .C(n_1817), .Y(n_1806) );
AOI211xp5_ASAP7_75t_L g1837 ( .A1(n_1713), .A2(n_1838), .B(n_1840), .C(n_1844), .Y(n_1837) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1714), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1714), .B(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
AOI322xp5_ASAP7_75t_L g1787 ( .A1(n_1717), .A2(n_1740), .A3(n_1788), .B1(n_1790), .B2(n_1793), .C1(n_1796), .C2(n_1801), .Y(n_1787) );
INVx2_ASAP7_75t_SL g1729 ( .A(n_1718), .Y(n_1729) );
HB1xp67_ASAP7_75t_L g1739 ( .A(n_1718), .Y(n_1739) );
AOI22xp5_ASAP7_75t_L g1722 ( .A1(n_1723), .A2(n_1727), .B1(n_1728), .B2(n_1730), .Y(n_1722) );
INVxp67_ASAP7_75t_L g1878 ( .A(n_1723), .Y(n_1878) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1725), .Y(n_1723) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1725), .Y(n_1789) );
NOR2xp33_ASAP7_75t_L g1872 ( .A(n_1725), .B(n_1873), .Y(n_1872) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1728), .Y(n_1856) );
INVx2_ASAP7_75t_SL g1767 ( .A(n_1729), .Y(n_1767) );
NOR2xp33_ASAP7_75t_L g1732 ( .A(n_1733), .B(n_1734), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1733), .B(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1734), .Y(n_1801) );
INVx1_ASAP7_75t_L g1819 ( .A(n_1735), .Y(n_1819) );
OAI21xp33_ASAP7_75t_SL g1830 ( .A1(n_1735), .A2(n_1831), .B(n_1833), .Y(n_1830) );
AOI21xp5_ASAP7_75t_L g1736 ( .A1(n_1737), .A2(n_1742), .B(n_1744), .Y(n_1736) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1738 ( .A(n_1739), .B(n_1740), .Y(n_1738) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1739), .Y(n_1770) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_1739), .B(n_1786), .Y(n_1785) );
NAND2xp5_ASAP7_75t_L g1814 ( .A(n_1739), .B(n_1815), .Y(n_1814) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1739), .Y(n_1835) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1739), .Y(n_1842) );
AOI211xp5_ASAP7_75t_SL g1857 ( .A1(n_1740), .A2(n_1858), .B(n_1859), .C(n_1860), .Y(n_1857) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
A2O1A1Ixp33_ASAP7_75t_L g1853 ( .A1(n_1743), .A2(n_1854), .B(n_1856), .C(n_1857), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1745), .B(n_1746), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1745), .B(n_1758), .Y(n_1757) );
AOI21xp5_ASAP7_75t_L g1817 ( .A1(n_1745), .A2(n_1818), .B(n_1819), .Y(n_1817) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1745), .Y(n_1823) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
NOR2xp33_ASAP7_75t_L g1779 ( .A(n_1747), .B(n_1780), .Y(n_1779) );
NAND2xp5_ASAP7_75t_L g1772 ( .A(n_1748), .B(n_1750), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1752), .Y(n_1749) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1750), .B(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
OAI211xp5_ASAP7_75t_L g1802 ( .A1(n_1752), .A2(n_1775), .B(n_1803), .C(n_1804), .Y(n_1802) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
OR2x2_ASAP7_75t_L g1753 ( .A(n_1754), .B(n_1756), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g1797 ( .A(n_1754), .B(n_1798), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1754), .B(n_1816), .Y(n_1815) );
NOR2x1_ASAP7_75t_L g1848 ( .A(n_1754), .B(n_1805), .Y(n_1848) );
INVx2_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1765 ( .A(n_1755), .B(n_1766), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1858 ( .A(n_1755), .B(n_1762), .Y(n_1858) );
INVx2_ASAP7_75t_L g1777 ( .A(n_1756), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1834 ( .A(n_1758), .B(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
NOR2xp33_ASAP7_75t_L g1870 ( .A(n_1759), .B(n_1835), .Y(n_1870) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1760), .Y(n_1795) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1764), .Y(n_1761) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1767), .Y(n_1781) );
OAI21xp33_ASAP7_75t_L g1868 ( .A1(n_1767), .A2(n_1794), .B(n_1869), .Y(n_1868) );
OAI221xp5_ASAP7_75t_L g1768 ( .A1(n_1769), .A2(n_1773), .B1(n_1774), .B2(n_1776), .C(n_1778), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1770), .B(n_1771), .Y(n_1769) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_SL g1784 ( .A(n_1775), .Y(n_1784) );
NOR3xp33_ASAP7_75t_L g1860 ( .A(n_1775), .B(n_1789), .C(n_1839), .Y(n_1860) );
INVxp67_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
NOR2xp33_ASAP7_75t_L g1811 ( .A(n_1781), .B(n_1812), .Y(n_1811) );
OAI211xp5_ASAP7_75t_SL g1782 ( .A1(n_1783), .A2(n_1785), .B(n_1787), .C(n_1802), .Y(n_1782) );
OAI311xp33_ASAP7_75t_L g1820 ( .A1(n_1783), .A2(n_1821), .A3(n_1822), .B1(n_1830), .C1(n_1836), .Y(n_1820) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1786), .Y(n_1825) );
OR2x2_ASAP7_75t_L g1794 ( .A(n_1789), .B(n_1795), .Y(n_1794) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
NAND2xp33_ASAP7_75t_L g1796 ( .A(n_1797), .B(n_1799), .Y(n_1796) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1812), .Y(n_1844) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1814), .Y(n_1821) );
INVxp67_ASAP7_75t_L g1864 ( .A(n_1815), .Y(n_1864) );
OAI21xp33_ASAP7_75t_L g1822 ( .A1(n_1823), .A2(n_1824), .B(n_1828), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1824 ( .A(n_1825), .B(n_1826), .Y(n_1824) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
A2O1A1Ixp33_ASAP7_75t_L g1863 ( .A1(n_1833), .A2(n_1864), .B(n_1865), .C(n_1867), .Y(n_1863) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
NAND2xp5_ASAP7_75t_L g1841 ( .A(n_1842), .B(n_1843), .Y(n_1841) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1846), .Y(n_1851) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1850), .B(n_1851), .Y(n_1849) );
AOI21xp5_ASAP7_75t_L g1852 ( .A1(n_1853), .A2(n_1861), .B(n_1863), .Y(n_1852) );
CKINVDCx14_ASAP7_75t_R g1861 ( .A(n_1862), .Y(n_1861) );
INVx1_ASAP7_75t_L g1865 ( .A(n_1866), .Y(n_1865) );
INVxp33_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1876), .Y(n_1875) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
AND2x2_ASAP7_75t_L g1882 ( .A(n_1883), .B(n_1910), .Y(n_1882) );
NOR3xp33_ASAP7_75t_SL g1883 ( .A(n_1884), .B(n_1891), .C(n_1894), .Y(n_1883) );
AOI211xp5_ASAP7_75t_L g1912 ( .A1(n_1905), .A2(n_1913), .B(n_1914), .C(n_1915), .Y(n_1912) );
AOI221xp5_ASAP7_75t_L g1921 ( .A1(n_1909), .A2(n_1922), .B1(n_1924), .B2(n_1928), .C(n_1930), .Y(n_1921) );
NAND3xp33_ASAP7_75t_L g1911 ( .A(n_1912), .B(n_1921), .C(n_1932), .Y(n_1911) );
INVx1_ASAP7_75t_L g1922 ( .A(n_1923), .Y(n_1922) );
INVx1_ASAP7_75t_L g1925 ( .A(n_1926), .Y(n_1925) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
INVx1_ASAP7_75t_L g1934 ( .A(n_1935), .Y(n_1934) );
INVx2_ASAP7_75t_L g1936 ( .A(n_1937), .Y(n_1936) );
INVx1_ASAP7_75t_L g1937 ( .A(n_1938), .Y(n_1937) );
INVx1_ASAP7_75t_L g1938 ( .A(n_1939), .Y(n_1938) );
INVx2_ASAP7_75t_L g1941 ( .A(n_1942), .Y(n_1941) );
CKINVDCx5p33_ASAP7_75t_R g1942 ( .A(n_1943), .Y(n_1942) );
INVxp33_ASAP7_75t_SL g1945 ( .A(n_1946), .Y(n_1945) );
HB1xp67_ASAP7_75t_L g1947 ( .A(n_1948), .Y(n_1947) );
endmodule