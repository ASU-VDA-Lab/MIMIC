module fake_jpeg_18838_n_12 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_12);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_12;

wire n_11;
wire n_10;
wire n_8;
wire n_9;
wire n_7;

A2O1A1Ixp33_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_6),
.B(n_4),
.C(n_2),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_7),
.B(n_8),
.Y(n_9)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_3),
.C(n_5),
.Y(n_12)
);


endmodule