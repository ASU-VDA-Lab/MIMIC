module real_aes_16463_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AND2x4_ASAP7_75t_L g837 ( .A(n_0), .B(n_838), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_1), .A2(n_4), .B1(n_247), .B2(n_248), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_2), .A2(n_43), .B1(n_148), .B2(n_196), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_3), .A2(n_25), .B1(n_196), .B2(n_230), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_5), .A2(n_16), .B1(n_498), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_6), .A2(n_60), .B1(n_133), .B2(n_134), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_7), .A2(n_17), .B1(n_148), .B2(n_149), .Y(n_147) );
INVx1_ASAP7_75t_L g838 ( .A(n_8), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_9), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_10), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_11), .A2(n_18), .B1(n_499), .B2(n_543), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_12), .A2(n_64), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_12), .Y(n_777) );
OR2x2_ASAP7_75t_L g791 ( .A(n_13), .B(n_39), .Y(n_791) );
BUFx2_ASAP7_75t_L g832 ( .A(n_13), .Y(n_832) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_14), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_15), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_19), .A2(n_100), .B1(n_248), .B2(n_498), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_20), .A2(n_38), .B1(n_126), .B2(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_21), .B(n_124), .Y(n_559) );
OAI22x1_ASAP7_75t_SL g774 ( .A1(n_22), .A2(n_775), .B1(n_776), .B2(n_779), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_22), .Y(n_779) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_23), .A2(n_58), .B(n_139), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_24), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_26), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_27), .B(n_121), .Y(n_188) );
INVx4_ASAP7_75t_R g172 ( .A(n_28), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_29), .A2(n_47), .B1(n_152), .B2(n_245), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_30), .A2(n_54), .B1(n_152), .B2(n_498), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_31), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_32), .B(n_523), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_33), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_34), .B(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g252 ( .A(n_35), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_SL g227 ( .A1(n_36), .A2(n_120), .B(n_148), .C(n_228), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_37), .A2(n_55), .B1(n_148), .B2(n_152), .Y(n_236) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_39), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_40), .A2(n_88), .B1(n_148), .B2(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_SL g795 ( .A1(n_41), .A2(n_53), .B1(n_796), .B2(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_41), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_42), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_44), .A2(n_46), .B1(n_148), .B2(n_149), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_45), .A2(n_59), .B1(n_498), .B2(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g192 ( .A(n_48), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_49), .B(n_148), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_50), .Y(n_206) );
INVx2_ASAP7_75t_L g786 ( .A(n_51), .Y(n_786) );
BUFx3_ASAP7_75t_L g789 ( .A(n_52), .Y(n_789) );
INVx1_ASAP7_75t_L g807 ( .A(n_52), .Y(n_807) );
INVx1_ASAP7_75t_L g796 ( .A(n_53), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_56), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_57), .A2(n_89), .B1(n_148), .B2(n_152), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_61), .A2(n_77), .B1(n_245), .B2(n_515), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_62), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_63), .A2(n_80), .B1(n_148), .B2(n_149), .Y(n_500) );
INVx1_ASAP7_75t_L g778 ( .A(n_64), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_65), .A2(n_99), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g139 ( .A(n_66), .Y(n_139) );
AND2x4_ASAP7_75t_L g142 ( .A(n_67), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_68), .A2(n_808), .B(n_820), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_69), .A2(n_91), .B1(n_152), .B2(n_245), .Y(n_244) );
AO22x1_ASAP7_75t_L g122 ( .A1(n_70), .A2(n_78), .B1(n_123), .B2(n_126), .Y(n_122) );
INVx1_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
AND2x2_ASAP7_75t_L g231 ( .A(n_72), .B(n_184), .Y(n_231) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_72), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_73), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_799) );
CKINVDCx14_ASAP7_75t_R g802 ( .A(n_73), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_74), .A2(n_105), .B1(n_827), .B2(n_840), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_75), .B(n_133), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_76), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_79), .B(n_196), .Y(n_207) );
INVx2_ASAP7_75t_L g121 ( .A(n_81), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_82), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_83), .B(n_184), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_84), .A2(n_98), .B1(n_133), .B2(n_152), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_85), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_86), .B(n_137), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_87), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_90), .B(n_184), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_92), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_93), .B(n_184), .Y(n_203) );
INVx1_ASAP7_75t_L g470 ( .A(n_94), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_94), .B(n_806), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g562 ( .A(n_95), .B(n_124), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_96), .A2(n_133), .B(n_154), .C(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g177 ( .A(n_97), .B(n_178), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_101), .A2(n_107), .B1(n_108), .B2(n_781), .Y(n_106) );
INVx1_ASAP7_75t_SL g781 ( .A(n_101), .Y(n_781) );
NAND2xp33_ASAP7_75t_L g211 ( .A(n_102), .B(n_173), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_103), .Y(n_809) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_782), .B(n_792), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_110), .B1(n_774), .B2(n_780), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_467), .B1(n_471), .B2(n_773), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_377), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_306), .C(n_348), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_280), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_179), .B1(n_255), .B2(n_266), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_160), .Y(n_116) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_117), .A2(n_300), .B(n_302), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_117), .A2(n_373), .B(n_374), .Y(n_372) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_144), .Y(n_117) );
INVx2_ASAP7_75t_L g292 ( .A(n_118), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_118), .B(n_145), .Y(n_322) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_122), .B(n_128), .C(n_140), .Y(n_119) );
INVx6_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_120), .A2(n_211), .B(n_212), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_120), .B(n_122), .Y(n_264) );
O2A1O1Ixp5_ASAP7_75t_L g557 ( .A1(n_120), .A2(n_149), .B(n_558), .C(n_559), .Y(n_557) );
BUFx8_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
INVx1_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
INVx1_ASAP7_75t_L g191 ( .A(n_121), .Y(n_191) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g498 ( .A(n_124), .Y(n_498) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g127 ( .A(n_125), .Y(n_127) );
INVx1_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_125), .Y(n_135) );
INVx3_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_125), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_125), .Y(n_196) );
INVx1_ASAP7_75t_L g224 ( .A(n_125), .Y(n_224) );
INVx2_ASAP7_75t_L g230 ( .A(n_125), .Y(n_230) );
OAI21xp33_ASAP7_75t_SL g187 ( .A1(n_126), .A2(n_188), .B(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g263 ( .A(n_128), .Y(n_263) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B(n_136), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_129), .A2(n_194), .B(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_129), .A2(n_150), .B1(n_235), .B2(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g481 ( .A(n_130), .Y(n_481) );
BUFx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
INVx1_ASAP7_75t_L g543 ( .A(n_134), .Y(n_543) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_135), .B(n_169), .Y(n_168) );
OAI21xp33_ASAP7_75t_L g140 ( .A1(n_136), .A2(n_137), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g155 ( .A(n_137), .Y(n_155) );
INVx2_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
INVx2_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
INVx1_ASAP7_75t_L g265 ( .A(n_140), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_141), .A2(n_220), .B(n_227), .Y(n_219) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx10_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
BUFx10_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
INVx1_ASAP7_75t_L g250 ( .A(n_142), .Y(n_250) );
AND2x2_ASAP7_75t_L g362 ( .A(n_144), .B(n_201), .Y(n_362) );
INVx1_ASAP7_75t_L g395 ( .A(n_144), .Y(n_395) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g257 ( .A(n_145), .B(n_202), .Y(n_257) );
AND2x2_ASAP7_75t_L g288 ( .A(n_145), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g297 ( .A(n_145), .Y(n_297) );
OR2x2_ASAP7_75t_L g316 ( .A(n_145), .B(n_162), .Y(n_316) );
AND2x2_ASAP7_75t_L g331 ( .A(n_145), .B(n_162), .Y(n_331) );
AO31x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_155), .A3(n_156), .B(n_157), .Y(n_145) );
OAI22x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B1(n_151), .B2(n_153), .Y(n_146) );
INVx4_ASAP7_75t_L g149 ( .A(n_148), .Y(n_149) );
INVx1_ASAP7_75t_L g499 ( .A(n_148), .Y(n_499) );
INVx1_ASAP7_75t_L g515 ( .A(n_148), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_149), .A2(n_206), .B(n_207), .C(n_208), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_150), .A2(n_153), .B1(n_244), .B2(n_246), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_150), .A2(n_480), .B1(n_481), .B2(n_482), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_150), .A2(n_153), .B1(n_489), .B2(n_491), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_150), .A2(n_497), .B1(n_500), .B2(n_501), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_150), .A2(n_481), .B1(n_513), .B2(n_514), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_150), .A2(n_481), .B1(n_522), .B2(n_524), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_150), .A2(n_481), .B1(n_532), .B2(n_533), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_150), .A2(n_501), .B1(n_542), .B2(n_544), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_150), .A2(n_561), .B(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_152), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g247 ( .A(n_152), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_153), .B(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g501 ( .A(n_154), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_155), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_155), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
AO31x2_ASAP7_75t_L g478 ( .A1(n_156), .A2(n_237), .A3(n_479), .B(n_483), .Y(n_478) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_156), .A2(n_487), .A3(n_521), .B(n_526), .Y(n_520) );
AO31x2_ASAP7_75t_L g540 ( .A1(n_156), .A2(n_218), .A3(n_541), .B(n_545), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx2_ASAP7_75t_L g178 ( .A(n_159), .Y(n_178) );
BUFx2_ASAP7_75t_L g218 ( .A(n_159), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_159), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_159), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_161), .B(n_330), .Y(n_373) );
OR2x2_ASAP7_75t_L g461 ( .A(n_161), .B(n_322), .Y(n_461) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g289 ( .A(n_162), .Y(n_289) );
AND2x2_ASAP7_75t_L g298 ( .A(n_162), .B(n_261), .Y(n_298) );
AND2x2_ASAP7_75t_L g301 ( .A(n_162), .B(n_202), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_162), .B(n_201), .Y(n_320) );
AND2x4_ASAP7_75t_L g339 ( .A(n_162), .B(n_262), .Y(n_339) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_177), .Y(n_162) );
AO31x2_ASAP7_75t_L g511 ( .A1(n_163), .A2(n_502), .A3(n_512), .B(n_516), .Y(n_511) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_163), .A2(n_249), .A3(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_165), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_SL g545 ( .A(n_165), .B(n_546), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_176), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_171) );
INVx2_ASAP7_75t_L g245 ( .A(n_173), .Y(n_245) );
INVx1_ASAP7_75t_L g523 ( .A(n_173), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_174), .Y(n_525) );
INVx1_ASAP7_75t_L g502 ( .A(n_176), .Y(n_502) );
OAI21xp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_199), .B(n_240), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_180), .B(n_334), .Y(n_437) );
CKINVDCx14_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_182), .B(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g270 ( .A(n_182), .Y(n_270) );
OR2x2_ASAP7_75t_L g278 ( .A(n_182), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_182), .B(n_271), .Y(n_303) );
AND2x2_ASAP7_75t_L g328 ( .A(n_182), .B(n_242), .Y(n_328) );
AND2x2_ASAP7_75t_L g346 ( .A(n_182), .B(n_276), .Y(n_346) );
INVx1_ASAP7_75t_L g385 ( .A(n_182), .Y(n_385) );
AND2x2_ASAP7_75t_L g387 ( .A(n_182), .B(n_388), .Y(n_387) );
NAND2x1p5_ASAP7_75t_SL g406 ( .A(n_182), .B(n_327), .Y(n_406) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_186), .Y(n_182) );
NOR2x1_ASAP7_75t_L g213 ( .A(n_184), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g197 ( .A(n_185), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_185), .B(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g487 ( .A(n_185), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_185), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_185), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g555 ( .A(n_185), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_193), .B(n_197), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
BUFx4f_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_196), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g214 ( .A(n_198), .Y(n_214) );
AO31x2_ASAP7_75t_L g233 ( .A1(n_198), .A2(n_234), .A3(n_237), .B(n_238), .Y(n_233) );
OAI32xp33_ASAP7_75t_L g290 ( .A1(n_199), .A2(n_282), .A3(n_291), .B1(n_293), .B2(n_295), .Y(n_290) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_215), .Y(n_199) );
INVx1_ASAP7_75t_L g330 ( .A(n_200), .Y(n_330) );
AND2x2_ASAP7_75t_L g338 ( .A(n_200), .B(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g337 ( .A(n_201), .B(n_261), .Y(n_337) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx3_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
AND2x2_ASAP7_75t_L g296 ( .A(n_202), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g402 ( .A(n_202), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_210), .B(n_213), .Y(n_204) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g272 ( .A(n_215), .Y(n_272) );
OR2x2_ASAP7_75t_L g282 ( .A(n_215), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g404 ( .A(n_215), .Y(n_404) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_232), .Y(n_215) );
AND2x2_ASAP7_75t_L g305 ( .A(n_216), .B(n_233), .Y(n_305) );
INVx2_ASAP7_75t_L g327 ( .A(n_216), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_216), .B(n_242), .Y(n_347) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g254 ( .A(n_217), .Y(n_254) );
AOI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_231), .Y(n_217) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_218), .A2(n_243), .A3(n_249), .B(n_251), .Y(n_242) );
AO31x2_ASAP7_75t_L g495 ( .A1(n_218), .A2(n_496), .A3(n_502), .B(n_503), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_223), .B(n_226), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g248 ( .A(n_224), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_SL g490 ( .A(n_230), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_232), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g336 ( .A(n_232), .Y(n_336) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
BUFx2_ASAP7_75t_L g276 ( .A(n_233), .Y(n_276) );
OR2x2_ASAP7_75t_L g342 ( .A(n_233), .B(n_242), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_233), .B(n_242), .Y(n_375) );
INVx2_ASAP7_75t_L g323 ( .A(n_240), .Y(n_323) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_253), .Y(n_240) );
OR2x2_ASAP7_75t_L g310 ( .A(n_241), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g388 ( .A(n_241), .Y(n_388) );
INVx1_ASAP7_75t_L g271 ( .A(n_242), .Y(n_271) );
INVx1_ASAP7_75t_L g279 ( .A(n_242), .Y(n_279) );
INVx1_ASAP7_75t_L g294 ( .A(n_242), .Y(n_294) );
AO31x2_ASAP7_75t_L g486 ( .A1(n_249), .A2(n_487), .A3(n_488), .B(n_492), .Y(n_486) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_SL g563 ( .A(n_250), .Y(n_563) );
OR2x2_ASAP7_75t_L g398 ( .A(n_253), .B(n_375), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_254), .B(n_270), .Y(n_311) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
OR2x2_ASAP7_75t_L g412 ( .A(n_254), .B(n_336), .Y(n_412) );
INVxp67_ASAP7_75t_L g436 ( .A(n_254), .Y(n_436) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_257), .B(n_298), .Y(n_365) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g314 ( .A(n_259), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g427 ( .A(n_260), .Y(n_427) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g456 ( .A(n_261), .B(n_289), .Y(n_456) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g382 ( .A(n_262), .B(n_289), .Y(n_382) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_273), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_269), .B(n_305), .Y(n_419) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g283 ( .A(n_270), .Y(n_283) );
AND2x2_ASAP7_75t_L g333 ( .A(n_270), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_270), .B(n_327), .Y(n_376) );
OR2x2_ASAP7_75t_L g448 ( .A(n_270), .B(n_335), .Y(n_448) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g368 ( .A(n_274), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx2_ASAP7_75t_L g359 ( .A(n_275), .Y(n_359) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g349 ( .A(n_278), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_278), .Y(n_360) );
OR2x2_ASAP7_75t_L g411 ( .A(n_278), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g466 ( .A(n_278), .Y(n_466) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B(n_290), .C(n_299), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g355 ( .A(n_283), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_283), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g428 ( .A(n_283), .B(n_305), .Y(n_428) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_286), .B(n_331), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_286), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g438 ( .A(n_286), .B(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g381 ( .A(n_287), .Y(n_381) );
AND2x2_ASAP7_75t_L g409 ( .A(n_288), .B(n_337), .Y(n_409) );
INVx2_ASAP7_75t_L g432 ( .A(n_288), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_288), .B(n_330), .Y(n_464) );
AND2x4_ASAP7_75t_SL g418 ( .A(n_291), .B(n_296), .Y(n_418) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g371 ( .A(n_292), .B(n_297), .Y(n_371) );
OR2x2_ASAP7_75t_L g423 ( .A(n_292), .B(n_316), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_293), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_293), .B(n_305), .Y(n_459) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g407 ( .A(n_294), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g390 ( .A(n_296), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_296), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g440 ( .A(n_297), .Y(n_440) );
BUFx2_ASAP7_75t_L g308 ( .A(n_298), .Y(n_308) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g426 ( .A(n_301), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_305), .Y(n_367) );
NAND3xp33_ASAP7_75t_SL g306 ( .A(n_307), .B(n_317), .C(n_332), .Y(n_306) );
AOI22xp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_309), .B1(n_312), .B2(n_314), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_314), .A2(n_340), .B1(n_421), .B2(n_424), .C1(n_426), .C2(n_428), .Y(n_420) );
AND2x2_ASAP7_75t_L g452 ( .A(n_315), .B(n_401), .Y(n_452) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g400 ( .A(n_316), .B(n_401), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_323), .B1(n_324), .B2(n_329), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx2_ASAP7_75t_SL g396 ( .A(n_320), .Y(n_396) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
AND2x2_ASAP7_75t_L g383 ( .A(n_325), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g341 ( .A(n_326), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g335 ( .A(n_327), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g450 ( .A(n_328), .Y(n_450) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_331), .B(n_427), .Y(n_446) );
INVx1_ASAP7_75t_L g463 ( .A(n_331), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_337), .B1(n_338), .B2(n_340), .C1(n_343), .C2(n_344), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_339), .Y(n_343) );
AND2x2_ASAP7_75t_L g361 ( .A(n_339), .B(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g392 ( .A(n_339), .Y(n_392) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g356 ( .A(n_342), .Y(n_356) );
OR2x2_ASAP7_75t_L g425 ( .A(n_342), .B(n_406), .Y(n_425) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_354), .C(n_363), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_361), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_355), .A2(n_393), .B1(n_442), .B2(n_445), .C(n_447), .Y(n_441) );
AND2x4_ASAP7_75t_L g384 ( .A(n_356), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
AOI211x1_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_368), .C(n_372), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_374), .B(n_422), .C(n_423), .Y(n_421) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g457 ( .A(n_375), .Y(n_457) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_429), .Y(n_377) );
NAND4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_386), .C(n_408), .D(n_420), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g439 ( .A(n_382), .B(n_440), .Y(n_439) );
AOI221x1_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_409), .B1(n_410), .B2(n_413), .C(n_416), .Y(n_408) );
AND2x2_ASAP7_75t_L g434 ( .A(n_384), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_393), .B2(n_397), .C(n_399), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_391), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_396), .A2(n_400), .B1(n_403), .B2(n_405), .Y(n_399) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_400), .A2(n_417), .B(n_419), .Y(n_416) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_425), .A2(n_463), .B1(n_464), .B2(n_465), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_441), .C(n_453), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B1(n_437), .B2(n_438), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g449 ( .A(n_436), .B(n_450), .Y(n_449) );
NAND2x1_ASAP7_75t_L g465 ( .A(n_436), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B1(n_458), .B2(n_460), .C(n_462), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx4_ASAP7_75t_L g773 ( .A(n_467), .Y(n_773) );
BUFx12f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g825 ( .A(n_469), .B(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g839 ( .A(n_470), .Y(n_839) );
XNOR2xp5_ASAP7_75t_L g794 ( .A(n_471), .B(n_795), .Y(n_794) );
NOR2x1p5_ASAP7_75t_L g471 ( .A(n_472), .B(n_683), .Y(n_471) );
NAND4xp75_ASAP7_75t_L g472 ( .A(n_473), .B(n_628), .C(n_648), .D(n_664), .Y(n_472) );
NOR2x1p5_ASAP7_75t_SL g473 ( .A(n_474), .B(n_598), .Y(n_473) );
NAND4xp75_ASAP7_75t_L g474 ( .A(n_475), .B(n_536), .C(n_575), .D(n_584), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_505), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
AND2x4_ASAP7_75t_L g708 ( .A(n_477), .B(n_635), .Y(n_708) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_478), .Y(n_551) );
INVx2_ASAP7_75t_L g569 ( .A(n_478), .Y(n_569) );
AND2x2_ASAP7_75t_L g592 ( .A(n_478), .B(n_554), .Y(n_592) );
OR2x2_ASAP7_75t_L g647 ( .A(n_478), .B(n_486), .Y(n_647) );
AND2x2_ASAP7_75t_L g565 ( .A(n_485), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g715 ( .A(n_485), .B(n_592), .Y(n_715) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
OR2x2_ASAP7_75t_L g552 ( .A(n_486), .B(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
AND2x2_ASAP7_75t_L g589 ( .A(n_486), .B(n_495), .Y(n_589) );
INVx1_ASAP7_75t_L g607 ( .A(n_486), .Y(n_607) );
INVx2_ASAP7_75t_L g636 ( .A(n_486), .Y(n_636) );
INVx3_ASAP7_75t_L g612 ( .A(n_494), .Y(n_612) );
INVx2_ASAP7_75t_L g617 ( .A(n_494), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_494), .B(n_568), .Y(n_622) );
AND2x2_ASAP7_75t_L g645 ( .A(n_494), .B(n_624), .Y(n_645) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_494), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_494), .B(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g634 ( .A(n_495), .Y(n_634) );
AND2x2_ASAP7_75t_L g682 ( .A(n_495), .B(n_636), .Y(n_682) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_507), .B(n_626), .Y(n_673) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_508), .B(n_626), .Y(n_670) );
INVx1_ASAP7_75t_L g771 ( .A(n_508), .Y(n_771) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g721 ( .A(n_509), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g574 ( .A(n_510), .Y(n_574) );
OR2x2_ASAP7_75t_L g655 ( .A(n_510), .B(n_529), .Y(n_655) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g597 ( .A(n_511), .Y(n_597) );
AND2x4_ASAP7_75t_L g603 ( .A(n_511), .B(n_604), .Y(n_603) );
AOI32xp33_ASAP7_75t_L g741 ( .A1(n_518), .A2(n_644), .A3(n_742), .B1(n_744), .B2(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g690 ( .A(n_519), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .Y(n_519) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_520), .Y(n_538) );
OR2x2_ASAP7_75t_L g572 ( .A(n_520), .B(n_530), .Y(n_572) );
INVx1_ASAP7_75t_L g587 ( .A(n_520), .Y(n_587) );
AND2x2_ASAP7_75t_L g596 ( .A(n_520), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g602 ( .A(n_520), .Y(n_602) );
INVx2_ASAP7_75t_L g627 ( .A(n_520), .Y(n_627) );
AND2x2_ASAP7_75t_L g746 ( .A(n_520), .B(n_540), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_528), .B(n_579), .Y(n_666) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g539 ( .A(n_530), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
INVx2_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
AND2x4_ASAP7_75t_L g626 ( .A(n_530), .B(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_530), .Y(n_718) );
AOI22x1_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_547), .B1(n_565), .B2(n_570), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_539), .B(n_696), .C(n_697), .D(n_698), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_539), .B(n_596), .Y(n_726) );
INVx4_ASAP7_75t_SL g579 ( .A(n_540), .Y(n_579) );
BUFx2_ASAP7_75t_L g642 ( .A(n_540), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_540), .B(n_587), .Y(n_705) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g667 ( .A(n_549), .B(n_616), .Y(n_667) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g590 ( .A(n_553), .B(n_568), .Y(n_590) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_554), .B(n_569), .Y(n_614) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_564), .Y(n_554) );
OAI21x1_ASAP7_75t_L g609 ( .A1(n_555), .A2(n_556), .B(n_564), .Y(n_609) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_563), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_566), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g632 ( .A(n_566), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g671 ( .A(n_567), .B(n_589), .Y(n_671) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g714 ( .A(n_569), .B(n_624), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_570), .A2(n_687), .B1(n_689), .B2(n_692), .C(n_694), .Y(n_686) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g580 ( .A(n_572), .Y(n_580) );
OR2x2_ASAP7_75t_L g680 ( .A(n_572), .B(n_619), .Y(n_680) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_581), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_576), .A2(n_702), .B1(n_706), .B2(n_709), .Y(n_701) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
AND2x4_ASAP7_75t_L g625 ( .A(n_577), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g737 ( .A(n_577), .B(n_655), .Y(n_737) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g585 ( .A(n_579), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g601 ( .A(n_579), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g660 ( .A(n_579), .B(n_597), .Y(n_660) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_579), .Y(n_677) );
INVx1_ASAP7_75t_L g691 ( .A(n_579), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_579), .B(n_604), .Y(n_734) );
AND2x4_ASAP7_75t_L g641 ( .A(n_580), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g639 ( .A(n_582), .Y(n_639) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_583), .B(n_624), .Y(n_623) );
NAND2x1_ASAP7_75t_L g743 ( .A(n_583), .B(n_645), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B1(n_591), .B2(n_593), .Y(n_584) );
AND2x2_ASAP7_75t_L g610 ( .A(n_585), .B(n_603), .Y(n_610) );
INVx1_ASAP7_75t_L g651 ( .A(n_585), .Y(n_651) );
AND2x2_ASAP7_75t_L g758 ( .A(n_585), .B(n_619), .Y(n_758) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g591 ( .A(n_589), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g731 ( .A(n_589), .Y(n_731) );
AND2x2_ASAP7_75t_L g748 ( .A(n_589), .B(n_608), .Y(n_748) );
AND2x2_ASAP7_75t_L g764 ( .A(n_589), .B(n_714), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_590), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g687 ( .A(n_590), .B(n_688), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_590), .A2(n_680), .B1(n_695), .B2(n_699), .Y(n_694) );
INVx1_ASAP7_75t_L g650 ( .A(n_592), .Y(n_650) );
AND2x2_ASAP7_75t_L g681 ( .A(n_592), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_592), .B(n_688), .Y(n_710) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g716 ( .A(n_596), .B(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_596), .A2(n_620), .B1(n_725), .B2(n_727), .Y(n_724) );
INVx3_ASAP7_75t_L g619 ( .A(n_597), .Y(n_619) );
AND2x2_ASAP7_75t_L g751 ( .A(n_597), .B(n_604), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_615), .Y(n_598) );
AOI32xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_605), .A3(n_608), .B1(n_610), .B2(n_611), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_602), .Y(n_697) );
INVx1_ASAP7_75t_L g722 ( .A(n_602), .Y(n_722) );
INVx3_ASAP7_75t_L g678 ( .A(n_603), .Y(n_678) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_606), .A2(n_754), .B1(n_755), .B2(n_756), .C(n_757), .Y(n_753) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g730 ( .A(n_608), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g766 ( .A(n_608), .B(n_727), .Y(n_766) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g624 ( .A(n_609), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g638 ( .A(n_611), .B(n_639), .Y(n_638) );
AO22x1_ASAP7_75t_L g668 ( .A1(n_611), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_668) );
NAND2x1p5_ASAP7_75t_L g772 ( .A(n_611), .B(n_639), .Y(n_772) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g688 ( .A(n_612), .Y(n_688) );
INVx1_ASAP7_75t_L g698 ( .A(n_612), .Y(n_698) );
AND2x2_ASAP7_75t_L g618 ( .A(n_613), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_614), .Y(n_700) );
INVx1_ASAP7_75t_L g740 ( .A(n_614), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_620), .C(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2x1p5_ASAP7_75t_L g727 ( .A(n_617), .B(n_647), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_618), .B(n_677), .Y(n_754) );
AOI31xp33_ASAP7_75t_L g637 ( .A1(n_619), .A2(n_638), .A3(n_640), .B(n_643), .Y(n_637) );
INVx4_ASAP7_75t_L g696 ( .A(n_619), .Y(n_696) );
OR2x2_ASAP7_75t_L g733 ( .A(n_619), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x4_ASAP7_75t_L g635 ( .A(n_624), .B(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_626), .Y(n_631) );
AND2x2_ASAP7_75t_L g662 ( .A(n_626), .B(n_660), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_629), .B(n_637), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g755 ( .A(n_632), .Y(n_755) );
INVx1_ASAP7_75t_L g663 ( .A(n_633), .Y(n_663) );
AND2x4_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g693 ( .A(n_634), .Y(n_693) );
AND2x2_ASAP7_75t_L g692 ( .A(n_635), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI322xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .A3(n_652), .B1(n_656), .B2(n_659), .C1(n_661), .C2(n_663), .Y(n_649) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI211x1_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_668), .C(n_674), .Y(n_664) );
INVx1_ASAP7_75t_L g769 ( .A(n_665), .Y(n_769) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g723 ( .A(n_667), .Y(n_723) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OA21x2_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B(n_681), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx2_ASAP7_75t_L g744 ( .A(n_678), .Y(n_744) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_682), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_752), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_719), .C(n_735), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_701), .C(n_711), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_688), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g747 ( .A1(n_692), .A2(n_748), .B(n_749), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_696), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_696), .B(n_746), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_697), .B(n_771), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_698), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_708), .A2(n_758), .B(n_759), .Y(n_757) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_724), .C(n_728), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_SL g738 ( .A(n_730), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_734), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B(n_741), .C(n_747), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_746), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g767 ( .A(n_746), .Y(n_767) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g763 ( .A(n_751), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_761), .C(n_768), .Y(n_752) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI21xp33_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_765), .B(n_767), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AOI21xp33_ASAP7_75t_R g768 ( .A1(n_769), .A2(n_770), .B(n_772), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_774), .Y(n_780) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx5_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AND2x6_ASAP7_75t_SL g784 ( .A(n_785), .B(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_L g818 ( .A(n_786), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_786), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_789), .B(n_791), .Y(n_826) );
NOR3x1_ASAP7_75t_L g835 ( .A(n_789), .B(n_836), .C(n_839), .Y(n_835) );
AND2x6_ASAP7_75t_SL g804 ( .A(n_790), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_817), .B(n_819), .Y(n_792) );
OAI21xp33_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_798), .B(n_811), .Y(n_793) );
NAND2xp33_ASAP7_75t_L g811 ( .A(n_794), .B(n_812), .Y(n_811) );
AO21x1_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_803), .B(n_808), .Y(n_798) );
INVxp67_ASAP7_75t_SL g816 ( .A(n_799), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_800), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
INVx5_ASAP7_75t_L g810 ( .A(n_804), .Y(n_810) );
INVx3_ASAP7_75t_L g815 ( .A(n_804), .Y(n_815) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_808), .A2(n_813), .B(n_816), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx10_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
CKINVDCx6p67_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
BUFx12f_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
BUFx12f_ASAP7_75t_L g841 ( .A(n_830), .Y(n_841) );
AND2x6_ASAP7_75t_L g830 ( .A(n_831), .B(n_835), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVxp33_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
CKINVDCx14_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
endmodule