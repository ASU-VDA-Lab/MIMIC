module real_jpeg_1706_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_1),
.B(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_1),
.B(n_40),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_76),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_3),
.B(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_3),
.B(n_45),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_3),
.B(n_27),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_3),
.B(n_91),
.Y(n_257)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_40),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_34),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_56),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_4),
.B(n_30),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_4),
.B(n_27),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_5),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_5),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_45),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_5),
.B(n_91),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_6),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_45),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_8),
.B(n_34),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_8),
.B(n_56),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_8),
.B(n_30),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_8),
.B(n_27),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_8),
.B(n_45),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_91),
.Y(n_270)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_13),
.B(n_34),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_13),
.B(n_40),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_13),
.B(n_56),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_13),
.B(n_30),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_14),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_56),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_14),
.B(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_14),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_153),
.B1(n_348),
.B2(n_349),
.Y(n_17)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_18),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_152),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_124),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_21),
.B(n_124),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_21),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_59),
.CI(n_94),
.CON(n_21),
.SN(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_38),
.C(n_43),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_25),
.A2(n_26),
.B1(n_43),
.B2(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_26),
.B1(n_188),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_26),
.B(n_188),
.C(n_189),
.Y(n_187)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_27),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_28),
.A2(n_29),
.B1(n_67),
.B2(n_97),
.Y(n_170)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_29),
.B(n_67),
.C(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_48),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_40),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_43),
.A2(n_44),
.B1(n_90),
.B2(n_103),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_43),
.A2(n_44),
.B1(n_149),
.B2(n_228),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_88),
.C(n_90),
.Y(n_87)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_46),
.B(n_146),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.C(n_54),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_52),
.A2(n_53),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_53),
.B(n_135),
.C(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_56),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.C(n_69),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_62),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_65),
.B(n_69),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_80),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_117),
.C(n_119),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_81),
.B1(n_117),
.B2(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.C(n_93),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_87),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_102),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_90),
.A2(n_103),
.B1(n_245),
.B2(n_246),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_91),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_93),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_116),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_113),
.B1(n_122),
.B2(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.C(n_115),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_110),
.CI(n_115),
.CON(n_125),
.SN(n_125)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_106),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_96),
.B(n_100),
.Y(n_334)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B(n_104),
.C(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_101),
.A2(n_102),
.B1(n_184),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_103),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_105),
.A2(n_160),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_106),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_121),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_121),
.B(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.C(n_129),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_125),
.B(n_126),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_125),
.Y(n_350)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_129),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_142),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_130),
.A2(n_131),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_137),
.Y(n_131)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_132),
.B(n_134),
.CI(n_137),
.CON(n_310),
.SN(n_310)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_135),
.A2(n_136),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_135),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_136),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_140),
.B(n_142),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.C(n_151),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_143),
.A2(n_144),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_149),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_145),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_148),
.A2(n_149),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_149),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_150),
.A2(n_151),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_151),
.Y(n_322)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_153),
.Y(n_349)
);

OAI31xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_324),
.A3(n_337),
.B(n_342),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_304),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_229),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_201),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_157),
.B(n_201),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_171),
.C(n_191),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_158),
.B(n_301),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_158),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_163),
.CI(n_167),
.CON(n_158),
.SN(n_158)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_159),
.B(n_163),
.C(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_161),
.B(n_162),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_169),
.B(n_185),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_169),
.B(n_212),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_171),
.B(n_191),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_181),
.B2(n_190),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_182),
.C(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_178),
.C(n_180),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_199),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_192),
.B(n_195),
.CI(n_199),
.CON(n_291),
.SN(n_291)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_198),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_240),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_201),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_219),
.CI(n_220),
.CON(n_201),
.SN(n_201)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_202),
.B(n_219),
.C(n_220),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_203),
.B(n_206),
.C(n_213),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_213),
.B2(n_214),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_222),
.B(n_223),
.C(n_225),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_299),
.B(n_303),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_287),
.B(n_298),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_259),
.B(n_286),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_250),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_250),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_243),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_235),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_237),
.CI(n_238),
.CON(n_251),
.SN(n_251)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_239),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_248),
.C(n_249),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.C(n_258),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_283),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_251),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_253),
.B1(n_258),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_280),
.B(n_285),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_271),
.B(n_279),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_267),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_274),
.B(n_278),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_289),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_294),
.C(n_295),
.Y(n_302)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_291),
.Y(n_352)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_323),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_323),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_309),
.C(n_312),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_310),
.Y(n_357)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_317),
.C(n_318),
.Y(n_331)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g342 ( 
.A1(n_325),
.A2(n_338),
.B(n_343),
.C(n_346),
.D(n_347),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_335),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_332),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_341),
.Y(n_346)
);


endmodule