module real_aes_17332_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_0), .B(n_5), .C(n_21), .Y(n_20) );
NOR5xp2_ASAP7_75t_SL g18 ( .A(n_1), .B(n_8), .C(n_19), .D(n_23), .E(n_24), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_1), .Y(n_38) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_2), .B(n_4), .Y(n_27) );
NAND2xp33_ASAP7_75t_R g28 ( .A(n_2), .B(n_4), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g31 ( .A(n_2), .B(n_32), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_2), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_3), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_4), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_4), .B(n_35), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g44 ( .A1(n_6), .A2(n_15), .B1(n_27), .B2(n_34), .Y(n_44) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_7), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g43 ( .A(n_8), .Y(n_43) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_9), .Y(n_23) );
OAI22xp33_ASAP7_75t_SL g25 ( .A1(n_10), .A2(n_12), .B1(n_26), .B2(n_28), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_11), .Y(n_21) );
OAI22xp33_ASAP7_75t_SL g29 ( .A1(n_13), .A2(n_14), .B1(n_30), .B2(n_33), .Y(n_29) );
OAI32xp33_ASAP7_75t_L g16 ( .A1(n_17), .A2(n_25), .A3(n_29), .B1(n_36), .B2(n_44), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_19), .Y(n_42) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_22), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g39 ( .A(n_23), .B(n_40), .Y(n_39) );
NAND2xp33_ASAP7_75t_R g41 ( .A(n_24), .B(n_42), .Y(n_41) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_27), .Y(n_26) );
INVxp33_ASAP7_75t_SL g30 ( .A(n_31), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
NAND2xp33_ASAP7_75t_R g36 ( .A(n_37), .B(n_43), .Y(n_36) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_38), .B(n_39), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_41), .Y(n_40) );
endmodule