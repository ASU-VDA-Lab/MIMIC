module fake_jpeg_31379_n_337 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_337);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_17),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx9p33_ASAP7_75t_R g107 ( 
.A(n_45),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_51),
.Y(n_73)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_68),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_54),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_65),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_34),
.B(n_20),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_0),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_26),
.Y(n_105)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_37),
.B1(n_39),
.B2(n_38),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_82),
.A2(n_87),
.B1(n_96),
.B2(n_97),
.Y(n_143)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_44),
.B1(n_55),
.B2(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_88),
.B1(n_70),
.B2(n_30),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_37),
.B1(n_32),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_45),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_28),
.B1(n_27),
.B2(n_38),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_92),
.A2(n_106),
.B1(n_30),
.B2(n_3),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_32),
.B1(n_31),
.B2(n_42),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_42),
.B1(n_35),
.B2(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_113),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_114),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_36),
.B1(n_28),
.B2(n_20),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_41),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_53),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_47),
.B(n_29),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_60),
.B(n_36),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_25),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_123),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_67),
.C(n_65),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_136),
.C(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_126),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_16),
.C(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_124),
.B(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_132),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_61),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_17),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_29),
.B(n_25),
.C(n_16),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_138),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_86),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_30),
.B(n_29),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_97),
.B(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_141),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_25),
.B(n_2),
.C(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_1),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_145),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_1),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_84),
.B1(n_101),
.B2(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_1),
.Y(n_148)
);

OR2x2_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_5),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_5),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_152),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_5),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_78),
.B(n_76),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_102),
.Y(n_175)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_93),
.A3(n_76),
.B1(n_94),
.B2(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_160),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_94),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_186),
.C(n_157),
.Y(n_192)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_103),
.A3(n_84),
.B1(n_100),
.B2(n_74),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_127),
.B1(n_117),
.B2(n_146),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_181),
.Y(n_191)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_102),
.B1(n_95),
.B2(n_111),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_184),
.B1(n_12),
.B2(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_95),
.Y(n_181)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_74),
.B1(n_101),
.B2(n_7),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_190),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_149),
.B1(n_145),
.B2(n_142),
.Y(n_207)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_166),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_126),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_207),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_125),
.B1(n_144),
.B2(n_137),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_130),
.B(n_136),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_198),
.A2(n_199),
.B(n_187),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_130),
.B(n_141),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_130),
.B(n_119),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_215),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_165),
.B(n_139),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_129),
.B1(n_131),
.B2(n_120),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_139),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_139),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_120),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_133),
.Y(n_217)
);

NOR4xp25_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_169),
.C(n_183),
.D(n_161),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_221),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_175),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_181),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_234),
.C(n_221),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_231),
.B(n_199),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_166),
.C(n_189),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_232),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_192),
.B(n_180),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_169),
.B(n_164),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_213),
.B(n_172),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_174),
.C(n_190),
.Y(n_234)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_193),
.Y(n_253)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_202),
.B1(n_211),
.B2(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_235),
.B(n_247),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_260),
.B(n_264),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_259),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_235),
.B(n_226),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_241),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_194),
.C(n_191),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_228),
.C(n_234),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_193),
.B1(n_220),
.B2(n_191),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_263),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_227),
.B(n_205),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_200),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_273),
.C(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_277),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_233),
.C(n_223),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_240),
.C(n_231),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_242),
.B(n_241),
.C(n_203),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_210),
.C(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_258),
.C(n_248),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_295),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_212),
.B(n_207),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_275),
.B1(n_284),
.B2(n_272),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_296),
.B1(n_298),
.B2(n_200),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_259),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_251),
.B(n_261),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_263),
.B1(n_254),
.B2(n_247),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_273),
.B1(n_271),
.B2(n_252),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_250),
.C(n_253),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_268),
.B1(n_260),
.B2(n_267),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_266),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

NAND2x1p5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_267),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_200),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_276),
.B1(n_251),
.B2(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_303),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_308),
.B(n_294),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_216),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_309),
.B(n_290),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_278),
.C(n_252),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_292),
.C(n_288),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_244),
.B(n_237),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_208),
.B1(n_161),
.B2(n_171),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_208),
.B1(n_299),
.B2(n_287),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_292),
.C(n_288),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_306),
.C(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_197),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_316),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_318),
.Y(n_325)
);

AOI31xp67_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_208),
.A3(n_206),
.B(n_197),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_156),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_311),
.B(n_319),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_320),
.B(n_321),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_171),
.C(n_178),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_324),
.C(n_197),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_332),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_331),
.B(n_334),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_336),
.Y(n_337)
);


endmodule