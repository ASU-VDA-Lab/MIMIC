module fake_jpeg_437_n_681 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_681);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_681;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_60),
.Y(n_223)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_65),
.B(n_69),
.Y(n_140)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_67),
.B(n_78),
.Y(n_170)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_15),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_70),
.Y(n_149)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_74),
.Y(n_180)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_81),
.B(n_97),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_89),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_0),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_99),
.Y(n_222)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_101),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_48),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_104),
.B(n_113),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_36),
.B(n_1),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_45),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_116),
.B(n_121),
.Y(n_228)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_50),
.B(n_1),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_43),
.Y(n_184)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_45),
.B(n_2),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_20),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_122),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_129),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_30),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_32),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_131),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_32),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_69),
.A2(n_32),
.B1(n_58),
.B2(n_49),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_133),
.A2(n_166),
.B1(n_169),
.B2(n_179),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_134),
.B(n_153),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_60),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_75),
.B(n_58),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_160),
.B(n_173),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_118),
.A2(n_21),
.B1(n_57),
.B2(n_53),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_62),
.A2(n_59),
.B1(n_42),
.B2(n_46),
.Y(n_169)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_68),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_93),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_205),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_84),
.A2(n_35),
.B1(n_59),
.B2(n_46),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_88),
.B(n_21),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_182),
.B(n_193),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_5),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_110),
.A2(n_35),
.B1(n_53),
.B2(n_41),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_122),
.B1(n_105),
.B2(n_91),
.Y(n_233)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_111),
.B(n_37),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_190),
.B(n_3),
.Y(n_247)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_191),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_106),
.B(n_57),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_195),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_63),
.A2(n_35),
.B1(n_43),
.B2(n_37),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_196),
.A2(n_226),
.B1(n_187),
.B2(n_179),
.Y(n_242)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_197),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_41),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_204),
.Y(n_241)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_114),
.B(n_2),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_112),
.Y(n_205)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_95),
.Y(n_208)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_117),
.B(n_2),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_225),
.Y(n_250)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_102),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_218),
.Y(n_313)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_108),
.Y(n_220)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_2),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_73),
.A2(n_39),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_230),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_233),
.Y(n_350)
);

CKINVDCx12_ASAP7_75t_R g235 ( 
.A(n_147),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_235),
.Y(n_330)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_183),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_239),
.B(n_244),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_91),
.B(n_132),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_240),
.B(n_252),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_242),
.A2(n_265),
.B1(n_309),
.B2(n_141),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_145),
.B(n_90),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_243),
.B(n_247),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_96),
.B(n_39),
.C(n_40),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_87),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_245),
.B(n_251),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_140),
.B(n_82),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_246),
.B(n_248),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_165),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_170),
.B(n_4),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_138),
.B(n_80),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_253),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_252),
.Y(n_315)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_142),
.Y(n_256)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_257),
.Y(n_338)
);

CKINVDCx12_ASAP7_75t_R g258 ( 
.A(n_147),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_6),
.B(n_7),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_259),
.B(n_279),
.Y(n_354)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_262),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_263),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_226),
.A2(n_76),
.B1(n_39),
.B2(n_40),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_171),
.Y(n_267)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_267),
.Y(n_363)
);

OR2x2_ASAP7_75t_SL g268 ( 
.A(n_135),
.B(n_39),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_268),
.B(n_214),
.C(n_151),
.Y(n_345)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_269),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_6),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_271),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_152),
.B(n_6),
.Y(n_271)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_171),
.Y(n_272)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_272),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_149),
.Y(n_273)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_154),
.B(n_7),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_275),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_156),
.B(n_7),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_139),
.A2(n_7),
.B(n_8),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_277),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_161),
.B(n_8),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_280),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_139),
.A2(n_8),
.B(n_9),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_163),
.B(n_9),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_189),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_285),
.Y(n_348)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_146),
.B(n_158),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_147),
.B(n_9),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_286),
.B(n_290),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_155),
.Y(n_288)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_148),
.B(n_10),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_155),
.Y(n_291)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_202),
.Y(n_292)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_180),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_297),
.B(n_298),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_144),
.B(n_10),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_299),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_185),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

CKINVDCx9p33_ASAP7_75t_R g302 ( 
.A(n_196),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_302),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_159),
.B(n_11),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_217),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_304),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_305),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_206),
.B(n_11),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_306),
.Y(n_364)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_157),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_168),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_308),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_162),
.A2(n_194),
.B1(n_176),
.B2(n_164),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_180),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_151),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_192),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_312),
.A2(n_214),
.B1(n_141),
.B2(n_219),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_315),
.B(n_259),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_254),
.B(n_194),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_321),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_250),
.B(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_192),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_332),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_328),
.A2(n_340),
.B1(n_344),
.B2(n_351),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_231),
.B(n_176),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_241),
.B(n_222),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_342),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_302),
.A2(n_164),
.B1(n_203),
.B2(n_186),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_252),
.B(n_224),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_232),
.A2(n_186),
.B1(n_203),
.B2(n_157),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_345),
.B(n_249),
.C(n_284),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_240),
.B(n_174),
.C(n_220),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_371),
.C(n_374),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_246),
.A2(n_236),
.B1(n_242),
.B2(n_244),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_265),
.A2(n_174),
.B1(n_200),
.B2(n_219),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_365),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_253),
.A2(n_177),
.B1(n_143),
.B2(n_167),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_367),
.A2(n_261),
.B1(n_288),
.B2(n_291),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_253),
.B(n_177),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_283),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_234),
.B(n_221),
.C(n_229),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_255),
.B(n_276),
.C(n_281),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_277),
.B1(n_279),
.B2(n_167),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_377),
.A2(n_393),
.B1(n_367),
.B2(n_373),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_270),
.B(n_297),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_378),
.A2(n_319),
.B(n_368),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_321),
.B(n_295),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_381),
.B(n_386),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_238),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_313),
.C(n_301),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_383),
.B(n_402),
.C(n_414),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_310),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_324),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_387),
.B(n_389),
.Y(n_447)
);

AO22x2_ASAP7_75t_SL g388 ( 
.A1(n_341),
.A2(n_309),
.B1(n_273),
.B2(n_301),
.Y(n_388)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_263),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_390),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_391),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_323),
.B(n_313),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_394),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_328),
.A2(n_137),
.B1(n_143),
.B2(n_307),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_372),
.B(n_260),
.Y(n_394)
);

BUFx12f_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_403),
.Y(n_439)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_396),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_230),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_397),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_333),
.B(n_237),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_399),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_324),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_311),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_400),
.B(n_401),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_330),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_314),
.B(n_349),
.C(n_315),
.Y(n_402)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_410),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_371),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_406),
.A2(n_353),
.B1(n_346),
.B2(n_326),
.Y(n_463)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_361),
.A2(n_304),
.B(n_293),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_408),
.A2(n_373),
.B(n_331),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_332),
.Y(n_409)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_409),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_316),
.B(n_264),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_337),
.B1(n_357),
.B2(n_318),
.Y(n_451)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_412),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_348),
.B(n_260),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_418),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_314),
.B(n_264),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_362),
.A2(n_269),
.B1(n_292),
.B2(n_256),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_415),
.A2(n_262),
.B1(n_331),
.B2(n_369),
.Y(n_437)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_417),
.Y(n_441)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_335),
.Y(n_423)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_345),
.B(n_294),
.C(n_287),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_374),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_327),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_SL g501 ( 
.A(n_427),
.B(n_435),
.Y(n_501)
);

OAI32xp33_ASAP7_75t_L g430 ( 
.A1(n_376),
.A2(n_355),
.A3(n_325),
.B1(n_370),
.B2(n_354),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_376),
.A2(n_354),
.B1(n_350),
.B2(n_355),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_431),
.A2(n_433),
.B1(n_377),
.B2(n_379),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_380),
.A2(n_354),
.B1(n_350),
.B2(n_360),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_436),
.A2(n_450),
.B1(n_457),
.B2(n_388),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_442),
.A2(n_464),
.B(n_417),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_385),
.A2(n_334),
.B1(n_342),
.B2(n_317),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_SL g486 ( 
.A1(n_451),
.A2(n_416),
.B(n_388),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_317),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_455),
.B(n_423),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_356),
.B1(n_336),
.B2(n_326),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_408),
.A2(n_357),
.B(n_356),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_458),
.A2(n_405),
.B(n_414),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_402),
.C(n_379),
.Y(n_472)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_421),
.Y(n_461)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_461),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_439),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_378),
.A2(n_353),
.B(n_346),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_466),
.A2(n_482),
.B1(n_492),
.B2(n_497),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_467),
.A2(n_485),
.B(n_490),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_452),
.B(n_401),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_468),
.B(n_470),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_392),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_431),
.C(n_448),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_426),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_475),
.Y(n_509)
);

OA22x2_ASAP7_75t_L g474 ( 
.A1(n_428),
.A2(n_411),
.B1(n_388),
.B2(n_420),
.Y(n_474)
);

AOI22x1_ASAP7_75t_L g540 ( 
.A1(n_474),
.A2(n_445),
.B1(n_363),
.B2(n_375),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_426),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_429),
.Y(n_476)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_383),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_480),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_425),
.B(n_438),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_481),
.B(n_495),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_428),
.A2(n_404),
.B1(n_420),
.B2(n_410),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_424),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_483),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_412),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_484),
.B(n_487),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_494),
.B1(n_502),
.B2(n_459),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_438),
.B(n_425),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_448),
.A2(n_381),
.B(n_422),
.C(n_407),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_496),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_489),
.Y(n_506)
);

HAxp5_ASAP7_75t_SL g490 ( 
.A(n_453),
.B(n_396),
.CON(n_490),
.SN(n_490)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_491),
.A2(n_447),
.B(n_444),
.Y(n_518)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_441),
.Y(n_493)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_436),
.A2(n_416),
.B1(n_423),
.B2(n_399),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_427),
.B(n_419),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_450),
.A2(n_427),
.B1(n_432),
.B2(n_453),
.Y(n_497)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_447),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_445),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_460),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_466),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_455),
.B(n_387),
.Y(n_500)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_500),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_433),
.A2(n_390),
.B1(n_336),
.B2(n_318),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_440),
.B(n_390),
.Y(n_503)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_499),
.B(n_465),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_505),
.B(n_483),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_507),
.B(n_512),
.C(n_525),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_501),
.A2(n_458),
.B(n_442),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_508),
.A2(n_518),
.B(n_520),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_463),
.C(n_440),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_432),
.Y(n_513)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_513),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_494),
.A2(n_451),
.B1(n_444),
.B2(n_439),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_519),
.A2(n_523),
.B1(n_529),
.B2(n_530),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_501),
.A2(n_479),
.B(n_485),
.Y(n_520)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_477),
.Y(n_522)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_522),
.Y(n_567)
);

OAI22x1_ASAP7_75t_L g524 ( 
.A1(n_482),
.A2(n_439),
.B1(n_430),
.B2(n_443),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_524),
.A2(n_483),
.B1(n_480),
.B2(n_502),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_481),
.B(n_434),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_526),
.B(n_491),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_479),
.A2(n_475),
.B1(n_473),
.B2(n_500),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_503),
.A2(n_441),
.B1(n_461),
.B2(n_449),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_467),
.A2(n_449),
.B1(n_446),
.B2(n_459),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_531),
.A2(n_540),
.B1(n_474),
.B2(n_456),
.Y(n_564)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_490),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_SL g568 ( 
.A(n_534),
.B(n_403),
.C(n_375),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_469),
.B(n_446),
.Y(n_536)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_536),
.Y(n_552)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_493),
.Y(n_543)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_543),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_509),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_544),
.B(n_547),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_551),
.Y(n_576)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_509),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_513),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_548),
.B(n_549),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_536),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_512),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_507),
.B(n_480),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_553),
.B(n_557),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_522),
.B(n_471),
.Y(n_554)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_556),
.A2(n_532),
.B1(n_539),
.B2(n_514),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_505),
.B(n_529),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_476),
.C(n_474),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_537),
.C(n_518),
.Y(n_573)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_560),
.Y(n_585)
);

AND3x1_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_474),
.C(n_478),
.Y(n_561)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_561),
.Y(n_580)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_562),
.Y(n_586)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_504),
.Y(n_563)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_563),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_564),
.A2(n_523),
.B1(n_524),
.B2(n_531),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_391),
.Y(n_565)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_565),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_514),
.A2(n_443),
.B(n_456),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_566),
.A2(n_535),
.B(n_517),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_508),
.B(n_489),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_570),
.B(n_540),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_532),
.B(n_510),
.Y(n_571)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_571),
.Y(n_596)
);

NOR2x1_ASAP7_75t_L g572 ( 
.A(n_510),
.B(n_395),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_572),
.A2(n_515),
.B(n_534),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_573),
.B(n_597),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_516),
.C(n_527),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_583),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_591),
.B1(n_556),
.B2(n_558),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_543),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_587),
.Y(n_612)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_589),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_559),
.A2(n_515),
.B1(n_540),
.B2(n_533),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_552),
.Y(n_610)
);

AO21x1_ASAP7_75t_L g615 ( 
.A1(n_594),
.A2(n_596),
.B(n_585),
.Y(n_615)
);

AOI21xp33_ASAP7_75t_L g595 ( 
.A1(n_569),
.A2(n_511),
.B(n_506),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_595),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_557),
.B(n_443),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_555),
.B(n_363),
.C(n_338),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_598),
.B(n_551),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_599),
.A2(n_506),
.B1(n_329),
.B2(n_352),
.Y(n_637)
);

AOI321xp33_ASAP7_75t_L g600 ( 
.A1(n_574),
.A2(n_569),
.A3(n_568),
.B1(n_541),
.B2(n_552),
.C(n_572),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g625 ( 
.A(n_600),
.Y(n_625)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_579),
.Y(n_603)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_603),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_604),
.B(n_618),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_553),
.C(n_545),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_605),
.B(n_606),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_575),
.B(n_570),
.C(n_566),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_594),
.Y(n_607)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_607),
.Y(n_623)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_577),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_608),
.B(n_609),
.Y(n_635)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_581),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_615),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_593),
.B(n_542),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_611),
.A2(n_616),
.B(n_550),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_554),
.C(n_541),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_613),
.B(n_614),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_576),
.C(n_573),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_578),
.B(n_571),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_591),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_589),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_622),
.B(n_624),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_602),
.A2(n_584),
.B1(n_582),
.B2(n_580),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_576),
.C(n_597),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_628),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_619),
.B(n_587),
.C(n_580),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_619),
.B(n_592),
.C(n_567),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_629),
.B(n_352),
.C(n_359),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_567),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_630),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_612),
.A2(n_588),
.B1(n_586),
.B2(n_561),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_636),
.Y(n_642)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_633),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_606),
.B(n_601),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_637),
.A2(n_610),
.B1(n_600),
.B2(n_615),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_634),
.A2(n_612),
.B(n_617),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_639),
.B(n_641),
.Y(n_654)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_640),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_632),
.B(n_395),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_645),
.B(n_646),
.Y(n_655)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_627),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_625),
.A2(n_359),
.B1(n_343),
.B2(n_395),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_647),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_626),
.B(n_343),
.C(n_249),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_648),
.B(n_649),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_L g649 ( 
.A1(n_625),
.A2(n_289),
.B(n_287),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_623),
.A2(n_627),
.B(n_622),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_650),
.B(n_651),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_636),
.A2(n_137),
.B1(n_305),
.B2(n_266),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_648),
.B(n_628),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_653),
.B(n_662),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_643),
.A2(n_620),
.B(n_635),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_657),
.A2(n_650),
.B(n_642),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_630),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_661),
.B(n_621),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_629),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_652),
.B(n_621),
.C(n_284),
.Y(n_663)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_663),
.B(n_649),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_664),
.B(n_667),
.C(n_660),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_638),
.C(n_641),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_665),
.B(n_666),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_654),
.B(n_647),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_668),
.B(n_669),
.C(n_663),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_655),
.B(n_257),
.C(n_289),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_671),
.B(n_674),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_672),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_670),
.B(n_659),
.C(n_658),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_675),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_677),
.B(n_670),
.C(n_673),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_678),
.A2(n_659),
.B1(n_267),
.B2(n_272),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_266),
.Y(n_680)
);

AO21x1_ASAP7_75t_L g681 ( 
.A1(n_680),
.A2(n_305),
.B(n_294),
.Y(n_681)
);


endmodule