module fake_jpeg_13916_n_546 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_546);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_58),
.Y(n_132)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_60),
.Y(n_135)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_65),
.B(n_87),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_15),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_41),
.B(n_75),
.C(n_24),
.Y(n_121)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_43),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_81),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_17),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_20),
.B(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_101),
.Y(n_129)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_24),
.Y(n_139)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_45),
.B1(n_39),
.B2(n_50),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_118),
.A2(n_136),
.B1(n_163),
.B2(n_42),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_121),
.B(n_125),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_66),
.A2(n_44),
.B(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_56),
.A2(n_46),
.B1(n_26),
.B2(n_45),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_24),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_141),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_24),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_23),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_144),
.B(n_91),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_63),
.A2(n_26),
.B1(n_50),
.B2(n_42),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_149),
.A2(n_21),
.B1(n_85),
.B2(n_83),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_75),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_41),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_104),
.Y(n_190)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_69),
.A2(n_50),
.B1(n_42),
.B2(n_44),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_178),
.Y(n_234)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_173),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_161),
.Y(n_175)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_88),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_177),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_100),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_199),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_180),
.Y(n_274)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_183),
.Y(n_245)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_108),
.B(n_23),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_188),
.B(n_197),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_190),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

OR2x4_ASAP7_75t_L g195 ( 
.A(n_112),
.B(n_104),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_226),
.Y(n_229)
);

CKINVDCx9p33_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_196),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_86),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_92),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_198),
.B(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_33),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_33),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_48),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_204),
.B(n_210),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_147),
.B1(n_138),
.B2(n_128),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_118),
.A2(n_90),
.B1(n_76),
.B2(n_79),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_206),
.A2(n_162),
.B1(n_119),
.B2(n_111),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_135),
.B(n_99),
.C(n_72),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_119),
.B1(n_162),
.B2(n_128),
.Y(n_247)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_38),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_126),
.B(n_38),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_211),
.B(n_213),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_91),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_212),
.B(n_214),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_0),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_133),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_62),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_219),
.Y(n_270)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_218),
.Y(n_273)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_142),
.B(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_221),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_62),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_145),
.B(n_21),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_160),
.C(n_146),
.Y(n_263)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

BUFx8_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_153),
.B(n_0),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_224),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_225),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_134),
.B(n_0),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_172),
.A2(n_82),
.B1(n_164),
.B2(n_111),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_236),
.A2(n_247),
.B1(n_259),
.B2(n_265),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_249),
.B1(n_196),
.B2(n_216),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_113),
.B(n_117),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_198),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_168),
.B(n_113),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_262),
.C(n_177),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_172),
.A2(n_147),
.B1(n_138),
.B2(n_143),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_143),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_254),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_211),
.A2(n_36),
.B1(n_160),
.B2(n_3),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_277),
.A2(n_279),
.B1(n_305),
.B2(n_177),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_278),
.A2(n_309),
.B(n_321),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_229),
.A2(n_205),
.B1(n_207),
.B2(n_206),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_188),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_280),
.B(n_283),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_180),
.B1(n_204),
.B2(n_171),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_189),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_284),
.Y(n_333)
);

OR2x2_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_195),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_320),
.C(n_223),
.Y(n_351)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_270),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_288),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_201),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_312),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_202),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_293),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_179),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_301),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_173),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_298),
.Y(n_332)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_272),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_299),
.B(n_300),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_239),
.B(n_235),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_307),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_239),
.B(n_192),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_311),
.Y(n_343)
);

AO21x2_ASAP7_75t_L g304 ( 
.A1(n_243),
.A2(n_182),
.B(n_209),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_257),
.B1(n_274),
.B2(n_182),
.Y(n_338)
);

OAI22x1_ASAP7_75t_SL g305 ( 
.A1(n_229),
.A2(n_263),
.B1(n_259),
.B2(n_254),
.Y(n_305)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_232),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_253),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_313),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_236),
.B(n_169),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_268),
.A2(n_175),
.B1(n_200),
.B2(n_198),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_310),
.A2(n_317),
.B1(n_203),
.B2(n_217),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_234),
.B(n_175),
.Y(n_311)
);

INVx2_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_238),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_319),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_176),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_318),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_231),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_316),
.A2(n_313),
.B(n_306),
.Y(n_354)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_231),
.B(n_181),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_184),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_238),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_325),
.A2(n_327),
.B1(n_348),
.B2(n_358),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_309),
.A2(n_186),
.B1(n_273),
.B2(n_242),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_326),
.A2(n_334),
.B1(n_335),
.B2(n_347),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_279),
.A2(n_305),
.B1(n_278),
.B2(n_315),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_295),
.A2(n_242),
.B1(n_244),
.B2(n_258),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_218),
.B1(n_244),
.B2(n_258),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_338),
.B(n_360),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_278),
.A2(n_274),
.B1(n_256),
.B2(n_264),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_350),
.B(n_354),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_293),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_346),
.B(n_304),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_304),
.A2(n_170),
.B1(n_193),
.B2(n_187),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_277),
.A2(n_264),
.B1(n_252),
.B2(n_261),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_285),
.A2(n_245),
.B(n_219),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_174),
.C(n_304),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_290),
.B(n_297),
.C(n_291),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_355),
.C(n_357),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_237),
.C(n_252),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_185),
.C(n_174),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_292),
.A2(n_261),
.B1(n_191),
.B2(n_271),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_316),
.A2(n_160),
.B1(n_194),
.B2(n_271),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_359),
.A2(n_354),
.B(n_341),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_282),
.A2(n_288),
.B(n_284),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_286),
.Y(n_363)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_304),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_364),
.A2(n_396),
.B(n_359),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_302),
.Y(n_365)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_360),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_343),
.B(n_307),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_372),
.Y(n_399)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_361),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_344),
.B(n_317),
.Y(n_372)
);

BUFx16f_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_353),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_385),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_327),
.Y(n_398)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_298),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_376),
.B(n_394),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_378),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_362),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_324),
.B(n_346),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_380),
.B(n_383),
.C(n_350),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_323),
.B(n_318),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_381),
.B(n_384),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_329),
.B(n_301),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_390),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_294),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_296),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_340),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_387),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_340),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_321),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_392),
.Y(n_407)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_314),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_375),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_362),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_339),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_398),
.B(n_403),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_325),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_404),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_379),
.Y(n_404)
);

XOR2x2_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_373),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_397),
.A2(n_331),
.B1(n_348),
.B2(n_355),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_411),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_416),
.B(n_418),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_347),
.B1(n_349),
.B2(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_393),
.A2(n_376),
.B(n_368),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_393),
.A2(n_368),
.B(n_396),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_366),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_420),
.B(n_424),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_351),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_428),
.C(n_429),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_335),
.B1(n_334),
.B2(n_326),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_423),
.A2(n_426),
.B1(n_388),
.B2(n_377),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_357),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_333),
.B1(n_349),
.B2(n_345),
.Y(n_425)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_425),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_389),
.A2(n_333),
.B1(n_345),
.B2(n_338),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_387),
.B(n_339),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_427),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_361),
.C(n_336),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_399),
.B(n_365),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_436),
.B(n_438),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_437),
.A2(n_447),
.B1(n_414),
.B2(n_406),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_401),
.B(n_390),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_418),
.A2(n_393),
.B(n_386),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_439),
.A2(n_441),
.B(n_446),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_421),
.A2(n_364),
.B(n_395),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_422),
.C(n_402),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_448),
.C(n_451),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_394),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_453),
.Y(n_471)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_385),
.B(n_388),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_420),
.A2(n_371),
.B1(n_338),
.B2(n_392),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_408),
.C(n_429),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_417),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_452),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_434),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_SL g451 ( 
.A(n_410),
.B(n_338),
.C(n_373),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_260),
.C(n_36),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_413),
.C(n_412),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_413),
.Y(n_454)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_454),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_260),
.C(n_2),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_407),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_456),
.B(n_403),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_426),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_460),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_464),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_453),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_431),
.A2(n_423),
.B1(n_400),
.B2(n_421),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_467),
.B1(n_450),
.B2(n_441),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_437),
.A2(n_409),
.B1(n_419),
.B2(n_414),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_473),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_433),
.A2(n_440),
.B1(n_419),
.B2(n_443),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_425),
.Y(n_468)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_405),
.Y(n_470)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_455),
.Y(n_472)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_405),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_478),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_411),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_458),
.A2(n_448),
.B1(n_451),
.B2(n_447),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_479),
.A2(n_481),
.B1(n_488),
.B2(n_464),
.Y(n_497)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_458),
.A2(n_435),
.B1(n_442),
.B2(n_430),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_430),
.C(n_444),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_469),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_462),
.A2(n_477),
.B1(n_461),
.B2(n_468),
.Y(n_488)
);

AOI322xp5_ASAP7_75t_L g489 ( 
.A1(n_474),
.A2(n_406),
.A3(n_446),
.B1(n_435),
.B2(n_456),
.C1(n_439),
.C2(n_452),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_489),
.B(n_475),
.Y(n_503)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_471),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_491),
.B(n_470),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_475),
.A2(n_260),
.B(n_2),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_1),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_494),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_498),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_497),
.A2(n_484),
.B1(n_6),
.B2(n_7),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_473),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_476),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_500),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_457),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_457),
.C(n_466),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_501),
.A2(n_503),
.B(n_507),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_504),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_486),
.A2(n_478),
.B1(n_459),
.B2(n_3),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_510),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_1),
.C(n_2),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_13),
.C(n_3),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_511),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_3),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_487),
.A2(n_5),
.B(n_6),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_483),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_514),
.A2(n_506),
.B(n_508),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_483),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_517),
.C(n_516),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_490),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_R g521 ( 
.A(n_507),
.B(n_492),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_521),
.B(n_505),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_509),
.Y(n_526)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_512),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_526),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_527),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_5),
.B(n_7),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_529),
.C(n_530),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_515),
.B(n_7),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_520),
.B(n_513),
.C(n_517),
.Y(n_531)
);

FAx1_ASAP7_75t_SL g532 ( 
.A(n_531),
.B(n_522),
.CI(n_516),
.CON(n_532),
.SN(n_532)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_532),
.A2(n_524),
.B(n_519),
.Y(n_537)
);

AOI322xp5_ASAP7_75t_L g540 ( 
.A1(n_537),
.A2(n_538),
.A3(n_539),
.B1(n_536),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_518),
.B(n_9),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_535),
.A2(n_8),
.B(n_9),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_541),
.C(n_10),
.Y(n_542)
);

AOI322xp5_ASAP7_75t_L g541 ( 
.A1(n_537),
.A2(n_534),
.A3(n_532),
.B1(n_533),
.B2(n_12),
.C1(n_9),
.C2(n_11),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_10),
.B(n_11),
.Y(n_543)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_543),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_10),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_545),
.Y(n_546)
);


endmodule