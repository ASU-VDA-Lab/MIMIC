module fake_jpeg_7442_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx9p33_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_0),
.C(n_1),
.Y(n_19)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_19),
.C(n_22),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_10),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_18),
.B1(n_16),
.B2(n_9),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_27),
.B2(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_15),
.B1(n_20),
.B2(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_14),
.B1(n_12),
.B2(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_27),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_0),
.B(n_2),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_41),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_42),
.A3(n_44),
.B1(n_6),
.B2(n_3),
.C1(n_5),
.C2(n_17),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_43),
.C(n_4),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_3),
.B1(n_5),
.B2(n_17),
.Y(n_51)
);


endmodule