module real_aes_7017_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_816;
wire n_400;
wire n_539;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_0), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_1), .Y(n_593) );
XOR2x2_ASAP7_75t_L g660 ( .A(n_2), .B(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_3), .A2(n_230), .B1(n_339), .B2(n_342), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_4), .A2(n_175), .B1(n_399), .B2(n_402), .Y(n_738) );
INVx1_ASAP7_75t_L g314 ( .A(n_5), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_6), .A2(n_59), .B1(n_395), .B2(n_396), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_7), .A2(n_185), .B1(n_383), .B2(n_619), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_8), .Y(n_542) );
INVx1_ASAP7_75t_L g733 ( .A(n_9), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_10), .A2(n_115), .B1(n_339), .B2(n_342), .C(n_345), .Y(n_338) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_11), .A2(n_31), .B1(n_222), .B2(n_358), .C1(n_569), .C2(n_575), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_12), .A2(n_246), .B1(n_324), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_13), .A2(n_173), .B1(n_287), .B2(n_376), .Y(n_434) );
INVx1_ASAP7_75t_L g520 ( .A(n_14), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_15), .B(n_422), .Y(n_736) );
OA22x2_ASAP7_75t_L g481 ( .A1(n_16), .A2(n_482), .B1(n_483), .B2(n_521), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_16), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_17), .A2(n_147), .B1(n_437), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_18), .A2(n_76), .B1(n_303), .B2(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_19), .A2(n_239), .B1(n_319), .B2(n_324), .C(n_328), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_20), .Y(n_841) );
INVx1_ASAP7_75t_L g346 ( .A(n_21), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_22), .A2(n_72), .B1(n_286), .B2(n_303), .C(n_307), .Y(n_285) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_23), .A2(n_34), .B1(n_247), .B2(n_358), .C1(n_360), .C2(n_364), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_24), .Y(n_638) );
XOR2x2_ASAP7_75t_L g679 ( .A(n_25), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g406 ( .A(n_26), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_27), .A2(n_94), .B1(n_457), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_28), .A2(n_79), .B1(n_473), .B2(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_29), .A2(n_259), .B1(n_478), .B2(n_858), .Y(n_857) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_30), .A2(n_83), .B1(n_292), .B2(n_297), .Y(n_300) );
INVx1_ASAP7_75t_L g787 ( .A(n_30), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_32), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_33), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_35), .A2(n_186), .B1(n_365), .B2(n_408), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_36), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_37), .A2(n_53), .B1(n_286), .B2(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g518 ( .A(n_38), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_39), .A2(n_43), .B1(n_395), .B2(n_422), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_40), .A2(n_206), .B1(n_327), .B2(n_376), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_41), .Y(n_543) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_42), .A2(n_87), .B1(n_292), .B2(n_293), .Y(n_302) );
INVx1_ASAP7_75t_L g788 ( .A(n_42), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_44), .A2(n_135), .B1(n_746), .B2(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g509 ( .A(n_45), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_46), .A2(n_120), .B1(n_303), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_47), .A2(n_48), .B1(n_335), .B2(n_499), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_49), .Y(n_601) );
INVx1_ASAP7_75t_L g492 ( .A(n_50), .Y(n_492) );
INVx1_ASAP7_75t_L g505 ( .A(n_51), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_52), .A2(n_256), .B1(n_568), .B2(n_569), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_54), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_55), .A2(n_151), .B1(n_471), .B2(n_472), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_56), .B(n_395), .Y(n_420) );
INVx1_ASAP7_75t_L g728 ( .A(n_57), .Y(n_728) );
AOI22xp5_ASAP7_75t_SL g378 ( .A1(n_58), .A2(n_253), .B1(n_379), .B2(n_383), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_60), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_61), .A2(n_197), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_62), .A2(n_233), .B1(n_617), .B2(n_704), .Y(n_703) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_63), .B(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_64), .A2(n_208), .B1(n_468), .B2(n_636), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_65), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_66), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_67), .B(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_68), .A2(n_249), .B1(n_398), .B2(n_401), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_69), .A2(n_205), .B1(n_287), .B2(n_468), .Y(n_673) );
OA22x2_ASAP7_75t_L g445 ( .A1(n_70), .A2(n_446), .B1(n_447), .B2(n_479), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_70), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_71), .A2(n_255), .B1(n_365), .B2(n_424), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_73), .B(n_339), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_74), .A2(n_791), .B1(n_823), .B2(n_824), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_74), .Y(n_823) );
INVx1_ASAP7_75t_L g659 ( .A(n_75), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_77), .A2(n_154), .B1(n_417), .B2(n_418), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_78), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_80), .A2(n_160), .B1(n_319), .B2(n_640), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_81), .A2(n_99), .B1(n_747), .B2(n_762), .Y(n_761) );
AO22x1_ASAP7_75t_L g752 ( .A1(n_82), .A2(n_753), .B1(n_754), .B2(n_771), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_82), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_84), .A2(n_179), .B1(n_478), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_85), .A2(n_90), .B1(n_402), .B2(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_86), .A2(n_224), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_88), .A2(n_210), .B1(n_428), .B2(n_430), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_89), .A2(n_204), .B1(n_389), .B2(n_392), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_91), .A2(n_149), .B1(n_384), .B2(n_468), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_92), .Y(n_815) );
INVx1_ASAP7_75t_L g833 ( .A(n_93), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_93), .A2(n_833), .B1(n_835), .B2(n_860), .Y(n_834) );
INVx1_ASAP7_75t_L g278 ( .A(n_95), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_96), .A2(n_128), .B1(n_578), .B2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_97), .A2(n_139), .B1(n_585), .B2(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_98), .B(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_100), .A2(n_187), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_101), .Y(n_596) );
INVx1_ASAP7_75t_L g274 ( .A(n_102), .Y(n_274) );
INVx1_ASAP7_75t_L g409 ( .A(n_103), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_104), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_105), .A2(n_184), .B1(n_619), .B2(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_106), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_107), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_108), .A2(n_152), .B1(n_428), .B2(n_640), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_109), .A2(n_234), .B1(n_376), .B2(n_384), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_110), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_111), .A2(n_192), .B1(n_498), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_112), .A2(n_223), .B1(n_615), .B2(n_852), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_113), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_114), .Y(n_711) );
AOI222xp33_ASAP7_75t_L g770 ( .A1(n_116), .A2(n_148), .B1(n_257), .B2(n_358), .C1(n_364), .C2(n_424), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_117), .A2(n_167), .B1(n_360), .B2(n_365), .Y(n_715) );
AOI222xp33_ASAP7_75t_L g553 ( .A1(n_118), .A2(n_132), .B1(n_215), .B2(n_554), .C1(n_555), .C2(n_556), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_119), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_121), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_122), .A2(n_217), .B1(n_463), .B2(n_464), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_123), .A2(n_131), .B1(n_360), .B2(n_665), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_124), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_125), .A2(n_178), .B1(n_383), .B2(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_126), .A2(n_284), .B1(n_368), .B2(n_369), .Y(n_283) );
INVx1_ASAP7_75t_L g368 ( .A(n_126), .Y(n_368) );
INVx1_ASAP7_75t_L g351 ( .A(n_127), .Y(n_351) );
AO22x2_ASAP7_75t_L g525 ( .A1(n_129), .A2(n_526), .B1(n_557), .B2(n_558), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_129), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_130), .A2(n_141), .B1(n_546), .B2(n_548), .C(n_549), .Y(n_545) );
INVx1_ASAP7_75t_L g486 ( .A(n_133), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_134), .A2(n_263), .B1(n_428), .B2(n_436), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_136), .A2(n_201), .B1(n_585), .B2(n_612), .Y(n_856) );
INVx1_ASAP7_75t_L g329 ( .A(n_137), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_138), .A2(n_172), .B1(n_615), .B2(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_140), .B(n_555), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_142), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_143), .A2(n_245), .B1(n_398), .B2(n_555), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_144), .A2(n_196), .B1(n_475), .B2(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_145), .A2(n_168), .B1(n_383), .B2(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g308 ( .A(n_146), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_150), .Y(n_842) );
AND2x2_ASAP7_75t_L g277 ( .A(n_153), .B(n_278), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_155), .A2(n_268), .B1(n_335), .B2(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_156), .A2(n_241), .B1(n_417), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_157), .A2(n_269), .B1(n_424), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_158), .A2(n_161), .B1(n_475), .B2(n_477), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_159), .A2(n_262), .B1(n_580), .B2(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g333 ( .A(n_162), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_163), .A2(n_218), .B1(n_619), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_164), .A2(n_264), .B1(n_383), .B2(n_467), .Y(n_466) );
AND2x6_ASAP7_75t_L g273 ( .A(n_165), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_165), .Y(n_781) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_166), .A2(n_229), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_169), .A2(n_227), .B1(n_547), .B2(n_548), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_170), .Y(n_839) );
INVx1_ASAP7_75t_L g438 ( .A(n_171), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_174), .A2(n_228), .B1(n_465), .B2(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_176), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_177), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_180), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_181), .Y(n_845) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_182), .A2(n_271), .B(n_279), .C(n_789), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_183), .A2(n_235), .B1(n_428), .B2(n_463), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_188), .A2(n_213), .B1(n_608), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_189), .A2(n_220), .B1(n_303), .B2(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_190), .B(n_422), .Y(n_421) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_191), .A2(n_243), .B1(n_292), .B2(n_297), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_193), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_194), .A2(n_244), .B1(n_610), .B2(n_727), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_195), .B(n_396), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_198), .A2(n_200), .B1(n_432), .B2(n_468), .Y(n_742) );
INVx1_ASAP7_75t_L g517 ( .A(n_199), .Y(n_517) );
INVx1_ASAP7_75t_L g718 ( .A(n_202), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_203), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_207), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_209), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_211), .A2(n_265), .B1(n_399), .B2(n_424), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_212), .Y(n_808) );
INVx1_ASAP7_75t_L g487 ( .A(n_214), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_216), .A2(n_261), .B1(n_326), .B2(n_585), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_219), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_221), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_225), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_226), .A2(n_238), .B1(n_402), .B2(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_229), .B(n_786), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_231), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_232), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_236), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_237), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_240), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_242), .Y(n_452) );
INVx1_ASAP7_75t_L g784 ( .A(n_243), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_248), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_250), .B(n_547), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_251), .A2(n_588), .B1(n_621), .B2(n_622), .Y(n_587) );
INVx1_ASAP7_75t_L g621 ( .A(n_251), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_252), .Y(n_843) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_258), .B(n_417), .Y(n_599) );
INVx1_ASAP7_75t_L g496 ( .A(n_260), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_266), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_267), .Y(n_712) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_274), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_275), .A2(n_779), .B(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_626), .B1(n_774), .B2(n_775), .C(n_776), .Y(n_279) );
INVx1_ASAP7_75t_L g774 ( .A(n_280), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_442), .B2(n_625), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OA22x2_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_370), .B1(n_371), .B2(n_441), .Y(n_282) );
INVx1_ASAP7_75t_L g441 ( .A(n_283), .Y(n_441) );
INVx1_ASAP7_75t_L g369 ( .A(n_284), .Y(n_369) );
AND4x1_ASAP7_75t_L g284 ( .A(n_285), .B(n_318), .C(n_338), .D(n_357), .Y(n_284) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g485 ( .A(n_287), .Y(n_485) );
BUFx3_ASAP7_75t_L g615 ( .A(n_287), .Y(n_615) );
BUFx3_ASAP7_75t_L g757 ( .A(n_287), .Y(n_757) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g476 ( .A(n_288), .Y(n_476) );
BUFx2_ASAP7_75t_SL g578 ( .A(n_288), .Y(n_578) );
BUFx2_ASAP7_75t_SL g722 ( .A(n_288), .Y(n_722) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_298), .Y(n_288) );
AND2x6_ASAP7_75t_L g321 ( .A(n_289), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g327 ( .A(n_289), .B(n_311), .Y(n_327) );
AND2x6_ASAP7_75t_L g359 ( .A(n_289), .B(n_354), .Y(n_359) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
AND2x2_ASAP7_75t_L g306 ( .A(n_290), .B(n_296), .Y(n_306) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g312 ( .A(n_291), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_291), .B(n_296), .Y(n_317) );
AND2x2_ASAP7_75t_L g349 ( .A(n_291), .B(n_300), .Y(n_349) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
INVx1_ASAP7_75t_L g363 ( .A(n_296), .Y(n_363) );
AND2x4_ASAP7_75t_L g305 ( .A(n_298), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_298), .B(n_312), .Y(n_332) );
AND2x4_ASAP7_75t_L g336 ( .A(n_298), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g377 ( .A(n_298), .B(n_312), .Y(n_377) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_299), .B(n_302), .Y(n_311) );
OR2x2_ASAP7_75t_L g323 ( .A(n_299), .B(n_302), .Y(n_323) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g354 ( .A(n_300), .B(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
AND2x2_ASAP7_75t_L g362 ( .A(n_301), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g316 ( .A(n_302), .Y(n_316) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g852 ( .A(n_304), .Y(n_852) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_305), .Y(n_391) );
BUFx3_ASAP7_75t_L g465 ( .A(n_305), .Y(n_465) );
BUFx3_ASAP7_75t_L g617 ( .A(n_305), .Y(n_617) );
BUFx3_ASAP7_75t_L g747 ( .A(n_305), .Y(n_747) );
AND2x4_ASAP7_75t_L g341 ( .A(n_306), .B(n_322), .Y(n_341) );
AND2x6_ASAP7_75t_L g344 ( .A(n_306), .B(n_311), .Y(n_344) );
INVx1_ASAP7_75t_L g504 ( .A(n_306), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_306), .B(n_311), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_314), .B2(n_315), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_309), .A2(n_533), .B1(n_534), .B2(n_535), .Y(n_532) );
BUFx2_ASAP7_75t_R g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g382 ( .A(n_311), .B(n_312), .Y(n_382) );
INVx1_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
INVx6_ASAP7_75t_SL g384 ( .A(n_315), .Y(n_384) );
INVx1_ASAP7_75t_L g636 ( .A(n_315), .Y(n_636) );
INVx1_ASAP7_75t_SL g817 ( .A(n_315), .Y(n_817) );
OR2x6_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g400 ( .A(n_316), .Y(n_400) );
INVx1_ASAP7_75t_L g337 ( .A(n_317), .Y(n_337) );
INVx4_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g387 ( .A(n_320), .Y(n_387) );
INVx2_ASAP7_75t_SL g697 ( .A(n_320), .Y(n_697) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_320), .Y(n_763) );
INVx11_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx11_ASAP7_75t_L g429 ( .A(n_321), .Y(n_429) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g503 ( .A(n_323), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g436 ( .A(n_327), .Y(n_436) );
BUFx3_ASAP7_75t_L g463 ( .A(n_327), .Y(n_463) );
INVx6_ASAP7_75t_L g495 ( .A(n_327), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_333), .B2(n_334), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_330), .A2(n_542), .B1(n_543), .B2(n_544), .Y(n_541) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g642 ( .A(n_331), .Y(n_642) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_334), .A2(n_390), .B1(n_644), .B2(n_645), .Y(n_643) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_336), .Y(n_392) );
BUFx3_ASAP7_75t_L g437 ( .A(n_336), .Y(n_437) );
BUFx3_ASAP7_75t_L g478 ( .A(n_336), .Y(n_478) );
INVx1_ASAP7_75t_L g670 ( .A(n_336), .Y(n_670) );
BUFx3_ASAP7_75t_L g699 ( .A(n_336), .Y(n_699) );
BUFx2_ASAP7_75t_L g727 ( .A(n_336), .Y(n_727) );
BUFx3_ASAP7_75t_L g759 ( .A(n_336), .Y(n_759) );
AND2x2_ASAP7_75t_L g432 ( .A(n_337), .B(n_350), .Y(n_432) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g395 ( .A(n_340), .Y(n_395) );
INVx5_ASAP7_75t_L g547 ( .A(n_340), .Y(n_547) );
INVx4_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g396 ( .A(n_343), .Y(n_396) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
BUFx4f_ASAP7_75t_L g422 ( .A(n_344), .Y(n_422) );
BUFx2_ASAP7_75t_L g548 ( .A(n_344), .Y(n_548) );
BUFx2_ASAP7_75t_L g692 ( .A(n_344), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_351), .B2(n_352), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_347), .A2(n_550), .B1(n_551), .B2(n_552), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_347), .A2(n_352), .B1(n_717), .B2(n_718), .Y(n_716) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g603 ( .A(n_348), .Y(n_603) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_348), .Y(n_846) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x4_ASAP7_75t_L g361 ( .A(n_349), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g366 ( .A(n_349), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g399 ( .A(n_349), .B(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g552 ( .A(n_352), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_352), .A2(n_602), .B1(n_648), .B2(n_649), .Y(n_647) );
CKINVDCx16_ASAP7_75t_R g810 ( .A(n_352), .Y(n_810) );
OR2x6_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g402 ( .A(n_354), .B(n_356), .Y(n_402) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g565 ( .A(n_358), .Y(n_565) );
INVx2_ASAP7_75t_L g802 ( .A(n_358), .Y(n_802) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx4_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
INVx2_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
BUFx3_ASAP7_75t_L g451 ( .A(n_359), .Y(n_451) );
INVx2_ASAP7_75t_SL g683 ( .A(n_359), .Y(n_683) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_360), .Y(n_568) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g408 ( .A(n_361), .Y(n_408) );
BUFx4f_ASAP7_75t_SL g424 ( .A(n_361), .Y(n_424) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_361), .Y(n_516) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_361), .Y(n_555) );
INVx1_ASAP7_75t_L g367 ( .A(n_363), .Y(n_367) );
INVx1_ASAP7_75t_L g519 ( .A(n_364), .Y(n_519) );
BUFx4f_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g570 ( .A(n_365), .Y(n_570) );
BUFx12f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_410), .B1(n_439), .B2(n_440), .Y(n_371) );
INVx2_ASAP7_75t_SL g439 ( .A(n_372), .Y(n_439) );
XOR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_409), .Y(n_372) );
NOR4xp75_ASAP7_75t_L g373 ( .A(n_374), .B(n_385), .C(n_393), .D(n_403), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_375), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g859 ( .A(n_376), .Y(n_859) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g473 ( .A(n_377), .Y(n_473) );
BUFx3_ASAP7_75t_L g499 ( .A(n_377), .Y(n_499) );
BUFx3_ASAP7_75t_L g610 ( .A(n_377), .Y(n_610) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g490 ( .A(n_380), .Y(n_490) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx5_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g468 ( .A(n_381), .Y(n_468) );
BUFx3_ASAP7_75t_L g620 ( .A(n_381), .Y(n_620) );
INVx3_ASAP7_75t_L g765 ( .A(n_381), .Y(n_765) );
INVx8_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVxp67_ASAP7_75t_L g535 ( .A(n_383), .Y(n_535) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g581 ( .A(n_384), .Y(n_581) );
BUFx2_ASAP7_75t_L g704 ( .A(n_384), .Y(n_704) );
BUFx4f_ASAP7_75t_SL g854 ( .A(n_384), .Y(n_854) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx4_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_390), .A2(n_485), .B1(n_486), .B2(n_487), .C(n_488), .Y(n_484) );
OAI221xp5_ASAP7_75t_SL g812 ( .A1(n_390), .A2(n_813), .B1(n_814), .B2(n_815), .C(n_816), .Y(n_812) );
INVx4_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_397), .Y(n_393) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g458 ( .A(n_399), .Y(n_458) );
BUFx3_ASAP7_75t_L g665 ( .A(n_399), .Y(n_665) );
BUFx2_ASAP7_75t_L g769 ( .A(n_399), .Y(n_769) );
INVx1_ASAP7_75t_SL g687 ( .A(n_401), .Y(n_687) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_SL g418 ( .A(n_402), .Y(n_418) );
BUFx3_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
BUFx2_ASAP7_75t_SL g575 ( .A(n_402), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_406), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g554 ( .A(n_404), .Y(n_554) );
OAI221xp5_ASAP7_75t_SL g595 ( .A1(n_404), .A2(n_596), .B1(n_597), .B2(n_598), .C(n_599), .Y(n_595) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g512 ( .A1(n_405), .A2(n_513), .B1(n_517), .B2(n_518), .C1(n_519), .C2(n_520), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_405), .A2(n_651), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
XOR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_438), .Y(n_410) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_425), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_419), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_415), .B(n_416), .Y(n_413) );
BUFx2_ASAP7_75t_L g454 ( .A(n_417), .Y(n_454) );
BUFx3_ASAP7_75t_L g556 ( .A(n_417), .Y(n_556) );
INVx2_ASAP7_75t_L g652 ( .A(n_417), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .C(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g597 ( .A(n_424), .Y(n_597) );
INVx1_ASAP7_75t_L g800 ( .A(n_424), .Y(n_800) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_433), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_431), .Y(n_426) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_429), .A2(n_492), .B1(n_493), .B2(n_496), .C(n_497), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_429), .A2(n_538), .B1(n_539), .B2(n_540), .Y(n_537) );
INVx2_ASAP7_75t_SL g585 ( .A(n_429), .Y(n_585) );
INVx3_ASAP7_75t_L g634 ( .A(n_429), .Y(n_634) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_430), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g625 ( .A(n_442), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_523), .B2(n_624), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_480), .B1(n_481), .B2(n_522), .Y(n_444) );
INVx1_ASAP7_75t_L g522 ( .A(n_445), .Y(n_522) );
INVx1_ASAP7_75t_SL g479 ( .A(n_447), .Y(n_479) );
NAND3x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_461), .C(n_469), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_455), .Y(n_448) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_452), .B(n_453), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_450), .A2(n_714), .B(n_715), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g732 ( .A1(n_450), .A2(n_733), .B(n_734), .Y(n_732) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g511 ( .A(n_458), .Y(n_511) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
INVx1_ASAP7_75t_L g540 ( .A(n_463), .Y(n_540) );
INVx1_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_476), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_528) );
INVx3_ASAP7_75t_L g746 ( .A(n_476), .Y(n_746) );
INVx1_ASAP7_75t_L g544 ( .A(n_477), .Y(n_544) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g521 ( .A(n_483), .Y(n_521) );
OR4x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_491), .C(n_500), .D(n_512), .Y(n_483) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g612 ( .A(n_495), .Y(n_612) );
INVx3_ASAP7_75t_L g640 ( .A(n_495), .Y(n_640) );
INVx2_ASAP7_75t_L g702 ( .A(n_495), .Y(n_702) );
BUFx4f_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g822 ( .A(n_499), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_505), .B1(n_506), .B2(n_509), .C(n_510), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_501), .A2(n_798), .B1(n_838), .B2(n_839), .Y(n_837) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_503), .Y(n_592) );
BUFx3_ASAP7_75t_L g657 ( .A(n_503), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_506), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_506), .A2(n_657), .B1(n_711), .B2(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_SL g594 ( .A(n_507), .Y(n_594) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g798 ( .A(n_508), .Y(n_798) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI222xp33_ASAP7_75t_L g840 ( .A1(n_515), .A2(n_565), .B1(n_652), .B2(n_841), .C1(n_842), .C2(n_843), .Y(n_840) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g624 ( .A(n_523), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_559), .B2(n_560), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g558 ( .A(n_526), .Y(n_558) );
AND4x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .C(n_545), .D(n_553), .Y(n_526) );
NOR2xp33_ASAP7_75t_SL g527 ( .A(n_528), .B(n_532), .Y(n_527) );
NOR2xp33_ASAP7_75t_SL g536 ( .A(n_537), .B(n_541), .Y(n_536) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_547), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_552), .A2(n_601), .B1(n_602), .B2(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_586), .B1(n_587), .B2(n_623), .Y(n_560) );
INVx1_ASAP7_75t_L g623 ( .A(n_561), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_576), .C(n_582), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_566), .B(n_567), .Y(n_564) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .C(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g622 ( .A(n_588), .Y(n_622) );
AND2x2_ASAP7_75t_SL g588 ( .A(n_589), .B(n_605), .Y(n_588) );
NOR3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_595), .C(n_600), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_592), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_793) );
INVx3_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g807 ( .A(n_603), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_613), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .Y(n_613) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g775 ( .A(n_626), .Y(n_775) );
AOI22xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_752), .B1(n_772), .B2(n_773), .Y(n_626) );
INVx1_ASAP7_75t_L g772 ( .A(n_627), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_675), .B1(n_676), .B2(n_751), .Y(n_627) );
INVx1_ASAP7_75t_L g751 ( .A(n_628), .Y(n_751) );
XOR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_660), .Y(n_628) );
XOR2xp5_ASAP7_75t_SL g629 ( .A(n_630), .B(n_659), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_646), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_637), .C(n_643), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_641), .B2(n_642), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .C(n_655), .Y(n_646) );
OAI222xp33_ASAP7_75t_L g799 ( .A1(n_652), .A2(n_800), .B1(n_801), .B2(n_802), .C1(n_803), .C2(n_804), .Y(n_799) );
XOR2x2_ASAP7_75t_L g678 ( .A(n_660), .B(n_679), .Y(n_678) );
NAND4xp75_ASAP7_75t_L g661 ( .A(n_662), .B(n_666), .C(n_671), .D(n_674), .Y(n_661) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_705), .B2(n_750), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_681), .B(n_694), .Y(n_680) );
NOR2xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_688), .Y(n_681) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .B(n_685), .Y(n_682) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .C(n_693), .Y(n_688) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g750 ( .A(n_705), .Y(n_750) );
AO22x1_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_729), .B2(n_749), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
XOR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_728), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_719), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .C(n_716), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g813 ( .A(n_722), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx3_ASAP7_75t_SL g749 ( .A(n_729), .Y(n_749) );
XOR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_748), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_731), .B(n_739), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .C(n_738), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g773 ( .A(n_752), .Y(n_773) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
NAND4xp75_ASAP7_75t_SL g754 ( .A(n_755), .B(n_760), .C(n_766), .D(n_770), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
NOR2x1_ASAP7_75t_L g777 ( .A(n_778), .B(n_782), .Y(n_777) );
OR2x2_ASAP7_75t_SL g863 ( .A(n_778), .B(n_783), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_780), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_780), .B(n_829), .Y(n_832) );
CKINVDCx16_ASAP7_75t_R g829 ( .A(n_781), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
OAI322xp33_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_825), .A3(n_826), .B1(n_830), .B2(n_833), .C1(n_834), .C2(n_861), .Y(n_789) );
INVx1_ASAP7_75t_L g824 ( .A(n_791), .Y(n_824) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_811), .Y(n_791) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_799), .C(n_805), .Y(n_792) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_805) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g848 ( .A(n_810), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_818), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g860 ( .A(n_835), .Y(n_860) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_849), .Y(n_835) );
NOR3xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_840), .C(n_844), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_855), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_853), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g855 ( .A(n_856), .B(n_857), .Y(n_855) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
endmodule