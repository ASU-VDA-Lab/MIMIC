module fake_jpeg_31383_n_101 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_5),
.B1(n_7),
.B2(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_35),
.C(n_33),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_11),
.C(n_12),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_57),
.B1(n_28),
.B2(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_8),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_13),
.Y(n_73)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_16),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_67),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_19),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_84),
.B1(n_22),
.B2(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_21),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_62),
.C(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_83),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_86),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_81),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_87),
.Y(n_101)
);


endmodule