module fake_netlist_6_3071_n_74 (n_7, n_6, n_12, n_4, n_2, n_15, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_10, n_74);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_74;

wire n_41;
wire n_52;
wire n_16;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_18;
wire n_21;
wire n_24;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_72;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_73;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_17;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_19;
wire n_48;
wire n_47;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_1),
.B(n_7),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_20),
.C(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_25),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_25),
.Y(n_34)
);

OR2x6_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_29),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_20),
.A2(n_21),
.B1(n_28),
.B2(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_25),
.Y(n_37)
);

NOR2x1_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_36),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_27),
.B(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_33),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_35),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_48),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_47),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_53),
.B(n_52),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_56),
.B(n_54),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_59),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_64),
.B(n_54),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_62),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_54),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI21x1_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_67),
.B(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_71),
.B(n_17),
.Y(n_73)
);

AO21x2_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_21),
.B(n_17),
.Y(n_74)
);


endmodule