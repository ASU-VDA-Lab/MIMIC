module fake_jpeg_11047_n_103 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_50),
.Y(n_54)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_4),
.B2(n_7),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_72),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_32),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_70),
.C(n_74),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_1),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_14),
.C(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_1),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_2),
.B(n_3),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

NAND2x1_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_8),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.C(n_10),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_11),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_77),
.B1(n_76),
.B2(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_92),
.B1(n_93),
.B2(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_88),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_99),
.A3(n_92),
.B1(n_98),
.B2(n_18),
.C(n_20),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_102),
.Y(n_103)
);


endmodule