module fake_jpeg_707_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_39),
.C(n_30),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_38),
.B1(n_46),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_51),
.B1(n_12),
.B2(n_14),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_37),
.B(n_1),
.C(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_37),
.B1(n_44),
.B2(n_41),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_21),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_64),
.B(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_17),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_89),
.B(n_22),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_86),
.B1(n_26),
.B2(n_28),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_81),
.B1(n_88),
.B2(n_83),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_100),
.C(n_94),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_91),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_97),
.B1(n_93),
.B2(n_92),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_96),
.B(n_95),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_106),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_8),
.Y(n_108)
);


endmodule