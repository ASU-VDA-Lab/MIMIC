module fake_jpeg_25509_n_144 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp33_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_10),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_21),
.Y(n_28)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_20),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_22),
.A2(n_18),
.B1(n_11),
.B2(n_14),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_37),
.B1(n_22),
.B2(n_27),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_22),
.A2(n_18),
.B1(n_11),
.B2(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_41),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_47),
.B1(n_16),
.B2(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_45),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_23),
.B(n_24),
.C(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_18),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_47),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_41),
.B1(n_42),
.B2(n_38),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_50),
.B(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_47),
.B1(n_30),
.B2(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_44),
.B1(n_33),
.B2(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_60),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_81),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_64),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_50),
.C(n_25),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_50),
.B(n_11),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_63),
.B1(n_71),
.B2(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_89),
.B1(n_93),
.B2(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_65),
.B1(n_16),
.B2(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_12),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_106),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_21),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_84),
.B1(n_93),
.B2(n_12),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_104),
.B1(n_19),
.B2(n_3),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_1),
.B(n_5),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_25),
.C(n_20),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_20),
.C(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_21),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_98),
.B(n_7),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_6),
.Y(n_128)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_107),
.B(n_115),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_128),
.A3(n_129),
.B1(n_121),
.B2(n_123),
.C(n_118),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_115),
.A3(n_7),
.B1(n_8),
.B2(n_6),
.C1(n_19),
.C2(n_25),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_120),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_133),
.B(n_19),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_117),
.B(n_8),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_8),
.B1(n_20),
.B2(n_19),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

AOI21x1_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_19),
.B(n_26),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_21),
.C(n_26),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_139),
.C(n_137),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_143),
.Y(n_144)
);


endmodule