module fake_jpeg_8759_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_22),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_17),
.B(n_9),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_27)
);

A2O1A1O1Ixp25_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_28),
.B(n_10),
.C(n_11),
.D(n_7),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_22),
.C(n_8),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_7),
.C(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_13),
.B(n_2),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_3),
.B(n_6),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_30),
.C(n_15),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_37),
.B(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_1),
.B1(n_16),
.B2(n_38),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_1),
.Y(n_41)
);


endmodule