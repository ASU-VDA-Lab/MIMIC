module fake_jpeg_13824_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_57),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_46),
.B(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_21),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_74),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_49),
.Y(n_135)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_6),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_66),
.Y(n_111)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_72),
.Y(n_113)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_75),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_77),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_8),
.B(n_13),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_83),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_26),
.B1(n_40),
.B2(n_17),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_42),
.B1(n_40),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_92),
.A2(n_96),
.B1(n_97),
.B2(n_132),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_26),
.B1(n_42),
.B2(n_24),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_118),
.B1(n_128),
.B2(n_87),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_43),
.A2(n_40),
.B1(n_24),
.B2(n_32),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_38),
.B1(n_23),
.B2(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_34),
.B1(n_35),
.B2(n_32),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_101),
.A2(n_116),
.B1(n_121),
.B2(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_123),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_38),
.B1(n_25),
.B2(n_23),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_37),
.B1(n_20),
.B2(n_3),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_69),
.A2(n_37),
.B1(n_20),
.B2(n_8),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_59),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_56),
.A2(n_74),
.B1(n_68),
.B2(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_0),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_2),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_2),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_57),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_136),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_66),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_140),
.Y(n_207)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_144),
.B(n_164),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_92),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_112),
.B1(n_103),
.B2(n_108),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_10),
.C(n_12),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_3),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_4),
.B(n_5),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_121),
.B1(n_124),
.B2(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_150),
.A2(n_174),
.B1(n_162),
.B2(n_173),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_151),
.A2(n_176),
.B1(n_158),
.B2(n_177),
.Y(n_213)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_133),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_159),
.C(n_164),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_163),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_157),
.A2(n_147),
.B1(n_172),
.B2(n_170),
.Y(n_209)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_88),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_111),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_167),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_161),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_87),
.A2(n_93),
.B1(n_129),
.B2(n_125),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_162),
.A2(n_170),
.B(n_140),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_94),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_88),
.B(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

BUFx6f_ASAP7_75t_SL g166 ( 
.A(n_120),
.Y(n_166)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_127),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_119),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_171),
.Y(n_187)
);

OR2x4_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_132),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_120),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_112),
.B1(n_108),
.B2(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_86),
.B(n_102),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_93),
.A2(n_114),
.B1(n_86),
.B2(n_110),
.Y(n_176)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_91),
.B(n_106),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_102),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_178),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_148),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_181),
.A2(n_211),
.B(n_204),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_99),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_208),
.B1(n_213),
.B2(n_157),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_103),
.Y(n_192)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_102),
.B1(n_106),
.B2(n_153),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_206),
.B1(n_209),
.B2(n_186),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_106),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_164),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_159),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_146),
.B1(n_145),
.B2(n_172),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_155),
.B(n_140),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_215),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_218),
.B(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_155),
.C(n_159),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_231),
.C(n_198),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_137),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_139),
.B(n_168),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_160),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_141),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_142),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_165),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_152),
.B1(n_161),
.B2(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_182),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_207),
.B1(n_191),
.B2(n_202),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_206),
.B1(n_181),
.B2(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_189),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_181),
.A2(n_195),
.B1(n_189),
.B2(n_199),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_240),
.B1(n_205),
.B2(n_199),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_186),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_200),
.B1(n_180),
.B2(n_212),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_205),
.B1(n_183),
.B2(n_190),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_186),
.B(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_198),
.B(n_180),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_263),
.B(n_253),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_242),
.C(n_228),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_200),
.B1(n_212),
.B2(n_180),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_256),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_217),
.B1(n_221),
.B2(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_217),
.A2(n_218),
.B1(n_215),
.B2(n_237),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_240),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_238),
.B(n_219),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_223),
.B1(n_236),
.B2(n_226),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_223),
.B(n_264),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_266),
.A2(n_278),
.B(n_246),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_220),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_269),
.C(n_270),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_260),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_SL g292 ( 
.A(n_268),
.B(n_275),
.C(n_277),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_223),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_224),
.C(n_230),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_246),
.C(n_254),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_281),
.B1(n_282),
.B2(n_244),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_227),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_251),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_229),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_263),
.B(n_262),
.Y(n_284)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_256),
.B1(n_248),
.B2(n_252),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_289),
.B1(n_281),
.B2(n_279),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_243),
.B1(n_255),
.B2(n_253),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_295),
.B1(n_283),
.B2(n_272),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_267),
.B(n_258),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_244),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_297),
.C(n_283),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_280),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_268),
.A2(n_281),
.B1(n_276),
.B2(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

AO221x1_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_278),
.B1(n_275),
.B2(n_266),
.C(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_288),
.C(n_291),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_295),
.B1(n_277),
.B2(n_273),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_309),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_282),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_308),
.Y(n_317)
);

BUFx12_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_309),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_288),
.C(n_290),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_300),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_307),
.B(n_300),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_319),
.B(n_318),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_306),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_317),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_306),
.Y(n_324)
);

BUFx4f_ASAP7_75t_SL g325 ( 
.A(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_317),
.B(n_309),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_315),
.B1(n_320),
.B2(n_325),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_330),
.B(n_325),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_323),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_330),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_229),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_229),
.Y(n_339)
);


endmodule