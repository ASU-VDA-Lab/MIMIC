module fake_jpeg_31282_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_46),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_49),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_50),
.B(n_59),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_51),
.Y(n_113)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g124 ( 
.A(n_54),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_33),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_14),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_13),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_16),
.B(n_13),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_86),
.Y(n_123)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_22),
.B1(n_38),
.B2(n_23),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_90),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_61),
.B1(n_59),
.B2(n_50),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_96),
.A2(n_102),
.B1(n_105),
.B2(n_134),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_16),
.B1(n_42),
.B2(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_97),
.A2(n_99),
.B1(n_106),
.B2(n_114),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_27),
.B1(n_25),
.B2(n_16),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_98),
.A2(n_100),
.B1(n_103),
.B2(n_117),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_42),
.B1(n_19),
.B2(n_41),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_27),
.B1(n_42),
.B2(n_23),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_86),
.B1(n_87),
.B2(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_42),
.B1(n_23),
.B2(n_38),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_48),
.A2(n_36),
.B1(n_29),
.B2(n_30),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_29),
.B1(n_36),
.B2(n_30),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_33),
.B1(n_37),
.B2(n_23),
.Y(n_110)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_110),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_33),
.B1(n_23),
.B2(n_43),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_43),
.B1(n_31),
.B2(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_115),
.A2(n_125),
.B1(n_128),
.B2(n_124),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_44),
.A2(n_22),
.B1(n_21),
.B2(n_11),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_43),
.B1(n_31),
.B2(n_10),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_24),
.B1(n_31),
.B2(n_3),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_52),
.B(n_74),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_60),
.B1(n_53),
.B2(n_71),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_84),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_142),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_67),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_141),
.B(n_145),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_84),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_144),
.A2(n_169),
.B1(n_177),
.B2(n_139),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g221 ( 
.A(n_146),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_147),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_58),
.Y(n_148)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_94),
.B(n_51),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_153),
.Y(n_190)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_152),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_159),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_187),
.B1(n_189),
.B2(n_93),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_81),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_51),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_161),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_49),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_162),
.A2(n_119),
.B1(n_138),
.B2(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_164),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_118),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_166),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_7),
.Y(n_166)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_7),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_131),
.Y(n_202)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_107),
.A2(n_8),
.B(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_188),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_8),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_176),
.C(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_109),
.C(n_107),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_89),
.A2(n_133),
.B1(n_105),
.B2(n_139),
.Y(n_177)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_180),
.Y(n_215)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_110),
.C(n_102),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_110),
.A2(n_89),
.B1(n_133),
.B2(n_104),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_155),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_110),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_195),
.B(n_196),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_93),
.B(n_111),
.C(n_120),
.Y(n_196)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_179),
.B1(n_165),
.B2(n_157),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_213),
.B1(n_220),
.B2(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_132),
.Y(n_205)
);

CKINVDCx12_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_206),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_132),
.B1(n_129),
.B2(n_101),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_129),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_227),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_119),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_223),
.B(n_224),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_140),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_169),
.A2(n_189),
.B1(n_179),
.B2(n_158),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_178),
.B(n_142),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_233),
.A2(n_226),
.B(n_232),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_191),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_241),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_140),
.B1(n_142),
.B2(n_169),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_236),
.A2(n_238),
.B1(n_240),
.B2(n_244),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_156),
.B1(n_184),
.B2(n_164),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_143),
.B1(n_151),
.B2(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_230),
.B1(n_192),
.B2(n_202),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_247),
.A2(n_256),
.B1(n_248),
.B2(n_238),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_175),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_181),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_255),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_172),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_192),
.A2(n_174),
.B1(n_185),
.B2(n_152),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_204),
.A2(n_146),
.B1(n_186),
.B2(n_155),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_261),
.B1(n_265),
.B2(n_219),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_149),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_167),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_192),
.A2(n_213),
.B1(n_210),
.B2(n_196),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_229),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_199),
.B(n_217),
.C(n_225),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_267),
.C(n_235),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_212),
.B(n_193),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_224),
.A2(n_222),
.B1(n_198),
.B2(n_228),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_209),
.B(n_197),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_221),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_272),
.A2(n_276),
.B(n_277),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_278),
.B(n_284),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_209),
.B(n_193),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_233),
.A2(n_212),
.B(n_209),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_221),
.B(n_197),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_249),
.B(n_228),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_286),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_269),
.Y(n_281)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_282),
.A2(n_297),
.B1(n_272),
.B2(n_291),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_197),
.B(n_219),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_263),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_236),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_247),
.B1(n_244),
.B2(n_257),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_255),
.B(n_262),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g320 ( 
.A1(n_290),
.A2(n_293),
.B(n_256),
.C(n_254),
.D(n_265),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_251),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_294),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_234),
.B(n_259),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_237),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_300),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_252),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_234),
.B(n_243),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_267),
.Y(n_318)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_239),
.B1(n_242),
.B2(n_245),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_282),
.B1(n_299),
.B2(n_289),
.Y(n_333)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

NAND4xp25_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_266),
.C(n_268),
.D(n_260),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_309),
.B(n_312),
.Y(n_330)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_285),
.B(n_246),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_300),
.B1(n_298),
.B2(n_296),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_315),
.A2(n_325),
.B1(n_288),
.B2(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_273),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_295),
.Y(n_322)
);

BUFx12f_ASAP7_75t_SL g323 ( 
.A(n_276),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_324),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_260),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_299),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_286),
.C(n_292),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_339),
.B1(n_320),
.B2(n_303),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_333),
.B(n_316),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_280),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_307),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_287),
.B1(n_288),
.B2(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_270),
.Y(n_342)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_270),
.C(n_290),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_346),
.C(n_338),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_278),
.C(n_284),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_274),
.Y(n_348)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_337),
.A2(n_323),
.B(n_314),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_356),
.B(n_335),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_354),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_360),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_348),
.A2(n_314),
.B(n_277),
.Y(n_356)
);

BUFx12_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_365),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_321),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_362),
.A2(n_367),
.B1(n_334),
.B2(n_346),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_334),
.A2(n_303),
.B1(n_316),
.B2(n_302),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_364),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_306),
.C(n_318),
.Y(n_365)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_366),
.A2(n_344),
.B1(n_349),
.B2(n_350),
.Y(n_382)
);

AOI221xp5_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_303),
.B1(n_302),
.B2(n_307),
.C(n_305),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_371),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_354),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_361),
.B(n_345),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_374),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_332),
.C(n_335),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_375),
.A2(n_380),
.B1(n_362),
.B2(n_367),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_377),
.A2(n_357),
.B(n_366),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_336),
.C(n_343),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_382),
.B(n_383),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_336),
.B1(n_343),
.B2(n_344),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_361),
.B(n_350),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_372),
.A2(n_358),
.B(n_355),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_385),
.B(n_371),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_377),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_394),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_389),
.B1(n_369),
.B2(n_380),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_381),
.A2(n_353),
.B(n_360),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_391),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_375),
.A2(n_368),
.B1(n_359),
.B2(n_363),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g391 ( 
.A1(n_381),
.A2(n_356),
.B(n_359),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_379),
.A2(n_363),
.B1(n_349),
.B2(n_308),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_392),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_400),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_393),
.B(n_370),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_401),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_390),
.A2(n_374),
.B(n_378),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_SL g406 ( 
.A1(n_398),
.A2(n_386),
.B(n_392),
.C(n_387),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_394),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_376),
.C(n_384),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_406),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_376),
.C(n_357),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_407),
.A2(n_403),
.B(n_402),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_399),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_409),
.B(n_404),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_410),
.A2(n_397),
.B(n_357),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_411),
.B(n_412),
.C(n_408),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_413),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_366),
.Y(n_415)
);


endmodule