module fake_jpeg_14793_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_2),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_34),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_3),
.C(n_4),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_25),
.C(n_19),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_3),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_62),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_67),
.Y(n_92)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_4),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_23),
.Y(n_79)
);

OR2x4_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_24),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_81),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_93),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_84),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_24),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_102),
.B1(n_103),
.B2(n_28),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_68),
.B1(n_63),
.B2(n_66),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_26),
.B1(n_28),
.B2(n_6),
.Y(n_122)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_33),
.B1(n_25),
.B2(n_19),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_33),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_60),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_55),
.B(n_29),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_128),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_122),
.B1(n_75),
.B2(n_72),
.Y(n_158)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_138),
.Y(n_179)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_131),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_15),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_79),
.B1(n_80),
.B2(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_136),
.B1(n_149),
.B2(n_116),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_104),
.B(n_98),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_137),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_78),
.B(n_5),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_108),
.C(n_91),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_86),
.A2(n_89),
.B(n_99),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_75),
.B(n_89),
.C(n_98),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_11),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_77),
.B(n_13),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_109),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_13),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_93),
.B(n_13),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_108),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_14),
.B1(n_82),
.B2(n_105),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_169),
.B(n_179),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_159),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_168),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_119),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_87),
.C(n_104),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_123),
.C(n_139),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_113),
.B1(n_144),
.B2(n_137),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_177),
.B1(n_134),
.B2(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_149),
.B1(n_122),
.B2(n_142),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_129),
.Y(n_191)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_99),
.B1(n_85),
.B2(n_74),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_115),
.B(n_135),
.C(n_118),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_189),
.B1(n_195),
.B2(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_150),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_203),
.B(n_169),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_124),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_201),
.C(n_164),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_157),
.A2(n_124),
.B1(n_136),
.B2(n_147),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_157),
.A2(n_140),
.B1(n_134),
.B2(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_123),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_163),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_139),
.B(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_178),
.B(n_153),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_219),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_209),
.C(n_222),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_153),
.B1(n_198),
.B2(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_211),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_201),
.C(n_196),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_167),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_221),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_160),
.C(n_152),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_173),
.B(n_160),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_203),
.A2(n_167),
.B(n_171),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_185),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_220),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_176),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_193),
.B1(n_198),
.B2(n_184),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_232),
.B1(n_218),
.B2(n_214),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_200),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_202),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.C(n_156),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_189),
.B1(n_183),
.B2(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_210),
.C(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_212),
.B1(n_213),
.B2(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_212),
.B1(n_213),
.B2(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_241),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_206),
.B(n_217),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_242),
.B(n_243),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_216),
.B(n_173),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_210),
.A3(n_199),
.B1(n_195),
.B2(n_156),
.C1(n_177),
.C2(n_162),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_247),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_162),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_223),
.C(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_188),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_253),
.C(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_223),
.C(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_228),
.B1(n_224),
.B2(n_235),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_172),
.B1(n_182),
.B2(n_175),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_260),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_240),
.B(n_242),
.C(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_262),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_174),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_249),
.Y(n_265)
);

OAI221xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_255),
.B1(n_239),
.B2(n_252),
.C(n_225),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_259),
.C(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_250),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

OAI321xp33_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.A3(n_269),
.B1(n_262),
.B2(n_259),
.C(n_166),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_269),
.B(n_263),
.CI(n_253),
.CON(n_270),
.SN(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);


endmodule