module fake_jpeg_26702_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_24),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_29),
.B1(n_15),
.B2(n_28),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_19),
.B1(n_24),
.B2(n_30),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_28),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_33),
.C(n_36),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_21),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_32),
.A2(n_25),
.B1(n_20),
.B2(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_27),
.B1(n_19),
.B2(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_0),
.Y(n_77)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_66),
.B(n_67),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_20),
.B1(n_40),
.B2(n_24),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_78),
.B1(n_58),
.B2(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_27),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_43),
.B1(n_51),
.B2(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_76),
.A2(n_52),
.B1(n_43),
.B2(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_86),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_61),
.B(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_90),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_54),
.C(n_48),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_67),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_43),
.B1(n_50),
.B2(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_67),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_56),
.B1(n_50),
.B2(n_35),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_99),
.B1(n_74),
.B2(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_84),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_45),
.B1(n_5),
.B2(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_112),
.Y(n_130)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_102),
.Y(n_133)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_66),
.A3(n_67),
.B1(n_68),
.B2(n_78),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_118),
.B(n_8),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_89),
.C(n_45),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_110),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_108),
.B(n_89),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_65),
.B(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_6),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_90),
.B(n_85),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_79),
.B1(n_93),
.B2(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_92),
.B1(n_85),
.B2(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_92),
.B1(n_106),
.B2(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_83),
.B(n_88),
.C(n_81),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_103),
.B(n_111),
.C(n_106),
.D(n_101),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_104),
.C(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_127),
.C(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_132),
.B(n_126),
.C(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_144),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_126),
.B1(n_129),
.B2(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_150),
.B1(n_140),
.B2(n_149),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_138),
.C(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_9),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_131),
.B(n_124),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_132),
.C(n_119),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_143),
.C(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_172),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_137),
.C(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_120),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_163),
.B(n_162),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_12),
.Y(n_188)
);

NAND2x1p5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_11),
.Y(n_186)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_165),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_155),
.C(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_101),
.C(n_13),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_12),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_158),
.B1(n_170),
.B2(n_154),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_179),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_187),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_177),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_180),
.C(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_188),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_180),
.C(n_189),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_190),
.B1(n_192),
.B2(n_13),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_192),
.B(n_14),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_198),
.B(n_14),
.Y(n_201)
);


endmodule