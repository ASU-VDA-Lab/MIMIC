module fake_netlist_6_1745_n_2153 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2153);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2153;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVxp67_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_71),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_62),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_54),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_65),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_40),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_173),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_39),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_36),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_2),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_67),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_21),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_100),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_81),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_4),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_160),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_95),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_132),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_168),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_117),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_182),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_188),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_151),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_69),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_206),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_81),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_85),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_215),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_57),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_43),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_109),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_193),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_153),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_147),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_0),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_16),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_126),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_28),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_122),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_70),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_61),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_75),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_23),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_13),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_194),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_178),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_54),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_210),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_78),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_74),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_158),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_164),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_39),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_148),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_101),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_55),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_185),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_127),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_80),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_128),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_141),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_121),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_5),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_91),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_130),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_74),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_169),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_115),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_183),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_90),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_9),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_139),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_179),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_16),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_198),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_162),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_19),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_114),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_55),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_56),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_83),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_61),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_25),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_82),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_192),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_42),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_197),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_105),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_143),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_149),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_78),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_167),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_9),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_125),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_29),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_118),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_152),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_142),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_43),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_208),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_200),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_31),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_41),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_6),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_11),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_213),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_190),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_52),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_120),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_13),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_205),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_72),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_176),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_7),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_96),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_79),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_29),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_146),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_36),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_79),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_201),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_88),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_50),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_89),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_112),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_123),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_116),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_150),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_174),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_19),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_113),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_196),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_97),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_92),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_106),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_203),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_163),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_4),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_68),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_124),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_191),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_70),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_30),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_44),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_186),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_57),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_145),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_6),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_87),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_18),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_214),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_71),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_131),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_217),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_45),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_28),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_166),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_171),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_195),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_58),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_33),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_98),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_52),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_59),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_82),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_133),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_189),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_49),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_180),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_144),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_59),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_212),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_202),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_41),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_165),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_119),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_40),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_108),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_50),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_156),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_129),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_49),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_170),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_135),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_24),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_47),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_199),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_137),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_44),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_216),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_140),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_155),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_8),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_72),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_42),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_83),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_211),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_209),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_231),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_222),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_228),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_433),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_433),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_289),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_300),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_300),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_233),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_237),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_324),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_240),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_324),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_284),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_238),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_238),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_238),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_293),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_298),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_293),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_293),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_404),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_437),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_404),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_234),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_286),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_234),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_236),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_243),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_236),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_244),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_254),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_254),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_245),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_272),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_288),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_373),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_272),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_399),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_396),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_273),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_273),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_247),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_408),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_279),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_408),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_399),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_288),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_302),
.Y(n_492)
);

BUFx2_ASAP7_75t_SL g493 ( 
.A(n_311),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_249),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_231),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_286),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_241),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_290),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_250),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_375),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_302),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_252),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_255),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_279),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_283),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_304),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_283),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_258),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_259),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_318),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_318),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_262),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_263),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_409),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_321),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_288),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_321),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_309),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_264),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_265),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_220),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_313),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_331),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_331),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_241),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_266),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_333),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_333),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_313),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_337),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_274),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_337),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_281),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_282),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_223),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_340),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_340),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_341),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_221),
.Y(n_539)
);

INVxp33_ASAP7_75t_SL g540 ( 
.A(n_224),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_287),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_341),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_342),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_291),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_313),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_342),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_242),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_242),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_292),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_350),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_294),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_297),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_350),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_358),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_358),
.Y(n_555)
);

INVx4_ASAP7_75t_R g556 ( 
.A(n_345),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_369),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_369),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_440),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_441),
.B(n_345),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_539),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_470),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_539),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_449),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_447),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_471),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_450),
.B(n_345),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_491),
.B(n_516),
.Y(n_573)
);

INVx6_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_521),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_529),
.B(n_347),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_452),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_479),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_472),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_474),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_454),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_461),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_444),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_473),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_477),
.B(n_347),
.Y(n_590)
);

BUFx8_ASAP7_75t_L g591 ( 
.A(n_522),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_446),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_475),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_439),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_495),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_476),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_545),
.B(n_493),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_497),
.B(n_347),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_525),
.B(n_311),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_457),
.B(n_377),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_493),
.B(n_372),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_518),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_535),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_540),
.B(n_482),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_480),
.B(n_227),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_469),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_548),
.B(n_372),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_458),
.B(n_380),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_458),
.B(n_380),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_459),
.B(n_420),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_478),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_448),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_448),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_451),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_483),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_459),
.B(n_420),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_481),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_451),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_506),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_453),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_481),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_453),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_460),
.B(n_462),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_498),
.B(n_225),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_486),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_460),
.B(n_438),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_500),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_455),
.A2(n_248),
.B(n_246),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_462),
.A2(n_299),
.B(n_221),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_463),
.B(n_303),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_484),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_494),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_499),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_456),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_502),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_490),
.B(n_366),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_484),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_456),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_463),
.B(n_377),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_485),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_485),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_503),
.B(n_299),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_488),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_464),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_488),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_563),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_606),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_563),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_562),
.B(n_508),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_606),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_606),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_572),
.B(n_509),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_565),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_573),
.B(n_464),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_565),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_512),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_576),
.B(n_221),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_565),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_652),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_652),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_652),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_600),
.A2(n_501),
.B1(n_492),
.B2(n_466),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_613),
.B(n_487),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_577),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_650),
.B(n_513),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_631),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_626),
.B(n_519),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_629),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_574),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_594),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_573),
.B(n_600),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_574),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_526),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_631),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_613),
.B(n_445),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_629),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_629),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_577),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_629),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_576),
.B(n_531),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_631),
.A2(n_496),
.B1(n_378),
.B2(n_385),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_604),
.B(n_465),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_626),
.B(n_534),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_615),
.A2(n_378),
.B1(n_385),
.B2(n_382),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_577),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_577),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_612),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_644),
.B(n_541),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_629),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_570),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_574),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_630),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_630),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_617),
.A2(n_415),
.B(n_330),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_574),
.B(n_330),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_630),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_585),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_594),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_544),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_609),
.B(n_552),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_630),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_594),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_594),
.Y(n_715)
);

AND3x2_ASAP7_75t_L g716 ( 
.A(n_622),
.B(n_280),
.C(n_253),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_581),
.B(n_393),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

NOR2x1p5_ASAP7_75t_L g719 ( 
.A(n_559),
.B(n_317),
.Y(n_719)
);

CKINVDCx14_ASAP7_75t_R g720 ( 
.A(n_587),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_603),
.B(n_330),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_632),
.B(n_489),
.C(n_608),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_594),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_604),
.B(n_465),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_630),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_SL g726 ( 
.A(n_607),
.B(n_520),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_642),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_601),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_594),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_581),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_626),
.A2(n_549),
.B1(n_551),
.B2(n_533),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_642),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_642),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_642),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_595),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_581),
.B(n_415),
.Y(n_736)
);

BUFx10_ASAP7_75t_L g737 ( 
.A(n_566),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_595),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_581),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_578),
.B(n_467),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_595),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_595),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_582),
.B(n_467),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_626),
.B(n_306),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_642),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_595),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_601),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_595),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_601),
.B(n_407),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_610),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_601),
.B(n_307),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_615),
.A2(n_387),
.B1(n_390),
.B2(n_382),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_610),
.Y(n_753)
);

BUFx10_ASAP7_75t_L g754 ( 
.A(n_584),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_642),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_615),
.A2(n_390),
.B1(n_392),
.B2(n_387),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_615),
.A2(n_403),
.B1(n_411),
.B2(n_392),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_567),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_635),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_610),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_626),
.B(n_308),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_610),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_626),
.B(n_310),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_567),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_617),
.A2(n_415),
.B(n_248),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_602),
.A2(n_268),
.B1(n_277),
.B2(n_235),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_607),
.A2(n_359),
.B1(n_435),
.B2(n_354),
.Y(n_767)
);

INVx11_ASAP7_75t_L g768 ( 
.A(n_591),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_567),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_568),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_601),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_314),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_626),
.B(n_323),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_568),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_591),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_647),
.B(n_504),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_610),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_634),
.B(n_325),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_610),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_568),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_579),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_560),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_579),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_579),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_560),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_561),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_633),
.B(n_326),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_616),
.A2(n_623),
.B1(n_602),
.B2(n_614),
.Y(n_788)
);

INVx8_ASAP7_75t_L g789 ( 
.A(n_640),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_638),
.B(n_256),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_636),
.B(n_524),
.C(n_251),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_641),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_636),
.B(n_251),
.C(n_246),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_638),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_643),
.B(n_256),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_647),
.B(n_504),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_602),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_602),
.B(n_514),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_612),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_616),
.B(n_219),
.Y(n_800)
);

BUFx6f_ASAP7_75t_SL g801 ( 
.A(n_603),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_636),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_256),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_583),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_583),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_616),
.B(n_269),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_616),
.B(n_505),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_623),
.A2(n_403),
.B1(n_434),
.B2(n_411),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_637),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_561),
.A2(n_320),
.B1(n_436),
.B2(n_362),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_583),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_564),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_564),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_569),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_SL g815 ( 
.A1(n_637),
.A2(n_422),
.B(n_419),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_666),
.B(n_721),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_675),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_797),
.B(n_623),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_654),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_794),
.B(n_603),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_681),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_672),
.B(n_608),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_654),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_680),
.B(n_591),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_718),
.B(n_256),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_701),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_797),
.A2(n_614),
.B1(n_623),
.B2(n_351),
.Y(n_828)
);

OAI22x1_ASAP7_75t_R g829 ( 
.A1(n_709),
.A2(n_400),
.B1(n_322),
.B2(n_759),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_656),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_728),
.A2(n_588),
.B(n_614),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_657),
.B(n_614),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_693),
.B(n_569),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_718),
.B(n_256),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_691),
.A2(n_334),
.B1(n_338),
.B2(n_327),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_656),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_666),
.A2(n_271),
.B1(n_295),
.B2(n_269),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_709),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_660),
.B(n_598),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_661),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_665),
.B(n_598),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_739),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_661),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_655),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_683),
.B(n_591),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_662),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_674),
.B(n_598),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_666),
.A2(n_295),
.B1(n_316),
.B2(n_271),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_658),
.B(n_598),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_693),
.B(n_571),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_659),
.B(n_619),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_718),
.B(n_256),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_726),
.A2(n_349),
.B1(n_353),
.B2(n_339),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_668),
.B(n_619),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_668),
.B(n_619),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_673),
.B(n_305),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_669),
.B(n_620),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_663),
.B(n_571),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_669),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_229),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_673),
.B(n_305),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_670),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_670),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_673),
.B(n_305),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_788),
.B(n_620),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_759),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_772),
.B(n_620),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_678),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_SL g869 ( 
.A(n_801),
.B(n_328),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_778),
.B(n_620),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_663),
.B(n_627),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_662),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_720),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_685),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_782),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_689),
.B(n_627),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_782),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_785),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_666),
.A2(n_365),
.B1(n_371),
.B2(n_361),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_689),
.B(n_627),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_701),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_785),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_807),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_689),
.B(n_305),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_666),
.A2(n_368),
.B1(n_332),
.B2(n_335),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_786),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_740),
.B(n_230),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_786),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_SL g889 ( 
.A(n_809),
.B(n_775),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_666),
.A2(n_423),
.B1(n_413),
.B2(n_416),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_812),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_815),
.A2(n_434),
.B(n_422),
.C(n_419),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_807),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_696),
.Y(n_894)
);

BUFx4f_ASAP7_75t_L g895 ( 
.A(n_789),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_664),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_791),
.A2(n_406),
.B1(n_335),
.B2(n_336),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_743),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_696),
.B(n_627),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_696),
.B(n_336),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_812),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_789),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_697),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_697),
.B(n_344),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_697),
.B(n_305),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_813),
.B(n_814),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_813),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_664),
.Y(n_908)
);

AND2x6_ASAP7_75t_L g909 ( 
.A(n_809),
.B(n_344),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_667),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_802),
.B(n_305),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_739),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_791),
.A2(n_356),
.B1(n_360),
.B2(n_364),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_814),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_776),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_711),
.B(n_232),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_776),
.B(n_356),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_796),
.B(n_360),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_796),
.B(n_364),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_724),
.B(n_367),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_667),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_747),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_758),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_724),
.B(n_367),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_802),
.B(n_363),
.Y(n_926)
);

INVx5_ASAP7_75t_L g927 ( 
.A(n_809),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_800),
.B(n_368),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_764),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_769),
.Y(n_930)
);

INVxp33_ASAP7_75t_L g931 ( 
.A(n_672),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_712),
.B(n_239),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_SL g933 ( 
.A1(n_789),
.A2(n_226),
.B1(n_376),
.B2(n_370),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_802),
.B(n_370),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_769),
.Y(n_935)
);

INVx4_ASAP7_75t_L g936 ( 
.A(n_747),
.Y(n_936)
);

CKINVDCx11_ASAP7_75t_R g937 ( 
.A(n_737),
.Y(n_937)
);

BUFx8_ASAP7_75t_L g938 ( 
.A(n_775),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_671),
.B(n_257),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_798),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_802),
.B(n_702),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_SL g942 ( 
.A(n_766),
.B(n_261),
.C(n_260),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_702),
.B(n_374),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_770),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_809),
.B(n_363),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_770),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_774),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_730),
.B(n_374),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_787),
.B(n_267),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_730),
.B(n_376),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_810),
.B(n_270),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_774),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_809),
.B(n_363),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_780),
.Y(n_954)
);

AND2x4_ASAP7_75t_SL g955 ( 
.A(n_737),
.B(n_226),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_806),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_771),
.B(n_386),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_719),
.A2(n_379),
.B1(n_384),
.B2(n_432),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_771),
.B(n_386),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_717),
.B(n_749),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_793),
.B(n_363),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_780),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_678),
.B(n_406),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_781),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_781),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_678),
.B(n_424),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_721),
.A2(n_424),
.B1(n_428),
.B2(n_363),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_793),
.B(n_363),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_815),
.B(n_388),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_783),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_806),
.B(n_676),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_783),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_784),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_784),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_789),
.B(n_428),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_804),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_682),
.B(n_580),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_737),
.B(n_580),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_682),
.B(n_586),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_716),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_804),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_956),
.B(n_806),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_927),
.Y(n_983)
);

AO22x1_ASAP7_75t_L g984 ( 
.A1(n_939),
.A2(n_722),
.B1(n_731),
.B2(n_698),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_897),
.A2(n_721),
.B1(n_752),
.B2(n_695),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_860),
.A2(n_719),
.B1(n_801),
.B2(n_721),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_827),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_832),
.B(n_806),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_860),
.B(n_806),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_916),
.A2(n_692),
.B(n_766),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_833),
.B(n_682),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_881),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_822),
.B(n_698),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_838),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_898),
.B(n_737),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_883),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_978),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_927),
.B(n_754),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_916),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_817),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_893),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_960),
.B(n_721),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_858),
.B(n_754),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_927),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_887),
.B(n_721),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_833),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_833),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_927),
.B(n_754),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_866),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_932),
.A2(n_801),
.B1(n_721),
.B2(n_694),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_915),
.B(n_707),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_868),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_868),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_850),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_818),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_887),
.B(n_932),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_903),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_847),
.B(n_754),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_913),
.A2(n_757),
.B1(n_808),
.B2(n_756),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_821),
.B(n_795),
.Y(n_1020)
);

AND2x6_ASAP7_75t_SL g1021 ( 
.A(n_939),
.B(n_505),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_850),
.B(n_707),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_940),
.B(n_792),
.Y(n_1023)
);

AND2x6_ASAP7_75t_L g1024 ( 
.A(n_902),
.B(n_677),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_824),
.B(n_751),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_937),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_874),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_923),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_850),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_818),
.B(n_792),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_816),
.A2(n_741),
.B(n_736),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_873),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_844),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_SL g1034 ( 
.A(n_942),
.B(n_767),
.C(n_276),
.Y(n_1034)
);

AND2x4_ASAP7_75t_SL g1035 ( 
.A(n_975),
.B(n_792),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_875),
.B(n_877),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_878),
.B(n_735),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_825),
.A2(n_761),
.B1(n_763),
.B2(n_744),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_909),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_820),
.B(n_799),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_947),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_941),
.A2(n_741),
.B(n_736),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_902),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_903),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_882),
.B(n_735),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_839),
.A2(n_741),
.B(n_736),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_947),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_886),
.B(n_888),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_931),
.B(n_951),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_891),
.B(n_735),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_909),
.A2(n_803),
.B1(n_790),
.B2(n_707),
.Y(n_1051)
);

NOR2x1p5_ASAP7_75t_L g1052 ( 
.A(n_917),
.B(n_768),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_918),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_818),
.B(n_707),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_868),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_931),
.B(n_792),
.Y(n_1056)
);

AND2x6_ASAP7_75t_SL g1057 ( 
.A(n_951),
.B(n_507),
.Y(n_1057)
);

AND2x6_ASAP7_75t_SL g1058 ( 
.A(n_949),
.B(n_507),
.Y(n_1058)
);

AND3x1_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_511),
.C(n_510),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_919),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_962),
.Y(n_1061)
);

AOI22x1_ASAP7_75t_L g1062 ( 
.A1(n_894),
.A2(n_714),
.B1(n_715),
.B2(n_710),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_859),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_938),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_901),
.B(n_777),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_962),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_862),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_912),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_965),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_907),
.B(n_777),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_955),
.B(n_799),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_914),
.B(n_906),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_825),
.B(n_789),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_955),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_841),
.B(n_895),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_845),
.B(n_773),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_871),
.B(n_777),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_863),
.B(n_710),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_975),
.B(n_707),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_971),
.A2(n_736),
.B1(n_753),
.B2(n_779),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_895),
.B(n_714),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_937),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_920),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_971),
.A2(n_736),
.B1(n_723),
.B2(n_753),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_938),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_938),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_928),
.B(n_715),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_909),
.A2(n_803),
.B1(n_811),
.B2(n_805),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_924),
.A2(n_723),
.B1(n_729),
.B2(n_746),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_869),
.B(n_765),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_912),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_SL g1092 ( 
.A(n_889),
.B(n_679),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_867),
.B(n_870),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_975),
.B(n_729),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_922),
.B(n_738),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_865),
.A2(n_768),
.B1(n_742),
.B2(n_779),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_868),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_934),
.B(n_738),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_922),
.B(n_742),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_876),
.B(n_746),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_842),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_970),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_980),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_828),
.B(n_589),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_977),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_909),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_970),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_826),
.A2(n_750),
.B1(n_762),
.B2(n_687),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_835),
.B(n_750),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_972),
.Y(n_1110)
);

BUFx4f_ASAP7_75t_L g1111 ( 
.A(n_909),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_972),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_880),
.B(n_762),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_933),
.B(n_589),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_911),
.B(n_805),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_974),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_842),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_974),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_936),
.B(n_677),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_936),
.B(n_686),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_911),
.B(n_811),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_976),
.Y(n_1122)
);

NOR2x1p5_ASAP7_75t_L g1123 ( 
.A(n_829),
.B(n_275),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_899),
.B(n_686),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_958),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_969),
.A2(n_803),
.B1(n_725),
.B2(n_755),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_981),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_926),
.B(n_687),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_853),
.B(n_593),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_969),
.A2(n_803),
.B1(n_226),
.B2(n_651),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_981),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_819),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_943),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_869),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_826),
.B(n_688),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_926),
.B(n_688),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_819),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_L g1138 ( 
.A1(n_834),
.A2(n_705),
.B(n_765),
.C(n_690),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_823),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_823),
.Y(n_1140)
);

BUFx4f_ASAP7_75t_L g1141 ( 
.A(n_963),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_830),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_900),
.B(n_593),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_963),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_966),
.B(n_705),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_834),
.A2(n_690),
.B1(n_700),
.B2(n_755),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_904),
.B(n_948),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_830),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_836),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_836),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_852),
.B(n_741),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_979),
.B(n_700),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_840),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_892),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_950),
.B(n_391),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_852),
.B(n_831),
.Y(n_1156)
);

AND3x2_ASAP7_75t_SL g1157 ( 
.A(n_892),
.B(n_226),
.C(n_0),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_SL g1158 ( 
.A1(n_957),
.A2(n_355),
.B1(n_285),
.B2(n_296),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_959),
.B(n_278),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_840),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_843),
.B(n_703),
.Y(n_1161)
);

AO22x1_ASAP7_75t_L g1162 ( 
.A1(n_849),
.A2(n_381),
.B1(n_426),
.B2(n_425),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_843),
.B(n_703),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_846),
.B(n_704),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_846),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_987),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1156),
.A2(n_953),
.B(n_945),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1156),
.A2(n_953),
.B(n_945),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1016),
.A2(n_968),
.B(n_961),
.C(n_884),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_990),
.A2(n_999),
.B(n_1049),
.C(n_1053),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1031),
.A2(n_967),
.B(n_851),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1019),
.A2(n_848),
.B1(n_837),
.B2(n_885),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1093),
.A2(n_968),
.B(n_961),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1060),
.B(n_872),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1040),
.B(n_854),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1072),
.B(n_872),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_992),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1125),
.A2(n_879),
.B1(n_890),
.B2(n_954),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1000),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1054),
.B(n_925),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1002),
.A2(n_857),
.B(n_855),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1098),
.A2(n_973),
.B(n_930),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_1026),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1019),
.A2(n_910),
.B1(n_896),
.B2(n_908),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_982),
.B(n_964),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1012),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_995),
.A2(n_301),
.B1(n_417),
.B2(n_414),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1083),
.A2(n_856),
.B(n_861),
.C(n_864),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1005),
.A2(n_748),
.B(n_679),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_982),
.B(n_1006),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1003),
.B(n_929),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_997),
.B(n_596),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_989),
.A2(n_856),
.B(n_861),
.C(n_864),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_R g1194 ( 
.A(n_1009),
.B(n_935),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_995),
.B(n_944),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1032),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_SL g1197 ( 
.A(n_1073),
.B(n_803),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_SL g1198 ( 
.A(n_1073),
.B(n_803),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1151),
.A2(n_748),
.B(n_679),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1103),
.A2(n_389),
.B1(n_315),
.B2(n_319),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_993),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1033),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1012),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1151),
.A2(n_748),
.B(n_679),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_1018),
.A2(n_905),
.B(n_884),
.C(n_952),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1093),
.A2(n_748),
.B(n_679),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1105),
.B(n_908),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1018),
.A2(n_905),
.B(n_946),
.C(n_910),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_R g1209 ( 
.A(n_1086),
.B(n_394),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1064),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1109),
.A2(n_921),
.B(n_745),
.C(n_734),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1046),
.A2(n_760),
.B(n_748),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_994),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1023),
.B(n_329),
.C(n_312),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1105),
.B(n_921),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1026),
.Y(n_1216)
);

CKINVDCx16_ASAP7_75t_R g1217 ( 
.A(n_1085),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1133),
.B(n_704),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1023),
.B(n_343),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1036),
.B(n_706),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1027),
.B(n_346),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_985),
.A2(n_352),
.B1(n_357),
.B2(n_383),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1075),
.A2(n_760),
.B(n_708),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1056),
.B(n_596),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_985),
.A2(n_405),
.B1(n_401),
.B2(n_395),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1063),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_996),
.B(n_348),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_R g1228 ( 
.A(n_1043),
.B(n_397),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1075),
.A2(n_760),
.B(n_706),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_996),
.B(n_398),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1109),
.A2(n_708),
.B(n_713),
.C(n_745),
.Y(n_1231)
);

AOI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1147),
.A2(n_713),
.B1(n_734),
.B2(n_733),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1085),
.B(n_597),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1022),
.B(n_402),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1001),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1042),
.A2(n_760),
.B(n_725),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1001),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1138),
.A2(n_733),
.B(n_732),
.Y(n_1238)
);

NOR3xp33_ASAP7_75t_L g1239 ( 
.A(n_984),
.B(n_1071),
.C(n_1030),
.Y(n_1239)
);

O2A1O1Ixp5_ASAP7_75t_L g1240 ( 
.A1(n_1096),
.A2(n_727),
.B(n_732),
.C(n_639),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1048),
.B(n_597),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1067),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1007),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1129),
.A2(n_599),
.B(n_653),
.C(n_651),
.Y(n_1244)
);

CKINVDCx6p67_ASAP7_75t_R g1245 ( 
.A(n_1082),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1030),
.A2(n_653),
.B(n_649),
.C(n_648),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1092),
.A2(n_410),
.B(n_430),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1043),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1034),
.A2(n_649),
.B(n_648),
.C(n_645),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1143),
.B(n_599),
.Y(n_1250)
);

BUFx5_ASAP7_75t_L g1251 ( 
.A(n_1024),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1012),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_982),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1110),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1059),
.A2(n_538),
.B1(n_537),
.B2(n_536),
.Y(n_1255)
);

INVx5_ASAP7_75t_L g1256 ( 
.A(n_983),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1159),
.B(n_1014),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_988),
.A2(n_1025),
.B(n_1077),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1159),
.A2(n_645),
.B(n_639),
.C(n_628),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1029),
.B(n_412),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1058),
.B(n_418),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1021),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1022),
.B(n_421),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1076),
.A2(n_427),
.B1(n_431),
.B2(n_803),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1095),
.A2(n_588),
.B(n_628),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1154),
.B(n_605),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1098),
.A2(n_646),
.B(n_625),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1099),
.A2(n_618),
.B(n_605),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1022),
.B(n_618),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1114),
.B(n_624),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1134),
.B(n_624),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1012),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1013),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1057),
.B(n_1),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1104),
.B(n_592),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1054),
.B(n_592),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1112),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1054),
.B(n_621),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1074),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1141),
.A2(n_542),
.B1(n_511),
.B2(n_515),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_R g1281 ( 
.A(n_1097),
.B(n_86),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1130),
.A2(n_558),
.B1(n_557),
.B2(n_510),
.Y(n_1282)
);

AND2x6_ASAP7_75t_L g1283 ( 
.A(n_1079),
.B(n_515),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1028),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1035),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1013),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1141),
.A2(n_543),
.B1(n_523),
.B2(n_527),
.Y(n_1287)
);

AND3x1_ASAP7_75t_SL g1288 ( 
.A(n_1123),
.B(n_558),
.C(n_557),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1015),
.A2(n_542),
.B(n_523),
.C(n_527),
.Y(n_1289)
);

NOR2x1_ASAP7_75t_L g1290 ( 
.A(n_998),
.B(n_517),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1015),
.B(n_1158),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1011),
.B(n_621),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1017),
.B(n_1044),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_991),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1011),
.A2(n_646),
.B1(n_625),
.B2(n_543),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1013),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1017),
.B(n_1),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1088),
.A2(n_538),
.B1(n_555),
.B2(n_554),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_L g1300 ( 
.A(n_1144),
.B(n_517),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1155),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1088),
.A2(n_546),
.B1(n_555),
.B2(n_554),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1038),
.A2(n_986),
.B(n_1010),
.C(n_1101),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1013),
.Y(n_1304)
);

AOI221xp5_ASAP7_75t_L g1305 ( 
.A1(n_1130),
.A2(n_537),
.B1(n_553),
.B2(n_550),
.C(n_546),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1055),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1118),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1152),
.A2(n_556),
.B(n_553),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_983),
.A2(n_1004),
.B(n_1128),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_991),
.B(n_528),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_983),
.A2(n_550),
.B(n_536),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_991),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1146),
.A2(n_532),
.B(n_530),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1238),
.A2(n_1124),
.B(n_1062),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1179),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1258),
.A2(n_1121),
.B(n_1115),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1201),
.B(n_1162),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1239),
.A2(n_1052),
.B1(n_1035),
.B2(n_1079),
.Y(n_1318)
);

O2A1O1Ixp5_ASAP7_75t_L g1319 ( 
.A1(n_1219),
.A2(n_1081),
.B(n_1106),
.C(n_1111),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1267),
.A2(n_1124),
.B(n_1113),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1205),
.A2(n_1087),
.B(n_1145),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1171),
.A2(n_1004),
.B(n_1106),
.Y(n_1322)
);

CKINVDCx14_ASAP7_75t_R g1323 ( 
.A(n_1196),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1167),
.A2(n_1004),
.B(n_1111),
.Y(n_1324)
);

NOR3xp33_ASAP7_75t_SL g1325 ( 
.A(n_1262),
.B(n_1008),
.C(n_998),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1224),
.B(n_1094),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1250),
.B(n_1041),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1236),
.A2(n_1100),
.B(n_1113),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_SL g1329 ( 
.A(n_1261),
.B(n_1155),
.C(n_1020),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1177),
.B(n_1122),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1168),
.A2(n_1081),
.B(n_1135),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1270),
.B(n_1068),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1274),
.A2(n_1157),
.B(n_1080),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1257),
.A2(n_1084),
.B(n_1089),
.C(n_1094),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1231),
.A2(n_1108),
.A3(n_1136),
.B(n_1078),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1166),
.B(n_1008),
.Y(n_1336)
);

AO32x2_ASAP7_75t_L g1337 ( 
.A1(n_1282),
.A2(n_1157),
.A3(n_1090),
.B1(n_1135),
.B2(n_1126),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1206),
.A2(n_1100),
.B(n_1164),
.Y(n_1338)
);

NAND2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1194),
.B(n_1117),
.Y(n_1339)
);

INVx6_ASAP7_75t_L g1340 ( 
.A(n_1217),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1169),
.A2(n_1117),
.B(n_1144),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1197),
.A2(n_1039),
.B(n_1051),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1214),
.A2(n_1144),
.B1(n_1091),
.B2(n_1097),
.Y(n_1343)
);

BUFx4f_ASAP7_75t_L g1344 ( 
.A(n_1216),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1175),
.B(n_1091),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1256),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1256),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1197),
.A2(n_1039),
.B(n_1051),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1212),
.A2(n_1090),
.B(n_1065),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1184),
.A2(n_1050),
.A3(n_1045),
.B(n_1037),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1235),
.B(n_1144),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1256),
.B(n_1055),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1172),
.A2(n_1070),
.B(n_1137),
.C(n_1132),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1210),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1291),
.A2(n_1119),
.B1(n_1120),
.B2(n_1024),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1213),
.Y(n_1356)
);

BUFx10_ASAP7_75t_L g1357 ( 
.A(n_1221),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1256),
.B(n_1285),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1241),
.B(n_1041),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1259),
.A2(n_1165),
.B(n_1127),
.C(n_1131),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1237),
.B(n_1140),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1301),
.A2(n_1263),
.B1(n_1234),
.B2(n_1230),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1198),
.A2(n_1039),
.B(n_1161),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1193),
.A2(n_1055),
.B(n_1119),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1189),
.A2(n_1163),
.B(n_1047),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1252),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1223),
.A2(n_1047),
.B(n_1061),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1181),
.A2(n_1102),
.B(n_1061),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1190),
.B(n_1055),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1266),
.A2(n_1039),
.B1(n_1160),
.B2(n_1153),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1190),
.B(n_1119),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1252),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1198),
.A2(n_1120),
.B(n_1149),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1271),
.B(n_1148),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1229),
.A2(n_1150),
.B(n_1149),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1240),
.A2(n_1150),
.B(n_1142),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1176),
.B(n_1066),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1275),
.B(n_1069),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1222),
.A2(n_528),
.B1(n_530),
.B2(n_532),
.C(n_1107),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1202),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1192),
.B(n_1207),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1199),
.A2(n_1120),
.B(n_1139),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1184),
.A2(n_1142),
.A3(n_1139),
.B(n_1107),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1204),
.A2(n_1102),
.B(n_1069),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1253),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1182),
.A2(n_1024),
.B(n_218),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1294),
.B(n_3),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1173),
.A2(n_1024),
.B(n_187),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1232),
.A2(n_184),
.B(n_181),
.Y(n_1389)
);

NAND3x1_ASAP7_75t_L g1390 ( 
.A(n_1227),
.B(n_3),
.C(n_10),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1309),
.A2(n_161),
.B(n_157),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1248),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1195),
.A2(n_111),
.B(n_104),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1215),
.B(n_12),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1295),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1226),
.B(n_14),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1244),
.A2(n_15),
.A3(n_18),
.B(n_20),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1249),
.B(n_20),
.C(n_21),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1242),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1308),
.A2(n_99),
.B(n_94),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1245),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1265),
.A2(n_93),
.B(n_23),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1208),
.A2(n_22),
.B(n_26),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1312),
.B(n_26),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1285),
.A2(n_1178),
.B1(n_1254),
.B2(n_1277),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1296),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1268),
.A2(n_27),
.B(n_30),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1248),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1307),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1313),
.A2(n_27),
.B(n_31),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1174),
.B(n_1284),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1298),
.A2(n_32),
.A3(n_33),
.B(n_34),
.Y(n_1412)
);

O2A1O1Ixp5_ASAP7_75t_L g1413 ( 
.A1(n_1247),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1233),
.B(n_35),
.Y(n_1414)
);

AND2x6_ASAP7_75t_L g1415 ( 
.A(n_1252),
.B(n_37),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1188),
.A2(n_38),
.B(n_46),
.C(n_47),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1246),
.A2(n_46),
.B(n_48),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1220),
.A2(n_51),
.B(n_53),
.Y(n_1418)
);

NAND2xp33_ASAP7_75t_L g1419 ( 
.A(n_1283),
.B(n_60),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1233),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1280),
.A2(n_60),
.A3(n_62),
.B(n_63),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1185),
.B(n_63),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1191),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1290),
.A2(n_64),
.B(n_66),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1300),
.A2(n_68),
.B(n_69),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1185),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1218),
.Y(n_1427)
);

AO31x2_ASAP7_75t_L g1428 ( 
.A1(n_1280),
.A2(n_73),
.A3(n_75),
.B(n_76),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1310),
.Y(n_1429)
);

AOI31xp67_ASAP7_75t_L g1430 ( 
.A1(n_1264),
.A2(n_73),
.A3(n_76),
.B(n_77),
.Y(n_1430)
);

OAI22x1_ASAP7_75t_L g1431 ( 
.A1(n_1180),
.A2(n_84),
.B1(n_77),
.B2(n_80),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1292),
.A2(n_84),
.B(n_1293),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1289),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1276),
.A2(n_1278),
.B(n_1269),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1222),
.A2(n_1225),
.B(n_1287),
.C(n_1243),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1260),
.A2(n_1225),
.B(n_1311),
.C(n_1287),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1283),
.B(n_1306),
.Y(n_1437)
);

NOR4xp25_ASAP7_75t_L g1438 ( 
.A(n_1305),
.B(n_1302),
.C(n_1299),
.D(n_1187),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1186),
.A2(n_1273),
.B(n_1304),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1299),
.A2(n_1302),
.B(n_1283),
.Y(n_1440)
);

CKINVDCx8_ASAP7_75t_R g1441 ( 
.A(n_1248),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1228),
.B(n_1279),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1203),
.A2(n_1233),
.B(n_1251),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1251),
.A2(n_1272),
.B(n_1286),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1251),
.A2(n_1272),
.B(n_1286),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1183),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1255),
.A2(n_1297),
.B1(n_1272),
.B2(n_1286),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1200),
.B(n_1297),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1251),
.A2(n_1288),
.B(n_1297),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1251),
.A2(n_1281),
.B(n_1209),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1183),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1256),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1231),
.A2(n_1211),
.A3(n_1168),
.B(n_1167),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1170),
.B(n_999),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1177),
.B(n_1003),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1222),
.A2(n_939),
.B1(n_990),
.B2(n_767),
.C(n_671),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1238),
.A2(n_1267),
.B(n_1236),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1303),
.A2(n_1212),
.B(n_1236),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1250),
.B(n_1016),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1238),
.A2(n_1267),
.B(n_1236),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1224),
.B(n_1003),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1170),
.B(n_999),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1177),
.B(n_1003),
.Y(n_1463)
);

O2A1O1Ixp5_ASAP7_75t_L g1464 ( 
.A1(n_1219),
.A2(n_1016),
.B(n_845),
.C(n_1073),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1170),
.A2(n_1016),
.B(n_999),
.C(n_990),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1248),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1258),
.A2(n_927),
.B(n_1016),
.Y(n_1467)
);

AO21x1_ASAP7_75t_L g1468 ( 
.A1(n_1258),
.A2(n_1016),
.B(n_989),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1238),
.A2(n_1267),
.B(n_1236),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1468),
.A2(n_1458),
.B(n_1388),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1370),
.A2(n_1416),
.A3(n_1467),
.B(n_1331),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1347),
.Y(n_1472)
);

BUFx2_ASAP7_75t_R g1473 ( 
.A(n_1441),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1356),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1456),
.A2(n_1362),
.B1(n_1329),
.B2(n_1333),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1341),
.A2(n_1348),
.B(n_1342),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1354),
.Y(n_1478)
);

AND2x4_ASAP7_75t_SL g1479 ( 
.A(n_1466),
.B(n_1347),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1365),
.A2(n_1322),
.B(n_1314),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1328),
.A2(n_1338),
.B(n_1384),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1333),
.B(n_1459),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1374),
.A2(n_1459),
.B1(n_1318),
.B2(n_1355),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1367),
.A2(n_1375),
.B(n_1324),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1315),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1401),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1376),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1346),
.B(n_1452),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1381),
.B(n_1461),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1420),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1323),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1462),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1407),
.A2(n_1398),
.B1(n_1417),
.B2(n_1395),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1370),
.A2(n_1353),
.A3(n_1465),
.B(n_1382),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1376),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1407),
.A2(n_1398),
.B1(n_1417),
.B2(n_1395),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1386),
.A2(n_1368),
.B(n_1320),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1357),
.A2(n_1405),
.B1(n_1326),
.B2(n_1463),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1357),
.A2(n_1405),
.B1(n_1455),
.B2(n_1448),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1451),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1389),
.A2(n_1391),
.B(n_1410),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1339),
.A2(n_1419),
.B1(n_1390),
.B2(n_1336),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1356),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1403),
.A2(n_1316),
.B(n_1373),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1446),
.Y(n_1505)
);

CKINVDCx8_ASAP7_75t_R g1506 ( 
.A(n_1466),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1316),
.A2(n_1363),
.B(n_1443),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1443),
.A2(n_1393),
.B(n_1364),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1402),
.A2(n_1464),
.B(n_1413),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1330),
.B(n_1385),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1392),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1380),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1399),
.Y(n_1513)
);

BUFx2_ASAP7_75t_SL g1514 ( 
.A(n_1408),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1451),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1440),
.A2(n_1431),
.B1(n_1414),
.B2(n_1425),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_SL g1517 ( 
.A1(n_1435),
.A2(n_1440),
.B(n_1450),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1444),
.A2(n_1445),
.B(n_1400),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1414),
.A2(n_1396),
.B1(n_1394),
.B2(n_1317),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1406),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1321),
.A2(n_1439),
.B(n_1319),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1321),
.A2(n_1377),
.B(n_1432),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1424),
.A2(n_1360),
.B(n_1436),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1344),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1349),
.A2(n_1334),
.B(n_1438),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1409),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1438),
.A2(n_1433),
.B(n_1377),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1427),
.B(n_1385),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1411),
.B(n_1426),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1345),
.A2(n_1359),
.B(n_1437),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1378),
.A2(n_1434),
.B(n_1327),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1411),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1327),
.A2(n_1447),
.B(n_1332),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1418),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1387),
.B(n_1404),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1418),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1447),
.A2(n_1369),
.B(n_1352),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1352),
.A2(n_1351),
.B(n_1343),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1429),
.A2(n_1325),
.B1(n_1442),
.B2(n_1361),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1358),
.A2(n_1371),
.B(n_1372),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1422),
.B(n_1379),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1340),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1366),
.B(n_1372),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1366),
.A2(n_1453),
.B(n_1383),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1344),
.B(n_1415),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1423),
.B(n_1340),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1453),
.A2(n_1335),
.B(n_1350),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1414),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1397),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1453),
.A2(n_1350),
.B(n_1430),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1397),
.B(n_1415),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1350),
.A2(n_1337),
.B(n_1335),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1415),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1415),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1335),
.A2(n_1337),
.B(n_1397),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1412),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1412),
.A2(n_1421),
.B(n_1428),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1356),
.Y(n_1558)
);

NAND2x1p5_ASAP7_75t_L g1559 ( 
.A(n_1347),
.B(n_1256),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_SL g1560 ( 
.A1(n_1436),
.A2(n_1016),
.B(n_1416),
.C(n_1465),
.Y(n_1560)
);

INVx4_ASAP7_75t_SL g1561 ( 
.A(n_1415),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1461),
.B(n_1326),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1315),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1376),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1364),
.B(n_1341),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1347),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1456),
.A2(n_1016),
.B1(n_990),
.B2(n_1407),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1466),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1456),
.A2(n_939),
.B1(n_990),
.B2(n_932),
.C(n_916),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1374),
.A2(n_1016),
.B1(n_999),
.B2(n_995),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1315),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1464),
.A2(n_1016),
.B(n_999),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1441),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1441),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1464),
.A2(n_1016),
.B(n_999),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1315),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1464),
.A2(n_1016),
.B(n_999),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1456),
.A2(n_1016),
.B1(n_990),
.B2(n_1407),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1323),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1333),
.A2(n_1016),
.B1(n_1456),
.B2(n_999),
.Y(n_1583)
);

NOR2xp67_ASAP7_75t_L g1584 ( 
.A(n_1329),
.B(n_1196),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1333),
.B(n_1016),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1586)
);

AO21x1_ASAP7_75t_L g1587 ( 
.A1(n_1417),
.A2(n_1016),
.B(n_1407),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_R g1588 ( 
.A(n_1339),
.B(n_1009),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1456),
.A2(n_1016),
.B(n_990),
.C(n_1440),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1347),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1364),
.B(n_1341),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1456),
.A2(n_1016),
.B1(n_990),
.B2(n_1407),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1315),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1315),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1315),
.Y(n_1596)
);

AO21x2_ASAP7_75t_L g1597 ( 
.A1(n_1468),
.A2(n_1458),
.B(n_1388),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1441),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_SL g1599 ( 
.A(n_1405),
.B(n_902),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1333),
.B(n_1016),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1376),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1374),
.A2(n_1016),
.B1(n_999),
.B2(n_995),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1456),
.B(n_1016),
.C(n_932),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1315),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1315),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1443),
.B(n_1426),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1374),
.A2(n_1016),
.B1(n_999),
.B2(n_995),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1456),
.A2(n_1016),
.B(n_990),
.C(n_1440),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1323),
.Y(n_1609)
);

OAI21xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1440),
.A2(n_1016),
.B(n_1342),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1464),
.A2(n_1016),
.B(n_999),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1456),
.A2(n_1016),
.B(n_990),
.C(n_1440),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1376),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1333),
.B(n_1016),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1456),
.A2(n_1016),
.B1(n_990),
.B2(n_1407),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_SL g1616 ( 
.A1(n_1407),
.A2(n_1449),
.B(n_1443),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1383),
.Y(n_1617)
);

OAI211xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1456),
.A2(n_940),
.B(n_898),
.C(n_999),
.Y(n_1618)
);

OR2x6_ASAP7_75t_L g1619 ( 
.A(n_1364),
.B(n_1341),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1460),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1347),
.B(n_1256),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1485),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1515),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1515),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1510),
.B(n_1489),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1492),
.B(n_1482),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1562),
.B(n_1482),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1492),
.B(n_1532),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1569),
.A2(n_1583),
.B1(n_1603),
.B2(n_1493),
.C(n_1496),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1585),
.B(n_1600),
.Y(n_1630)
);

AND2x6_ASAP7_75t_L g1631 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1585),
.B(n_1600),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1614),
.B(n_1529),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1547),
.A2(n_1504),
.B(n_1557),
.Y(n_1634)
);

O2A1O1Ixp5_ASAP7_75t_L g1635 ( 
.A1(n_1587),
.A2(n_1614),
.B(n_1608),
.C(n_1612),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1583),
.B(n_1570),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1474),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_SL g1638 ( 
.A1(n_1589),
.A2(n_1612),
.B(n_1608),
.Y(n_1638)
);

O2A1O1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1589),
.A2(n_1560),
.B(n_1607),
.C(n_1602),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1476),
.A2(n_1592),
.B(n_1565),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1503),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1573),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1527),
.B(n_1483),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1547),
.A2(n_1504),
.B(n_1484),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1535),
.B(n_1528),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1478),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1475),
.B(n_1519),
.Y(n_1647)
);

OA22x2_ASAP7_75t_L g1648 ( 
.A1(n_1502),
.A2(n_1499),
.B1(n_1498),
.B2(n_1539),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1505),
.Y(n_1649)
);

NOR2xp67_ASAP7_75t_L g1650 ( 
.A(n_1542),
.B(n_1500),
.Y(n_1650)
);

AOI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1519),
.A2(n_1618),
.B(n_1560),
.C(n_1610),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1558),
.B(n_1567),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1561),
.B(n_1606),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1493),
.A2(n_1496),
.B1(n_1578),
.B2(n_1567),
.Y(n_1654)
);

NOR2xp67_ASAP7_75t_L g1655 ( 
.A(n_1542),
.B(n_1486),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1511),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1512),
.Y(n_1657)
);

OA21x2_ASAP7_75t_L g1658 ( 
.A1(n_1522),
.A2(n_1497),
.B(n_1481),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1578),
.B(n_1593),
.Y(n_1659)
);

O2A1O1Ixp5_ASAP7_75t_L g1660 ( 
.A1(n_1572),
.A2(n_1575),
.B(n_1577),
.C(n_1611),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1513),
.Y(n_1661)
);

O2A1O1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1593),
.A2(n_1615),
.B(n_1541),
.C(n_1546),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1565),
.A2(n_1619),
.B(n_1592),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1615),
.A2(n_1517),
.B(n_1516),
.C(n_1545),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1527),
.B(n_1530),
.Y(n_1665)
);

AND2x6_ASAP7_75t_L g1666 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1516),
.A2(n_1619),
.B1(n_1553),
.B2(n_1545),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1551),
.B(n_1553),
.Y(n_1668)
);

BUFx12f_ASAP7_75t_L g1669 ( 
.A(n_1478),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1520),
.A2(n_1595),
.B1(n_1563),
.B2(n_1576),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1584),
.A2(n_1524),
.B1(n_1548),
.B2(n_1491),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1526),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1514),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1559),
.A2(n_1621),
.B(n_1599),
.Y(n_1674)
);

AND2x4_ASAP7_75t_SL g1675 ( 
.A(n_1505),
.B(n_1491),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1525),
.B(n_1571),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1537),
.B(n_1533),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1594),
.B(n_1596),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1604),
.B(n_1605),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1543),
.B(n_1568),
.Y(n_1680)
);

NAND2x1_ASAP7_75t_L g1681 ( 
.A(n_1616),
.B(n_1566),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1540),
.B(n_1479),
.Y(n_1682)
);

OAI211xp5_ASAP7_75t_L g1683 ( 
.A1(n_1588),
.A2(n_1509),
.B(n_1490),
.C(n_1536),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1473),
.A2(n_1598),
.B1(n_1574),
.B2(n_1573),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1574),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1598),
.A2(n_1506),
.B1(n_1524),
.B2(n_1556),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1540),
.B(n_1479),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1534),
.B(n_1549),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1588),
.B(n_1488),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1531),
.B(n_1591),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1509),
.A2(n_1552),
.B1(n_1609),
.B2(n_1580),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1617),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1490),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1509),
.A2(n_1552),
.B1(n_1609),
.B2(n_1580),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1486),
.Y(n_1695)
);

AOI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1507),
.A2(n_1508),
.B(n_1555),
.C(n_1538),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1472),
.B(n_1544),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1487),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1552),
.A2(n_1523),
.B1(n_1559),
.B2(n_1621),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1494),
.B(n_1471),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1494),
.B(n_1471),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1494),
.B(n_1471),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1523),
.B(n_1471),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1487),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1470),
.B(n_1597),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1501),
.A2(n_1521),
.B(n_1518),
.C(n_1480),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1550),
.A2(n_1601),
.B1(n_1495),
.B2(n_1613),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1521),
.B(n_1564),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1477),
.A2(n_1579),
.B(n_1581),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1620),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1582),
.B(n_1586),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1590),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1561),
.B(n_1606),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1562),
.B(n_1482),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1562),
.B(n_1482),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1510),
.Y(n_1716)
);

O2A1O1Ixp5_ASAP7_75t_L g1717 ( 
.A1(n_1587),
.A2(n_1016),
.B(n_1464),
.C(n_1417),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1492),
.B(n_1482),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1510),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1505),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1506),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1493),
.A2(n_1496),
.B1(n_1578),
.B2(n_1567),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1510),
.B(n_1489),
.Y(n_1723)
);

O2A1O1Ixp5_ASAP7_75t_L g1724 ( 
.A1(n_1587),
.A2(n_1016),
.B(n_1464),
.C(n_1417),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1505),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1515),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1562),
.B(n_1482),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1562),
.B(n_1482),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1492),
.B(n_1489),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1475),
.A2(n_1585),
.B1(n_1614),
.B2(n_1600),
.Y(n_1730)
);

O2A1O1Ixp5_ASAP7_75t_L g1731 ( 
.A1(n_1587),
.A2(n_1016),
.B(n_1464),
.C(n_1417),
.Y(n_1731)
);

AND2x6_ASAP7_75t_L g1732 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1476),
.A2(n_1016),
.B(n_1603),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_SL g1734 ( 
.A1(n_1589),
.A2(n_902),
.B(n_1073),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1561),
.B(n_1606),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1493),
.A2(n_1496),
.B1(n_1578),
.B2(n_1567),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1506),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1562),
.B(n_1482),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_SL g1739 ( 
.A1(n_1585),
.A2(n_845),
.B(n_1614),
.C(n_1600),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1589),
.A2(n_902),
.B(n_1073),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1506),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1515),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1703),
.B(n_1704),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1692),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1676),
.B(n_1643),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1688),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1708),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1698),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1676),
.B(n_1643),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1716),
.Y(n_1751)
);

AND2x4_ASAP7_75t_SL g1752 ( 
.A(n_1668),
.B(n_1653),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1665),
.B(n_1700),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1730),
.A2(n_1629),
.B1(n_1722),
.B2(n_1736),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1622),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1665),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1733),
.A2(n_1724),
.B(n_1717),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1630),
.B(n_1632),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1627),
.B(n_1714),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1711),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1715),
.B(n_1727),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1654),
.A2(n_1736),
.B(n_1722),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1626),
.B(n_1718),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1705),
.B(n_1701),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1702),
.B(n_1691),
.Y(n_1765)
);

OAI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1651),
.A2(n_1647),
.B(n_1638),
.C(n_1639),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1738),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_L g1768 ( 
.A(n_1683),
.B(n_1690),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1682),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1707),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1626),
.B(n_1718),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1729),
.B(n_1625),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1628),
.B(n_1633),
.Y(n_1773)
);

OR2x6_ASAP7_75t_L g1774 ( 
.A(n_1640),
.B(n_1663),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1657),
.B(n_1661),
.Y(n_1775)
);

OA21x2_ASAP7_75t_L g1776 ( 
.A1(n_1731),
.A2(n_1660),
.B(n_1635),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1651),
.B(n_1662),
.C(n_1739),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1628),
.B(n_1716),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1654),
.A2(n_1648),
.B1(n_1659),
.B2(n_1636),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1709),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1709),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1696),
.B(n_1712),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1719),
.B(n_1672),
.Y(n_1783)
);

CKINVDCx16_ASAP7_75t_R g1784 ( 
.A(n_1693),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1678),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1723),
.B(n_1645),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1664),
.B(n_1667),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1678),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1687),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1694),
.B(n_1677),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1637),
.B(n_1641),
.Y(n_1791)
);

NOR2xp67_ASAP7_75t_SL g1792 ( 
.A(n_1734),
.B(n_1740),
.Y(n_1792)
);

INVx4_ASAP7_75t_L g1793 ( 
.A(n_1631),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1634),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1649),
.B(n_1720),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1697),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1634),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1668),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1699),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1696),
.B(n_1653),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1670),
.B(n_1679),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1670),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1658),
.Y(n_1803)
);

OR2x6_ASAP7_75t_L g1804 ( 
.A(n_1674),
.B(n_1681),
.Y(n_1804)
);

AO21x2_ASAP7_75t_L g1805 ( 
.A1(n_1667),
.A2(n_1652),
.B(n_1686),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1713),
.B(n_1735),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1644),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1656),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1648),
.B(n_1686),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1631),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1769),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1744),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1744),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1744),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1780),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1751),
.B(n_1671),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1755),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1764),
.B(n_1760),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1793),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1760),
.B(n_1746),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1751),
.B(n_1689),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1760),
.B(n_1746),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1811),
.B(n_1685),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1811),
.B(n_1642),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1811),
.B(n_1673),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1754),
.A2(n_1669),
.B1(n_1732),
.B2(n_1631),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1745),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1745),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1750),
.B(n_1684),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1791),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1774),
.B(n_1655),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1743),
.B(n_1748),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1791),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1781),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1763),
.B(n_1666),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1756),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1749),
.Y(n_1838)
);

OAI21xp33_ASAP7_75t_L g1839 ( 
.A1(n_1762),
.A2(n_1779),
.B(n_1777),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1771),
.B(n_1666),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1756),
.Y(n_1841)
);

OAI33xp33_ASAP7_75t_L g1842 ( 
.A1(n_1777),
.A2(n_1684),
.A3(n_1646),
.B1(n_1695),
.B2(n_1650),
.B3(n_1666),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1750),
.B(n_1741),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1796),
.B(n_1623),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1804),
.Y(n_1845)
);

INVx5_ASAP7_75t_L g1846 ( 
.A(n_1774),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1775),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1796),
.B(n_1624),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1783),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_L g1850 ( 
.A(n_1774),
.B(n_1741),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1786),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1772),
.B(n_1675),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1778),
.B(n_1721),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1753),
.B(n_1721),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1778),
.B(n_1737),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1775),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1762),
.A2(n_1737),
.B1(n_1725),
.B2(n_1726),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1813),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1839),
.A2(n_1787),
.B1(n_1792),
.B2(n_1809),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1813),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1814),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1857),
.A2(n_1766),
.B1(n_1809),
.B2(n_1793),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1845),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1838),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1819),
.B(n_1782),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1839),
.A2(n_1787),
.B1(n_1792),
.B2(n_1805),
.Y(n_1866)
);

INVx3_ASAP7_75t_SL g1867 ( 
.A(n_1845),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1816),
.A2(n_1803),
.B(n_1797),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1842),
.A2(n_1766),
.B1(n_1757),
.B2(n_1773),
.C(n_1801),
.Y(n_1869)
);

INVx8_ASAP7_75t_L g1870 ( 
.A(n_1848),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1849),
.B(n_1831),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1833),
.B(n_1782),
.Y(n_1872)
);

AOI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1832),
.A2(n_1807),
.B(n_1768),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1826),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1837),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1815),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1834),
.B(n_1758),
.Y(n_1877)
);

NAND3xp33_ASAP7_75t_L g1878 ( 
.A(n_1857),
.B(n_1757),
.C(n_1776),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1827),
.A2(n_1784),
.B1(n_1749),
.B2(n_1793),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1826),
.A2(n_1805),
.B1(n_1774),
.B2(n_1768),
.Y(n_1880)
);

INVx5_ASAP7_75t_SL g1881 ( 
.A(n_1845),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1851),
.A2(n_1773),
.B1(n_1801),
.B2(n_1770),
.C(n_1758),
.Y(n_1882)
);

AOI211xp5_ASAP7_75t_L g1883 ( 
.A1(n_1830),
.A2(n_1799),
.B(n_1790),
.C(n_1765),
.Y(n_1883)
);

NOR3xp33_ASAP7_75t_SL g1884 ( 
.A(n_1817),
.B(n_1784),
.C(n_1795),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1850),
.A2(n_1774),
.B1(n_1805),
.B2(n_1793),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1853),
.A2(n_1770),
.B1(n_1808),
.B2(n_1799),
.C(n_1783),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1830),
.A2(n_1805),
.B1(n_1774),
.B2(n_1800),
.Y(n_1887)
);

OAI33xp33_ASAP7_75t_L g1888 ( 
.A1(n_1855),
.A2(n_1753),
.A3(n_1802),
.B1(n_1747),
.B2(n_1785),
.B3(n_1788),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1844),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1822),
.A2(n_1808),
.B1(n_1767),
.B2(n_1761),
.C(n_1759),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1843),
.B(n_1785),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1852),
.B(n_1759),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1843),
.Y(n_1893)
);

AOI33xp33_ASAP7_75t_L g1894 ( 
.A1(n_1838),
.A2(n_1788),
.A3(n_1802),
.B1(n_1747),
.B2(n_1761),
.B3(n_1767),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1818),
.Y(n_1895)
);

AO21x2_ASAP7_75t_L g1896 ( 
.A1(n_1835),
.A2(n_1794),
.B(n_1797),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1812),
.B(n_1789),
.Y(n_1897)
);

CKINVDCx20_ASAP7_75t_R g1898 ( 
.A(n_1836),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1841),
.Y(n_1899)
);

NAND3xp33_ASAP7_75t_L g1900 ( 
.A(n_1832),
.B(n_1776),
.C(n_1846),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1840),
.A2(n_1810),
.B1(n_1798),
.B2(n_1752),
.Y(n_1901)
);

INVxp67_ASAP7_75t_SL g1902 ( 
.A(n_1828),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1829),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1818),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1858),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1861),
.B(n_1821),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1882),
.B(n_1847),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1895),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1895),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1863),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1868),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_R g1912 ( 
.A(n_1884),
.B(n_1776),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1864),
.Y(n_1913)
);

AND4x1_ASAP7_75t_L g1914 ( 
.A(n_1866),
.B(n_1824),
.C(n_1825),
.D(n_1806),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1859),
.B(n_1878),
.C(n_1869),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1886),
.B(n_1847),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1896),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1894),
.B(n_1846),
.Y(n_1918)
);

OR2x6_ASAP7_75t_L g1919 ( 
.A(n_1900),
.B(n_1804),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1904),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1896),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1870),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1860),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1885),
.A2(n_1862),
.B(n_1804),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1873),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1902),
.B(n_1856),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1860),
.Y(n_1927)
);

INVx4_ASAP7_75t_SL g1928 ( 
.A(n_1867),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1875),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1867),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1899),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1870),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1865),
.B(n_1824),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1876),
.B(n_1821),
.Y(n_1934)
);

BUFx8_ASAP7_75t_L g1935 ( 
.A(n_1863),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1872),
.B(n_1825),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1867),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1863),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1905),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1911),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1918),
.B(n_1929),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1918),
.B(n_1903),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1915),
.A2(n_1879),
.B1(n_1887),
.B2(n_1880),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1913),
.B(n_1890),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1913),
.B(n_1883),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1915),
.B(n_1892),
.Y(n_1946)
);

NAND4xp25_ASAP7_75t_L g1947 ( 
.A(n_1912),
.B(n_1854),
.C(n_1871),
.D(n_1901),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1905),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1928),
.B(n_1872),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1928),
.B(n_1863),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1908),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1928),
.B(n_1863),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1928),
.B(n_1881),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1929),
.B(n_1893),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1909),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1931),
.B(n_1891),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1911),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1907),
.B(n_1898),
.Y(n_1958)
);

INVx5_ASAP7_75t_L g1959 ( 
.A(n_1925),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1907),
.B(n_1874),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1937),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1916),
.B(n_1877),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1928),
.B(n_1930),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1937),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1928),
.B(n_1881),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1920),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1911),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1930),
.B(n_1881),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1930),
.B(n_1889),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1931),
.B(n_1823),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1935),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1937),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1930),
.B(n_1881),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1933),
.B(n_1897),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1911),
.Y(n_1975)
);

INVx5_ASAP7_75t_L g1976 ( 
.A(n_1925),
.Y(n_1976)
);

OR2x6_ASAP7_75t_L g1977 ( 
.A(n_1924),
.B(n_1910),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1911),
.Y(n_1978)
);

INVx4_ASAP7_75t_L g1979 ( 
.A(n_1938),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1936),
.B(n_1922),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1923),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1923),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1922),
.B(n_1898),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1951),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1951),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_SL g1986 ( 
.A(n_1953),
.B(n_1965),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1954),
.B(n_1906),
.Y(n_1987)
);

NOR2xp67_ASAP7_75t_SL g1988 ( 
.A(n_1959),
.B(n_1624),
.Y(n_1988)
);

OA21x2_ASAP7_75t_L g1989 ( 
.A1(n_1972),
.A2(n_1921),
.B(n_1917),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1955),
.Y(n_1990)
);

OR2x6_ASAP7_75t_L g1991 ( 
.A(n_1977),
.B(n_1925),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1963),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1963),
.Y(n_1993)
);

OAI21xp33_ASAP7_75t_L g1994 ( 
.A1(n_1946),
.A2(n_1914),
.B(n_1919),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1979),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1954),
.B(n_1906),
.Y(n_1996)
);

NAND2x1_ASAP7_75t_L g1997 ( 
.A(n_1977),
.B(n_1910),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1955),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1953),
.B(n_1910),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1956),
.B(n_1934),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_SL g2001 ( 
.A(n_1965),
.B(n_1820),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1949),
.B(n_1910),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1979),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1949),
.B(n_1910),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1950),
.B(n_1922),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1966),
.Y(n_2006)
);

OAI21xp33_ASAP7_75t_L g2007 ( 
.A1(n_1943),
.A2(n_1914),
.B(n_1919),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1956),
.B(n_1934),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1979),
.Y(n_2009)
);

NAND2x1p5_ASAP7_75t_L g2010 ( 
.A(n_1959),
.B(n_1925),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1958),
.B(n_1936),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_L g2012 ( 
.A(n_1961),
.B(n_1888),
.C(n_1932),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1945),
.B(n_1926),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1977),
.B(n_1938),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1959),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1966),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1964),
.B(n_1934),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1941),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1977),
.B(n_1925),
.Y(n_2019)
);

INVxp67_ASAP7_75t_L g2020 ( 
.A(n_1944),
.Y(n_2020)
);

NOR4xp25_ASAP7_75t_L g2021 ( 
.A(n_1947),
.B(n_1926),
.C(n_1932),
.D(n_1927),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1950),
.B(n_1938),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1952),
.B(n_1938),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1981),
.Y(n_2024)
);

INVxp67_ASAP7_75t_SL g2025 ( 
.A(n_1941),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1981),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_2010),
.Y(n_2027)
);

BUFx2_ASAP7_75t_R g2028 ( 
.A(n_2013),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2022),
.B(n_1980),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_2007),
.A2(n_1919),
.B1(n_1973),
.B2(n_1968),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1994),
.B(n_1969),
.Y(n_2031)
);

NAND2xp33_ASAP7_75t_L g2032 ( 
.A(n_2019),
.B(n_1942),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2022),
.B(n_1980),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2023),
.B(n_1952),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2023),
.B(n_1968),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_2020),
.A2(n_1919),
.B1(n_1973),
.B2(n_1969),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_1993),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_2018),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2002),
.B(n_1969),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2025),
.B(n_1962),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1984),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2002),
.B(n_1974),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2021),
.B(n_1960),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1992),
.B(n_1939),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1992),
.B(n_2012),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_1999),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2004),
.B(n_1974),
.Y(n_2047)
);

INVxp67_ASAP7_75t_L g2048 ( 
.A(n_1986),
.Y(n_2048)
);

NOR2x1_ASAP7_75t_L g2049 ( 
.A(n_1991),
.B(n_1971),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_2011),
.A2(n_1919),
.B1(n_1971),
.B2(n_1983),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1987),
.B(n_1942),
.Y(n_2051)
);

INVxp67_ASAP7_75t_SL g2052 ( 
.A(n_2010),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1987),
.B(n_1970),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1985),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1996),
.B(n_1970),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1990),
.Y(n_2056)
);

INVx1_ASAP7_75t_SL g2057 ( 
.A(n_2028),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_2027),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2038),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2038),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2041),
.Y(n_2061)
);

OAI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_2043),
.A2(n_1997),
.B1(n_1991),
.B2(n_2001),
.C(n_1912),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2053),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_2028),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2037),
.B(n_1995),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2034),
.B(n_1999),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2027),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_2051),
.B(n_1996),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_2049),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2034),
.B(n_2005),
.Y(n_2070)
);

OAI21xp33_ASAP7_75t_L g2071 ( 
.A1(n_2043),
.A2(n_2004),
.B(n_1991),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2032),
.A2(n_1991),
.B(n_1997),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2041),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2048),
.A2(n_2031),
.B1(n_2035),
.B2(n_2045),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2030),
.A2(n_1976),
.B1(n_1959),
.B2(n_1919),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2054),
.Y(n_2076)
);

OAI21xp33_ASAP7_75t_L g2077 ( 
.A1(n_2045),
.A2(n_2003),
.B(n_1995),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_2049),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2027),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2057),
.B(n_2037),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2070),
.B(n_2035),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2068),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_2064),
.B(n_2048),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2059),
.B(n_2046),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_2060),
.B(n_2040),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_2070),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2066),
.B(n_2039),
.Y(n_2087)
);

OAI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2074),
.A2(n_2050),
.B1(n_2036),
.B2(n_2046),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2063),
.B(n_2029),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2068),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2063),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2071),
.A2(n_2040),
.B1(n_2052),
.B2(n_2039),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2065),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2066),
.B(n_2029),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2061),
.Y(n_2095)
);

OAI211xp5_ASAP7_75t_SL g2096 ( 
.A1(n_2092),
.A2(n_2078),
.B(n_2069),
.C(n_2062),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_SL g2097 ( 
.A(n_2090),
.B(n_1988),
.Y(n_2097)
);

NOR3xp33_ASAP7_75t_L g2098 ( 
.A(n_2083),
.B(n_2077),
.C(n_2072),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2088),
.A2(n_2075),
.B(n_2058),
.Y(n_2099)
);

AOI221xp5_ASAP7_75t_L g2100 ( 
.A1(n_2085),
.A2(n_2076),
.B1(n_2073),
.B2(n_2058),
.C(n_2067),
.Y(n_2100)
);

OAI221xp5_ASAP7_75t_L g2101 ( 
.A1(n_2092),
.A2(n_2051),
.B1(n_2027),
.B2(n_2067),
.C(n_2079),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_2083),
.A2(n_2079),
.B1(n_2044),
.B2(n_2055),
.C(n_2053),
.Y(n_2102)
);

AOI221x1_ASAP7_75t_L g2103 ( 
.A1(n_2080),
.A2(n_2015),
.B1(n_2009),
.B2(n_2003),
.C(n_2044),
.Y(n_2103)
);

AOI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_2085),
.A2(n_2015),
.B(n_2014),
.Y(n_2104)
);

AOI211xp5_ASAP7_75t_SL g2105 ( 
.A1(n_2084),
.A2(n_2014),
.B(n_2009),
.C(n_2054),
.Y(n_2105)
);

NAND3xp33_ASAP7_75t_L g2106 ( 
.A(n_2090),
.B(n_1976),
.C(n_1959),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2082),
.A2(n_1976),
.B(n_2033),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_2093),
.B(n_2055),
.Y(n_2108)
);

NAND5xp2_ASAP7_75t_L g2109 ( 
.A(n_2081),
.B(n_2033),
.C(n_2047),
.D(n_2042),
.E(n_2056),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_2094),
.A2(n_1976),
.B(n_2056),
.Y(n_2110)
);

NAND3xp33_ASAP7_75t_SL g2111 ( 
.A(n_2089),
.B(n_2091),
.C(n_2087),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2096),
.A2(n_2086),
.B(n_2095),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2102),
.Y(n_2113)
);

XNOR2x1_ASAP7_75t_L g2114 ( 
.A(n_2107),
.B(n_1624),
.Y(n_2114)
);

AOI221xp5_ASAP7_75t_L g2115 ( 
.A1(n_2098),
.A2(n_2101),
.B1(n_2099),
.B2(n_2100),
.C(n_2111),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2104),
.B(n_2105),
.Y(n_2116)
);

OA21x2_ASAP7_75t_SL g2117 ( 
.A1(n_2097),
.A2(n_2005),
.B(n_1976),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2103),
.B(n_2108),
.Y(n_2118)
);

INVxp67_ASAP7_75t_L g2119 ( 
.A(n_2109),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_2106),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2114),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2119),
.B(n_2110),
.Y(n_2122)
);

OAI221xp5_ASAP7_75t_L g2123 ( 
.A1(n_2115),
.A2(n_2118),
.B1(n_2116),
.B2(n_2112),
.C(n_2113),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2120),
.B(n_2042),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2117),
.B(n_2047),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2116),
.B(n_2017),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2119),
.B(n_2005),
.Y(n_2127)
);

OAI21xp5_ASAP7_75t_SL g2128 ( 
.A1(n_2115),
.A2(n_1726),
.B(n_1742),
.Y(n_2128)
);

AOI211xp5_ASAP7_75t_L g2129 ( 
.A1(n_2123),
.A2(n_1726),
.B(n_1742),
.C(n_1988),
.Y(n_2129)
);

XOR2xp5_ASAP7_75t_L g2130 ( 
.A(n_2127),
.B(n_1742),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2125),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2121),
.B(n_2126),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2124),
.Y(n_2133)
);

XNOR2xp5_ASAP7_75t_L g2134 ( 
.A(n_2122),
.B(n_2017),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2128),
.A2(n_2006),
.B(n_1998),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2134),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2131),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2129),
.A2(n_2026),
.B1(n_2024),
.B2(n_2016),
.Y(n_2138)
);

AOI221xp5_ASAP7_75t_L g2139 ( 
.A1(n_2130),
.A2(n_1925),
.B1(n_1939),
.B2(n_1948),
.C(n_1938),
.Y(n_2139)
);

NAND4xp75_ASAP7_75t_L g2140 ( 
.A(n_2137),
.B(n_2132),
.C(n_2133),
.D(n_2135),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2140),
.A2(n_2139),
.B1(n_2129),
.B2(n_2136),
.C(n_2138),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_2141),
.Y(n_2142)
);

OAI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2141),
.A2(n_1948),
.B1(n_2000),
.B2(n_2008),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2142),
.A2(n_2143),
.B1(n_2008),
.B2(n_2000),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2143),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2145),
.A2(n_1989),
.B1(n_1957),
.B2(n_1978),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2144),
.A2(n_1989),
.B1(n_1957),
.B2(n_1978),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2147),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2148),
.B(n_2146),
.Y(n_2149)
);

OR2x6_ASAP7_75t_L g2150 ( 
.A(n_2149),
.B(n_1932),
.Y(n_2150)
);

AOI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_2150),
.A2(n_1989),
.B1(n_1940),
.B2(n_1975),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_SL g2152 ( 
.A1(n_2151),
.A2(n_1925),
.B1(n_1975),
.B2(n_1940),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_2152),
.A2(n_1967),
.B1(n_1938),
.B2(n_1982),
.Y(n_2153)
);


endmodule