module fake_jpeg_22631_n_136 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_1),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_29),
.Y(n_33)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_25),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_20),
.B1(n_21),
.B2(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_19),
.B1(n_26),
.B2(n_23),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_19),
.B1(n_20),
.B2(n_11),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_13),
.C(n_11),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_42),
.C(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_22),
.A2(n_21),
.B1(n_16),
.B2(n_15),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_14),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_R g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_27),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_26),
.B1(n_25),
.B2(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_48),
.B1(n_46),
.B2(n_25),
.Y(n_71)
);

A2O1A1O1Ixp25_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_54),
.B(n_53),
.C(n_42),
.D(n_49),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_27),
.CI(n_24),
.CON(n_77),
.SN(n_77)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_53),
.B(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_76),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_79),
.B1(n_58),
.B2(n_67),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_64),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_36),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_27),
.Y(n_75)
);

NAND2x1_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_63),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_27),
.B(n_24),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_34),
.B1(n_12),
.B2(n_18),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.C(n_75),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_58),
.B1(n_56),
.B2(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_90),
.B1(n_77),
.B2(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_56),
.B1(n_34),
.B2(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_71),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_102),
.C(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_32),
.B1(n_70),
.B2(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_90),
.Y(n_100)
);

BUFx6f_ASAP7_75t_SL g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_18),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_106),
.B(n_18),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_83),
.C(n_88),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_108),
.Y(n_113)
);

XOR2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_99),
.B1(n_97),
.B2(n_96),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_84),
.C(n_32),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_103),
.B1(n_109),
.B2(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_117),
.B(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_8),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_3),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_7),
.B(n_10),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_12),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_12),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_5),
.C(n_6),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_4),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_5),
.B(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_113),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_124),
.B(n_113),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

AOI21x1_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_127),
.B(n_5),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_132),
.B(n_134),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_135),
.Y(n_136)
);


endmodule