module real_jpeg_6184_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_1),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_2),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_91),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_2),
.A2(n_91),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_2),
.A2(n_40),
.B1(n_91),
.B2(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_47),
.B1(n_63),
.B2(n_85),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_47),
.B1(n_137),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_47),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_5),
.A2(n_28),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_7),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_12),
.A2(n_64),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_64),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_12),
.A2(n_64),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_12),
.B(n_75),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_12),
.A2(n_104),
.B(n_260),
.C(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_12),
.B(n_293),
.C(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_12),
.B(n_151),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_12),
.B(n_187),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_12),
.B(n_168),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_13),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_230),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_228),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_197),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_23),
.B(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_140),
.C(n_182),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_24),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_72),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_25),
.B(n_73),
.C(n_100),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_51),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_26),
.B(n_51),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_35),
.B(n_38),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_27),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_37),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_38),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_39),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_39),
.B(n_205),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_39),
.A2(n_205),
.B(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_39),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_41),
.Y(n_209)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_41),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_45),
.B(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_50),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.A3(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_126)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_61),
.A2(n_64),
.B(n_95),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_64),
.A2(n_261),
.B(n_264),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_100),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_88),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_75),
.B(n_89),
.Y(n_155)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_84),
.B(n_93),
.Y(n_225)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_123),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_106),
.Y(n_279)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_108),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_108),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_110),
.Y(n_266)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_116),
.A2(n_124),
.B(n_151),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_116),
.B(n_124),
.Y(n_341)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_122),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_123),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_134),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_128),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_140),
.B(n_182),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_152),
.C(n_156),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_141),
.A2(n_156),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_141),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_150),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_145),
.B(n_151),
.Y(n_241)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_150),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_152),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_155),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_176),
.B(n_177),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_158),
.B(n_278),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_168),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_162),
.B1(n_164),
.B2(n_167),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AO22x2_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_169),
.B1(n_171),
.B2(n_174),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_168),
.B(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_212),
.B(n_219),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_176),
.B(n_177),
.Y(n_276)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_188),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_185),
.B(n_301),
.Y(n_329)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_189),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_190),
.B(n_277),
.Y(n_306)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_220),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_211),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_210),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_202),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_208),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_210),
.B(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_219),
.B(n_297),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_248),
.B(n_353),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_232),
.B(n_246),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_239),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_244),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_316),
.Y(n_327)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_283),
.B(n_352),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_251),
.B(n_254),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_273),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_255),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_258),
.A2(n_273),
.B1(n_274),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_270),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_259),
.A2(n_270),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_346),
.B(n_351),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_334),
.B(n_345),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_310),
.B(n_333),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_298),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_298),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_296),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_289),
.B1(n_296),
.B2(n_313),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.Y(n_298)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_308),
.C(n_336),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_311),
.A2(n_319),
.B(n_332),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_314),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_328),
.B(n_331),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_327),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_337),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_340),
.C(n_342),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_347),
.B(n_350),
.Y(n_351)
);


endmodule