module fake_jpeg_2326_n_287 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_16),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_63),
.B(n_81),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_0),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_2),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NAND2xp67_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_85),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_77),
.Y(n_95)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_80),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_82),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_2),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_25),
.Y(n_92)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_86),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_36),
.B1(n_31),
.B2(n_27),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_92),
.B(n_4),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_36),
.B1(n_31),
.B2(n_27),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_23),
.B(n_35),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_24),
.B1(n_35),
.B2(n_34),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_103),
.B1(n_110),
.B2(n_120),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_29),
.B1(n_34),
.B2(n_33),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_54),
.A2(n_44),
.B1(n_33),
.B2(n_30),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_105),
.B1(n_125),
.B2(n_131),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_44),
.B1(n_24),
.B2(n_30),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_61),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_53),
.B(n_19),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_26),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_41),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_41),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_133),
.B1(n_91),
.B2(n_122),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_41),
.C(n_8),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_41),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_143),
.Y(n_181)
);

AND2x4_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_60),
.Y(n_139)
);

AND2x4_ASAP7_75t_SL g185 ( 
.A(n_139),
.B(n_136),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_151),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_80),
.B1(n_85),
.B2(n_77),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_145),
.B1(n_154),
.B2(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_124),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_14),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_160),
.Y(n_169)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_127),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_109),
.B1(n_91),
.B2(n_122),
.Y(n_154)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_166),
.B1(n_107),
.B2(n_132),
.Y(n_170)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_9),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_106),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_159),
.A2(n_116),
.B1(n_121),
.B2(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_89),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_114),
.A2(n_13),
.B1(n_113),
.B2(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_93),
.B(n_108),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_132),
.B1(n_121),
.B2(n_99),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_173),
.B1(n_179),
.B2(n_155),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_180),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_125),
.B1(n_113),
.B2(n_100),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_126),
.B1(n_100),
.B2(n_129),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_182),
.B1(n_141),
.B2(n_156),
.Y(n_203)
);

AOI22x1_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_126),
.B1(n_107),
.B2(n_127),
.Y(n_179)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_139),
.B(n_116),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_135),
.B1(n_154),
.B2(n_148),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_157),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_142),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_139),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_149),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_180),
.C(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_185),
.B(n_192),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_206),
.B1(n_167),
.B2(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_204),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_213),
.B1(n_214),
.B2(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_207),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_138),
.B1(n_145),
.B2(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_211),
.B(n_212),
.Y(n_225)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_152),
.B(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_205),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_191),
.C(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_220),
.C(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_191),
.C(n_187),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_204),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_193),
.B1(n_201),
.B2(n_197),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_167),
.B(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_229),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_200),
.A2(n_187),
.B1(n_185),
.B2(n_174),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_210),
.B1(n_172),
.B2(n_147),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_234),
.Y(n_257)
);

AOI221xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_209),
.B1(n_185),
.B2(n_212),
.C(n_169),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_183),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_211),
.B(n_195),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_238),
.B(n_221),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_216),
.B1(n_227),
.B2(n_228),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_231),
.B1(n_230),
.B2(n_222),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_172),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_233),
.A2(n_226),
.B1(n_229),
.B2(n_224),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_215),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_254),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_226),
.B1(n_238),
.B2(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_240),
.C(n_226),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_261),
.C(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_243),
.C(n_242),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_250),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_221),
.C(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_218),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_262),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_268),
.B(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_255),
.C(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_255),
.C(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_253),
.C(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_247),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_259),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_258),
.B(n_267),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_265),
.C(n_246),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_281),
.A2(n_274),
.B1(n_276),
.B2(n_278),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_264),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_282),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_246),
.C(n_252),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_218),
.Y(n_287)
);


endmodule