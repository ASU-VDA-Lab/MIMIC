module real_jpeg_8179_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_203;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_63),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_2),
.A2(n_11),
.B(n_52),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_57),
.B1(n_62),
.B2(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_38),
.B(n_42),
.C(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_10),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_11),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_11),
.A2(n_62),
.B1(n_67),
.B2(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_155),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_38),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_38),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_208),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_11),
.A2(n_51),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_51),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_12),
.A2(n_62),
.B1(n_67),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_12),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_128),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_128),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_14),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_15),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_16),
.A2(n_62),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_16),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_16),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_17),
.A2(n_62),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_17),
.A2(n_51),
.B1(n_52),
.B2(n_88),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_88),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_17),
.A2(n_38),
.B1(n_39),
.B2(n_88),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_21),
.B(n_92),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_78),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_47),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_59),
.C(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_36),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_26),
.A2(n_33),
.B(n_34),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_26),
.A2(n_33),
.B1(n_81),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_26),
.A2(n_33),
.B1(n_191),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_26),
.A2(n_33),
.B1(n_193),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_26),
.A2(n_33),
.B1(n_224),
.B2(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_27),
.A2(n_28),
.B1(n_136),
.B2(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_27),
.A2(n_28),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_29),
.B(n_44),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_29),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_30),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_33),
.B(n_132),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_50),
.B2(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_38),
.B(n_55),
.Y(n_236)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_39),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_41),
.A2(n_43),
.B1(n_76),
.B2(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_41),
.A2(n_43),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_41),
.A2(n_43),
.B1(n_199),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_41),
.A2(n_43),
.B1(n_222),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_41),
.A2(n_43),
.B1(n_158),
.B2(n_229),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_42),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_43),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_43),
.B(n_132),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_59),
.B1(n_60),
.B2(n_71),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_54),
.B1(n_58),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_49),
.A2(n_54),
.B1(n_91),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_49),
.A2(n_54),
.B1(n_123),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_49),
.A2(n_54),
.B1(n_151),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_49),
.A2(n_54),
.B1(n_177),
.B2(n_231),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_53),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_54),
.B(n_132),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_65),
.B1(n_69),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_65),
.B1(n_87),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_63),
.B(n_132),
.C(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_72),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_74),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.C(n_89),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_82),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_109),
.B2(n_110),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_100),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_98),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_140),
.B(n_263),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_137),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_115),
.B(n_137),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_119),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_118),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_120),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_124),
.C(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_182),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_164),
.B(n_181),
.Y(n_142)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_161),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_148),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_156),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_150),
.B1(n_156),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_165),
.B(n_167),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_173),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_168),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_171),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_176),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_261),
.C(n_262),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_255),
.B(n_260),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_241),
.B(n_254),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_226),
.B(n_240),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_216),
.B(n_225),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_205),
.B(n_215),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_194),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_204),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_204),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_210),
.B(n_214),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_227),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.CI(n_223),
.CON(n_219),
.SN(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.CI(n_233),
.CON(n_227),
.SN(n_227)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_232),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_243),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_251),
.C(n_252),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_250),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_251),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);


endmodule