module real_aes_8364_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g534 ( .A(n_1), .Y(n_534) );
INVx1_ASAP7_75t_L g155 ( .A(n_2), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_3), .A2(n_38), .B1(n_180), .B2(n_480), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g187 ( .A1(n_4), .A2(n_171), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_5), .B(n_169), .Y(n_546) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_7), .A2(n_258), .B(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_39), .Y(n_114) );
INVx1_ASAP7_75t_L g193 ( .A(n_9), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_10), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g140 ( .A(n_11), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_12), .B(n_161), .Y(n_489) );
INVx1_ASAP7_75t_L g264 ( .A(n_13), .Y(n_264) );
INVx1_ASAP7_75t_L g528 ( .A(n_14), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_15), .B(n_136), .Y(n_517) );
AO32x2_ASAP7_75t_L g501 ( .A1(n_16), .A2(n_135), .A3(n_169), .B1(n_482), .B2(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_17), .B(n_180), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_18), .B(n_176), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_19), .B(n_136), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_20), .A2(n_50), .B1(n_180), .B2(n_480), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_21), .B(n_171), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_22), .A2(n_98), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_22), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_23), .A2(n_76), .B1(n_161), .B2(n_180), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_24), .B(n_180), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_25), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_26), .A2(n_262), .B(n_263), .C(n_265), .Y(n_261) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_27), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_28), .B(n_166), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_29), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_30), .B(n_117), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_31), .A2(n_88), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_31), .Y(n_126) );
INVx1_ASAP7_75t_L g208 ( .A(n_32), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_33), .B(n_166), .Y(n_473) );
INVx2_ASAP7_75t_L g146 ( .A(n_34), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_35), .B(n_180), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_36), .B(n_166), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_37), .A2(n_148), .B(n_151), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g206 ( .A(n_40), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_41), .A2(n_104), .B1(n_115), .B2(n_744), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_42), .B(n_159), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_43), .B(n_180), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_44), .A2(n_86), .B1(n_228), .B2(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_45), .B(n_180), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_46), .B(n_180), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_47), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_48), .B(n_533), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_49), .B(n_171), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_51), .A2(n_61), .B1(n_161), .B2(n_180), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_52), .A2(n_734), .B1(n_735), .B2(n_738), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_52), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_53), .A2(n_151), .B1(n_161), .B2(n_204), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_54), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_55), .B(n_180), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_56), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_57), .B(n_180), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_58), .A2(n_179), .B(n_191), .C(n_192), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_59), .Y(n_241) );
INVx1_ASAP7_75t_L g189 ( .A(n_60), .Y(n_189) );
INVx1_ASAP7_75t_L g149 ( .A(n_62), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_63), .B(n_180), .Y(n_535) );
INVx1_ASAP7_75t_L g139 ( .A(n_64), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_65), .Y(n_445) );
AO32x2_ASAP7_75t_L g477 ( .A1(n_66), .A2(n_169), .A3(n_244), .B1(n_478), .B2(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g553 ( .A(n_67), .Y(n_553) );
INVx1_ASAP7_75t_L g468 ( .A(n_68), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_69), .A2(n_124), .B1(n_440), .B2(n_441), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_69), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_70), .A2(n_176), .B(n_177), .C(n_179), .Y(n_175) );
INVxp67_ASAP7_75t_L g178 ( .A(n_71), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_72), .B(n_161), .Y(n_469) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_74), .Y(n_211) );
INVx1_ASAP7_75t_L g234 ( .A(n_75), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_77), .A2(n_148), .B(n_151), .C(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_78), .B(n_480), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_79), .B(n_161), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_80), .B(n_156), .Y(n_224) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_82), .B(n_176), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_83), .B(n_161), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_84), .A2(n_148), .B(n_151), .C(n_154), .Y(n_150) );
INVx2_ASAP7_75t_L g109 ( .A(n_85), .Y(n_109) );
OR2x2_ASAP7_75t_L g119 ( .A(n_85), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g451 ( .A(n_85), .B(n_121), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_87), .A2(n_102), .B1(n_161), .B2(n_162), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_88), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_89), .B(n_166), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_90), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_91), .A2(n_148), .B(n_151), .C(n_247), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_92), .Y(n_254) );
INVx1_ASAP7_75t_L g174 ( .A(n_93), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_94), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_95), .B(n_156), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_96), .B(n_161), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_97), .B(n_169), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_98), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_100), .A2(n_171), .B(n_172), .Y(n_170) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_101), .A2(n_448), .B1(n_732), .B2(n_733), .C1(n_739), .C2(n_742), .Y(n_447) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_107), .Y(n_745) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
OR2x2_ASAP7_75t_L g455 ( .A(n_109), .B(n_121), .Y(n_455) );
NOR2x2_ASAP7_75t_L g741 ( .A(n_109), .B(n_120), .Y(n_741) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g121 ( .A(n_114), .B(n_122), .Y(n_121) );
AO21x1_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_443), .B(n_446), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_123), .B(n_442), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g441 ( .A(n_124), .Y(n_441) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
INVx1_ASAP7_75t_L g452 ( .A(n_128), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_128), .A2(n_453), .B1(n_457), .B2(n_743), .Y(n_742) );
NAND2x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_356), .Y(n_128) );
NOR5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_279), .C(n_311), .D(n_326), .E(n_343), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_195), .B(n_216), .C(n_267), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_167), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_132), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_132), .B(n_331), .Y(n_394) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_133), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_133), .B(n_213), .Y(n_280) );
AND2x2_ASAP7_75t_L g321 ( .A(n_133), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_133), .B(n_290), .Y(n_325) );
OR2x2_ASAP7_75t_L g362 ( .A(n_133), .B(n_201), .Y(n_362) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g200 ( .A(n_134), .B(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g270 ( .A(n_134), .Y(n_270) );
OR2x2_ASAP7_75t_L g433 ( .A(n_134), .B(n_273), .Y(n_433) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_141), .B(n_163), .Y(n_134) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_135), .A2(n_202), .B(n_210), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_135), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g229 ( .A(n_135), .Y(n_229) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_137), .B(n_138), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_150), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_143), .A2(n_181), .B1(n_203), .B2(n_209), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_143), .A2(n_234), .B(n_235), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
AND2x4_ASAP7_75t_L g171 ( .A(n_144), .B(n_148), .Y(n_171) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g533 ( .A(n_145), .Y(n_533) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx3_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_147), .Y(n_159) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
INVx4_ASAP7_75t_SL g181 ( .A(n_148), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_148), .A2(n_467), .B(n_470), .Y(n_466) );
BUFx3_ASAP7_75t_L g482 ( .A(n_148), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_148), .A2(n_487), .B(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_148), .A2(n_527), .B(n_531), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_148), .A2(n_540), .B(n_543), .Y(n_539) );
INVx5_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
BUFx3_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
INVx1_ASAP7_75t_L g480 ( .A(n_152), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_158), .C(n_160), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_SL g467 ( .A1(n_156), .A2(n_179), .B(n_468), .C(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g504 ( .A(n_156), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_156), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_156), .A2(n_550), .B(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_157), .B(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_157), .B(n_193), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g478 ( .A1(n_157), .A2(n_159), .B1(n_479), .B2(n_481), .Y(n_478) );
INVx2_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVx4_ASAP7_75t_L g250 ( .A(n_159), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_159), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_159), .A2(n_504), .B1(n_520), .B2(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_160), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_165), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_165), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g244 ( .A(n_166), .Y(n_244) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_166), .A2(n_257), .B(n_266), .Y(n_256) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_166), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_166), .A2(n_486), .B(n_494), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_167), .A2(n_336), .B1(n_337), .B2(n_340), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_167), .B(n_270), .Y(n_419) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_185), .Y(n_167) );
AND2x2_ASAP7_75t_L g215 ( .A(n_168), .B(n_201), .Y(n_215) );
AND2x2_ASAP7_75t_L g272 ( .A(n_168), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g277 ( .A(n_168), .Y(n_277) );
INVx3_ASAP7_75t_L g290 ( .A(n_168), .Y(n_290) );
OR2x2_ASAP7_75t_L g310 ( .A(n_168), .B(n_273), .Y(n_310) );
AND2x2_ASAP7_75t_L g329 ( .A(n_168), .B(n_186), .Y(n_329) );
BUFx2_ASAP7_75t_L g361 ( .A(n_168), .Y(n_361) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_182), .Y(n_168) );
INVx4_ASAP7_75t_L g184 ( .A(n_169), .Y(n_184) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_169), .A2(n_539), .B(n_546), .Y(n_538) );
BUFx2_ASAP7_75t_L g258 ( .A(n_171), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_181), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_181), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_173), .A2(n_181), .B(n_260), .C(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g490 ( .A(n_176), .Y(n_490) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_180), .Y(n_251) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_183), .A2(n_187), .B(n_194), .Y(n_186) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_184), .B(n_231), .Y(n_230) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_184), .B(n_482), .C(n_519), .Y(n_518) );
AO21x1_ASAP7_75t_L g608 ( .A1(n_184), .A2(n_519), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g276 ( .A(n_185), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
BUFx2_ASAP7_75t_L g199 ( .A(n_186), .Y(n_199) );
INVx2_ASAP7_75t_L g214 ( .A(n_186), .Y(n_214) );
OR2x2_ASAP7_75t_L g292 ( .A(n_186), .B(n_273), .Y(n_292) );
AND2x2_ASAP7_75t_L g322 ( .A(n_186), .B(n_201), .Y(n_322) );
AND2x2_ASAP7_75t_L g339 ( .A(n_186), .B(n_270), .Y(n_339) );
AND2x2_ASAP7_75t_L g379 ( .A(n_186), .B(n_290), .Y(n_379) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_186), .B(n_215), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_191), .A2(n_492), .B(n_493), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g552 ( .A1(n_191), .A2(n_532), .B(n_553), .C(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp33_ASAP7_75t_SL g196 ( .A(n_197), .B(n_212), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_198), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_199), .A2(n_215), .B(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_199), .B(n_201), .Y(n_409) );
AND2x2_ASAP7_75t_L g345 ( .A(n_200), .B(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_201), .Y(n_371) );
OAI22xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_204) );
INVx2_ASAP7_75t_L g207 ( .A(n_205), .Y(n_207) );
INVx4_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_212), .B(n_270), .Y(n_438) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_213), .A2(n_381), .B1(n_382), .B2(n_387), .Y(n_380) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x2_ASAP7_75t_L g271 ( .A(n_214), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g309 ( .A(n_214), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g346 ( .A(n_214), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_215), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g400 ( .A(n_215), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_242), .Y(n_217) );
INVx4_ASAP7_75t_L g286 ( .A(n_218), .Y(n_286) );
AND2x2_ASAP7_75t_L g364 ( .A(n_218), .B(n_331), .Y(n_364) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_232), .Y(n_218) );
INVx3_ASAP7_75t_L g283 ( .A(n_219), .Y(n_283) );
AND2x2_ASAP7_75t_L g297 ( .A(n_219), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g301 ( .A(n_219), .Y(n_301) );
INVx2_ASAP7_75t_L g315 ( .A(n_219), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_219), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g372 ( .A(n_219), .B(n_367), .Y(n_372) );
AND2x2_ASAP7_75t_L g437 ( .A(n_219), .B(n_407), .Y(n_437) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_230), .Y(n_219) );
AOI21xp5_ASAP7_75t_SL g220 ( .A1(n_221), .A2(n_222), .B(n_229), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_226), .A2(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
INVx1_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_229), .A2(n_526), .B(n_536), .Y(n_525) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_229), .A2(n_548), .B(n_555), .Y(n_547) );
AND2x2_ASAP7_75t_L g278 ( .A(n_232), .B(n_256), .Y(n_278) );
INVx2_ASAP7_75t_L g298 ( .A(n_232), .Y(n_298) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_239), .B(n_240), .Y(n_232) );
INVx1_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
AND2x2_ASAP7_75t_L g349 ( .A(n_242), .B(n_297), .Y(n_349) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_255), .Y(n_242) );
INVx2_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
INVx1_ASAP7_75t_L g296 ( .A(n_243), .Y(n_296) );
AND2x2_ASAP7_75t_L g314 ( .A(n_243), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_243), .B(n_298), .Y(n_352) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_253), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_252), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_251), .Y(n_247) );
AND2x2_ASAP7_75t_L g331 ( .A(n_255), .B(n_288), .Y(n_331) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
AND2x2_ASAP7_75t_L g367 ( .A(n_256), .B(n_298), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_262), .B(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_262), .A2(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g530 ( .A(n_262), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_274), .B(n_278), .Y(n_267) );
INVx1_ASAP7_75t_SL g312 ( .A(n_268), .Y(n_312) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_269), .B(n_276), .Y(n_369) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g318 ( .A(n_270), .B(n_273), .Y(n_318) );
AND2x2_ASAP7_75t_L g347 ( .A(n_270), .B(n_291), .Y(n_347) );
OR2x2_ASAP7_75t_L g350 ( .A(n_270), .B(n_310), .Y(n_350) );
AOI222xp33_ASAP7_75t_L g414 ( .A1(n_271), .A2(n_363), .B1(n_415), .B2(n_416), .C1(n_418), .C2(n_420), .Y(n_414) );
BUFx2_ASAP7_75t_L g328 ( .A(n_273), .Y(n_328) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g317 ( .A(n_276), .B(n_318), .Y(n_317) );
INVx3_ASAP7_75t_SL g334 ( .A(n_276), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_276), .B(n_328), .Y(n_388) );
AND2x2_ASAP7_75t_L g323 ( .A(n_278), .B(n_283), .Y(n_323) );
INVx1_ASAP7_75t_L g342 ( .A(n_278), .Y(n_342) );
OAI221xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_281), .B1(n_285), .B2(n_289), .C(n_293), .Y(n_279) );
OR2x2_ASAP7_75t_L g351 ( .A(n_281), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x2_ASAP7_75t_L g336 ( .A(n_283), .B(n_306), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_283), .B(n_296), .Y(n_376) );
AND2x2_ASAP7_75t_L g381 ( .A(n_283), .B(n_331), .Y(n_381) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_283), .Y(n_391) );
NAND2x1_ASAP7_75t_SL g402 ( .A(n_283), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g287 ( .A(n_284), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_284), .B(n_302), .Y(n_333) );
INVx1_ASAP7_75t_L g399 ( .A(n_284), .Y(n_399) );
INVx1_ASAP7_75t_L g374 ( .A(n_285), .Y(n_374) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g386 ( .A(n_286), .Y(n_386) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_286), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g403 ( .A(n_287), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_287), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g306 ( .A(n_288), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_288), .B(n_298), .Y(n_319) );
INVx1_ASAP7_75t_L g385 ( .A(n_288), .Y(n_385) );
INVx1_ASAP7_75t_L g406 ( .A(n_289), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI21xp5_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_299), .B(n_308), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x2_ASAP7_75t_L g439 ( .A(n_295), .B(n_372), .Y(n_439) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g407 ( .A(n_296), .B(n_367), .Y(n_407) );
AOI32xp33_ASAP7_75t_L g320 ( .A1(n_297), .A2(n_303), .A3(n_321), .B1(n_323), .B2(n_324), .Y(n_320) );
AOI322xp5_ASAP7_75t_L g422 ( .A1(n_297), .A2(n_329), .A3(n_412), .B1(n_423), .B2(n_424), .C1(n_425), .C2(n_427), .Y(n_422) );
INVx2_ASAP7_75t_L g302 ( .A(n_298), .Y(n_302) );
INVx1_ASAP7_75t_L g412 ( .A(n_298), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B1(n_304), .B2(n_305), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_300), .B(n_306), .Y(n_355) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_301), .B(n_367), .Y(n_417) );
INVx1_ASAP7_75t_L g304 ( .A(n_302), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_302), .B(n_331), .Y(n_421) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_310), .B(n_405), .Y(n_404) );
OAI221xp5_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_313), .B1(n_316), .B2(n_319), .C(n_320), .Y(n_311) );
OR2x2_ASAP7_75t_L g332 ( .A(n_313), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g341 ( .A(n_313), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g366 ( .A(n_314), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g370 ( .A(n_324), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_332), .B2(n_334), .C(n_335), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_328), .A2(n_359), .B1(n_363), .B2(n_364), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_329), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_329), .Y(n_434) );
INVx1_ASAP7_75t_L g428 ( .A(n_331), .Y(n_428) );
INVx1_ASAP7_75t_SL g363 ( .A(n_332), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_334), .B(n_362), .Y(n_424) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_339), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g405 ( .A(n_339), .Y(n_405) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
OAI221xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_348), .B1(n_350), .B2(n_351), .C(n_353), .Y(n_343) );
NOR2xp33_ASAP7_75t_SL g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_345), .A2(n_363), .B1(n_409), .B2(n_410), .Y(n_408) );
CKINVDCx14_ASAP7_75t_R g348 ( .A(n_349), .Y(n_348) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_350), .A2(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR3xp33_ASAP7_75t_SL g356 ( .A(n_357), .B(n_389), .C(n_413), .Y(n_356) );
NAND4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_365), .C(n_373), .D(n_380), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g436 ( .A(n_361), .Y(n_436) );
INVx3_ASAP7_75t_SL g430 ( .A(n_362), .Y(n_430) );
OR2x2_ASAP7_75t_L g435 ( .A(n_362), .B(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_370), .B2(n_372), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_367), .B(n_385), .Y(n_426) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B(n_377), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_392), .B(n_395), .C(n_408), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_400), .B1(n_401), .B2(n_404), .C1(n_406), .C2(n_407), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND4xp25_ASAP7_75t_SL g432 ( .A(n_405), .B(n_433), .C(n_434), .D(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND3xp33_ASAP7_75t_SL g413 ( .A(n_414), .B(n_422), .C(n_431), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_437), .B1(n_438), .B2(n_439), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_442), .A2(n_443), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B1(n_453), .B2(n_456), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g743 ( .A(n_450), .Y(n_743) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_653), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_602), .C(n_644), .Y(n_458) );
AOI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_511), .B(n_556), .C(n_578), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_474), .B(n_495), .C(n_506), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_462), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g665 ( .A(n_462), .B(n_582), .Y(n_665) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g567 ( .A(n_463), .B(n_498), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_463), .B(n_485), .Y(n_684) );
INVx1_ASAP7_75t_L g702 ( .A(n_463), .Y(n_702) );
AND2x2_ASAP7_75t_L g711 ( .A(n_463), .B(n_599), .Y(n_711) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g594 ( .A(n_464), .B(n_485), .Y(n_594) );
AND2x2_ASAP7_75t_L g652 ( .A(n_464), .B(n_599), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_464), .Y(n_696) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g573 ( .A(n_465), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g581 ( .A(n_465), .Y(n_581) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_465), .Y(n_621) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
AND2x2_ASAP7_75t_L g560 ( .A(n_476), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g593 ( .A(n_476), .Y(n_593) );
OR2x2_ASAP7_75t_L g719 ( .A(n_476), .B(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_476), .B(n_485), .Y(n_723) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx1_ASAP7_75t_L g509 ( .A(n_477), .Y(n_509) );
AND2x2_ASAP7_75t_L g582 ( .A(n_477), .B(n_500), .Y(n_582) );
AND2x2_ASAP7_75t_L g622 ( .A(n_477), .B(n_501), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_482), .A2(n_549), .B(n_552), .Y(n_548) );
INVxp67_ASAP7_75t_L g664 ( .A(n_483), .Y(n_664) );
AND2x4_ASAP7_75t_L g689 ( .A(n_483), .B(n_582), .Y(n_689) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_484), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g499 ( .A(n_485), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g568 ( .A(n_485), .B(n_501), .Y(n_568) );
INVx1_ASAP7_75t_L g574 ( .A(n_485), .Y(n_574) );
INVx2_ASAP7_75t_L g600 ( .A(n_485), .Y(n_600) );
AND2x2_ASAP7_75t_L g616 ( .A(n_485), .B(n_617), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_496), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
AND2x2_ASAP7_75t_L g679 ( .A(n_498), .B(n_500), .Y(n_679) );
AND2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_581), .Y(n_596) );
AND2x2_ASAP7_75t_L g695 ( .A(n_499), .B(n_696), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_500), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g720 ( .A(n_500), .B(n_581), .Y(n_720) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g510 ( .A(n_501), .Y(n_510) );
AND2x2_ASAP7_75t_L g599 ( .A(n_501), .B(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_504), .A2(n_532), .B(n_534), .C(n_535), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_504), .A2(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AND2x2_ASAP7_75t_L g645 ( .A(n_508), .B(n_580), .Y(n_645) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_509), .B(n_581), .Y(n_630) );
INVx2_ASAP7_75t_L g629 ( .A(n_510), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_510), .A2(n_573), .B1(n_634), .B2(n_636), .C1(n_637), .C2(n_640), .Y(n_633) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g558 ( .A(n_515), .Y(n_558) );
OR2x2_ASAP7_75t_L g669 ( .A(n_515), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_516), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g648 ( .A(n_516), .B(n_562), .Y(n_648) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_522), .A2(n_612), .B1(n_651), .B2(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_537), .Y(n_522) );
INVx3_ASAP7_75t_L g584 ( .A(n_523), .Y(n_584) );
OR2x2_ASAP7_75t_L g717 ( .A(n_523), .B(n_593), .Y(n_717) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g590 ( .A(n_524), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g606 ( .A(n_524), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g614 ( .A(n_524), .B(n_562), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_524), .B(n_538), .Y(n_670) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g561 ( .A(n_525), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g565 ( .A(n_525), .B(n_538), .Y(n_565) );
AND2x2_ASAP7_75t_L g641 ( .A(n_525), .B(n_588), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_525), .B(n_547), .Y(n_681) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_537), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_558), .Y(n_597) );
AND2x2_ASAP7_75t_L g601 ( .A(n_537), .B(n_591), .Y(n_601) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
INVx3_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
AND2x2_ASAP7_75t_L g587 ( .A(n_538), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g722 ( .A(n_538), .B(n_705), .Y(n_722) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_547), .Y(n_576) );
INVx2_ASAP7_75t_L g588 ( .A(n_547), .Y(n_588) );
AND2x2_ASAP7_75t_L g632 ( .A(n_547), .B(n_608), .Y(n_632) );
INVx1_ASAP7_75t_L g675 ( .A(n_547), .Y(n_675) );
OR2x2_ASAP7_75t_L g706 ( .A(n_547), .B(n_608), .Y(n_706) );
AND2x2_ASAP7_75t_L g726 ( .A(n_547), .B(n_562), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g564 ( .A(n_558), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_558), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g683 ( .A(n_560), .Y(n_683) );
INVx2_ASAP7_75t_SL g577 ( .A(n_561), .Y(n_577) );
AND2x2_ASAP7_75t_L g697 ( .A(n_561), .B(n_591), .Y(n_697) );
INVx2_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_562), .B(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_569), .B2(n_575), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_565), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g731 ( .A(n_565), .Y(n_731) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g656 ( .A(n_567), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_567), .B(n_599), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_568), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_568), .B(n_621), .Y(n_672) );
INVx2_ASAP7_75t_L g728 ( .A(n_568), .Y(n_728) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_571), .B(n_616), .Y(n_649) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_573), .B(n_593), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g710 ( .A(n_576), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_577), .A2(n_661), .B(n_663), .C(n_666), .Y(n_660) );
OR2x2_ASAP7_75t_L g687 ( .A(n_577), .B(n_591), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_583), .B1(n_585), .B2(n_592), .C(n_595), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_580), .B(n_629), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_580), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g714 ( .A(n_580), .Y(n_714) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_581), .Y(n_605) );
INVx1_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_584), .B(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g692 ( .A(n_584), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_584), .B(n_632), .Y(n_708) );
INVx2_ASAP7_75t_L g694 ( .A(n_585), .Y(n_694) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g635 ( .A(n_587), .B(n_606), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_587), .A2(n_603), .B(n_645), .C(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g613 ( .A(n_588), .B(n_608), .Y(n_613) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_592), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g661 ( .A(n_593), .B(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_598), .B2(n_601), .Y(n_595) );
INVx1_ASAP7_75t_L g715 ( .A(n_597), .Y(n_715) );
INVx1_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
AOI211xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_606), .B(n_610), .C(n_633), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g625 ( .A(n_605), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g676 ( .A(n_606), .Y(n_676) );
AND2x2_ASAP7_75t_L g725 ( .A(n_606), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_615), .B(n_623), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx2_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_613), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g631 ( .A(n_614), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g707 ( .A(n_614), .Y(n_707) );
OAI32xp33_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_666), .A3(n_673), .B1(n_714), .B2(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_SL g686 ( .A(n_616), .Y(n_686) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g626 ( .A(n_622), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_631), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_625), .A2(n_673), .B1(n_699), .B2(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_629), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g666 ( .A(n_632), .Y(n_666) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_652), .A2(n_694), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g653 ( .A(n_654), .B(n_677), .C(n_693), .D(n_703), .E(n_721), .Y(n_653) );
AOI211xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_667), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g724 ( .A(n_661), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_SL g700 ( .A(n_670), .Y(n_700) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_673), .A2(n_683), .A3(n_684), .B1(n_685), .B2(n_686), .C1(n_687), .C2(n_688), .Y(n_682) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g685 ( .A(n_675), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_675), .B(n_700), .Y(n_699) );
AOI211xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_680), .B(n_682), .C(n_690), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_686), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g729 ( .A(n_696), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_711), .B1(n_712), .B2(n_716), .C(n_718), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_708), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g730 ( .A(n_706), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .C(n_727), .Y(n_721) );
AOI21xp33_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_729), .B(n_730), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
endmodule