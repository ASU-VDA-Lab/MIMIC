module fake_jpeg_1478_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_36),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_45),
.B1(n_48),
.B2(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_48),
.B1(n_47),
.B2(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_63),
.B1(n_38),
.B2(n_2),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_0),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_46),
.B1(n_40),
.B2(n_39),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_45),
.B1(n_38),
.B2(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_56),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_52),
.B1(n_51),
.B2(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_1),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_71),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_31),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_43),
.B1(n_37),
.B2(n_39),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_43),
.B1(n_37),
.B2(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_34),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_38),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_84),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_65),
.B1(n_66),
.B2(n_64),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_74),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_66),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_100),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_85),
.B(n_92),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_17),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_104),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_5),
.CI(n_7),
.CON(n_98),
.SN(n_98)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_7),
.B(n_8),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_19),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_107),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_108),
.Y(n_113)
);

XOR2x2_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_18),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_11),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_20),
.C(n_29),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_110),
.B(n_98),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_22),
.B(n_26),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_102),
.C(n_121),
.Y(n_124)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_12),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_13),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_107),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_97),
.C(n_23),
.Y(n_128)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_130),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_123),
.B(n_115),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_123),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.C(n_125),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_113),
.B(n_131),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_109),
.A3(n_111),
.B1(n_132),
.B2(n_112),
.C1(n_115),
.C2(n_24),
.Y(n_142)
);

NAND4xp25_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_30),
.C(n_14),
.D(n_15),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_13),
.Y(n_144)
);


endmodule