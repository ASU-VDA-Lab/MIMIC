module fake_netlist_6_2812_n_1867 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1867);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1867;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_50),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_17),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_81),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_29),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_90),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_25),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_48),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_49),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_70),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_68),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_77),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_61),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_2),
.Y(n_206)
);

BUFx2_ASAP7_75t_SL g207 ( 
.A(n_170),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_113),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_26),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_107),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_86),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_9),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_35),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_83),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_43),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_63),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_97),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_85),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_32),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_67),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_54),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_34),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_42),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_100),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_84),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_37),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_59),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_123),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_110),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_10),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_19),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_93),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_50),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_141),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_151),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_72),
.Y(n_253)
);

BUFx2_ASAP7_75t_SL g254 ( 
.A(n_124),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_16),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_87),
.Y(n_257)
);

BUFx8_ASAP7_75t_SL g258 ( 
.A(n_92),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_66),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_89),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_75),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_133),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_46),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_179),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_94),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_169),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_153),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_147),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_31),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_135),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_31),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_162),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_38),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_55),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_15),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_36),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_99),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_62),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_80),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_114),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_35),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_171),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_12),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_173),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_52),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_6),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_28),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_180),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_160),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_55),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_166),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_109),
.Y(n_301)
);

BUFx8_ASAP7_75t_SL g302 ( 
.A(n_36),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_60),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_43),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_150),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_134),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_131),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_5),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_74),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_14),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_49),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_148),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_126),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_125),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_167),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_79),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_139),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_105),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_33),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_33),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_46),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_24),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_27),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_45),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_25),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_32),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_175),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_57),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_118),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_120),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_156),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_95),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_24),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_16),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_42),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_143),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_78),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_64),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_22),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_117),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_98),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_129),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_149),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_65),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_56),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_18),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_103),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_76),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_41),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_54),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_168),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_62),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_106),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_71),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_2),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_17),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_91),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_206),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_302),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_206),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_305),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_185),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_3),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_193),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_230),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_221),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_200),
.B(n_321),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_230),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_239),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_237),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_230),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_230),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_220),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_200),
.B(n_321),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_200),
.B(n_4),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_181),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_225),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_215),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_217),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_230),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_228),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_272),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_R g392 ( 
.A(n_347),
.B(n_128),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_197),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_181),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_240),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_243),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_248),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_364),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_258),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_186),
.B(n_6),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_218),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_249),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_216),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_219),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_223),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_224),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_204),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_226),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_256),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_204),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_259),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_233),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_265),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_245),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_283),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_225),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_283),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_286),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_288),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_273),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_231),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_293),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_232),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_298),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_275),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_235),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_310),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_183),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_234),
.B(n_7),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_227),
.B(n_8),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_241),
.B(n_8),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_276),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_253),
.B(n_10),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_278),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_280),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_282),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_184),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_236),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_188),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_262),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_326),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_242),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_195),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_289),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_292),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_183),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_203),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_205),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_295),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_212),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_326),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_326),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_214),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_262),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_399),
.B(n_401),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_373),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_421),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_377),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_385),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_423),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_383),
.B(n_410),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_229),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_246),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_447),
.Y(n_485)
);

AND2x6_ASAP7_75t_L g486 ( 
.A(n_375),
.B(n_225),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_416),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_416),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_426),
.Y(n_491)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_416),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_416),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_370),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_415),
.B(n_279),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_404),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_372),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_444),
.Y(n_501)
);

BUFx8_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_378),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_386),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_382),
.B(n_371),
.C(n_388),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_448),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_367),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_367),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_414),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_386),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_410),
.B(n_255),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_449),
.B(n_269),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_422),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_387),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_387),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_390),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_458),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_390),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_453),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_456),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_437),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_395),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_439),
.A2(n_297),
.B(n_291),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_440),
.A2(n_311),
.B(n_304),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_395),
.Y(n_538)
);

BUFx8_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_506),
.B(n_484),
.C(n_397),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_535),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_384),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_535),
.B(n_384),
.Y(n_544)
);

INVx4_ASAP7_75t_SL g545 ( 
.A(n_486),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_471),
.B(n_396),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_530),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_487),
.B(n_381),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_532),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_497),
.B(n_396),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_486),
.B(n_225),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_471),
.B(n_225),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_535),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_532),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_495),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_471),
.B(n_397),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_497),
.A2(n_400),
.B1(n_431),
.B2(n_432),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_R g562 ( 
.A1(n_504),
.A2(n_222),
.B1(n_294),
.B2(n_277),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_485),
.B(n_452),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_495),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_494),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_512),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_472),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_496),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_462),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_471),
.B(n_402),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_482),
.B(n_402),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_486),
.B(n_238),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_482),
.B(n_409),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_472),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_482),
.B(n_238),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_513),
.B(n_394),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_472),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_482),
.B(n_409),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_463),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_499),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_516),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_516),
.B(n_411),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_516),
.B(n_238),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_520),
.B(n_411),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_509),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_516),
.B(n_413),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_522),
.A2(n_434),
.B1(n_394),
.B2(n_430),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_485),
.B(n_413),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_513),
.B(n_420),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_463),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_515),
.B(n_425),
.C(n_420),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_521),
.A2(n_438),
.B1(n_455),
.B2(n_451),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_533),
.B(n_441),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_533),
.B(n_425),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_512),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_467),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_486),
.B(n_433),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_496),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_498),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_465),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_433),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_526),
.B(n_438),
.C(n_435),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_498),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_534),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_486),
.B(n_435),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_500),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_500),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_476),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_513),
.B(n_442),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_486),
.B(n_442),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_468),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_512),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_505),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_488),
.B(n_489),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_505),
.B(n_238),
.Y(n_624)
);

BUFx10_ASAP7_75t_L g625 ( 
.A(n_538),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_529),
.B(n_450),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_512),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_510),
.B(n_417),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_510),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_512),
.B(n_450),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_476),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_473),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_480),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_474),
.B(n_451),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

INVx4_ASAP7_75t_SL g637 ( 
.A(n_492),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_488),
.B(n_455),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_475),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_511),
.B(n_366),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_536),
.A2(n_271),
.B1(n_279),
.B2(n_244),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_511),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_514),
.A2(n_369),
.B1(n_300),
.B2(n_303),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_480),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_475),
.B(n_457),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_492),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_518),
.Y(n_649)
);

BUFx4f_ASAP7_75t_L g650 ( 
.A(n_536),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_493),
.B(n_247),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_529),
.B(n_238),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_483),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_503),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_476),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_523),
.B(n_368),
.Y(n_656)
);

INVx8_ASAP7_75t_L g657 ( 
.A(n_464),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_518),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_519),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_519),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_480),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_490),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_502),
.B(n_313),
.C(n_309),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_469),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_492),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_531),
.B(n_182),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_524),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_493),
.B(n_251),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_525),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_525),
.A2(n_209),
.B1(n_365),
.B2(n_190),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_490),
.B(n_252),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_466),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_490),
.B(n_257),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_490),
.B(n_260),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_492),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_527),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_470),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_527),
.B(n_322),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_531),
.B(n_392),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_469),
.B(n_261),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_536),
.A2(n_271),
.B1(n_250),
.B2(n_244),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_528),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_528),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_523),
.B(n_391),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_477),
.B(n_263),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_478),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_539),
.A2(n_398),
.B1(n_213),
.B2(n_208),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_536),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_656),
.B(n_491),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_628),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_554),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_657),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_684),
.B(n_537),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_546),
.B(n_501),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_543),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_558),
.B(n_244),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_684),
.B(n_537),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_558),
.B(n_244),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_565),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_591),
.B(n_537),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_591),
.B(n_537),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_628),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_607),
.B(n_332),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_607),
.B(n_342),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_548),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_541),
.B(n_478),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_593),
.B(n_507),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_558),
.B(n_650),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_550),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_542),
.A2(n_582),
.B1(n_560),
.B2(n_682),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_600),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_551),
.B(n_461),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_556),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_542),
.B(n_182),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_650),
.A2(n_479),
.B(n_481),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_617),
.B(n_346),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_617),
.A2(n_307),
.B1(n_308),
.B2(n_306),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_540),
.B(n_187),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_576),
.A2(n_354),
.B(n_355),
.C(n_360),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_609),
.B(n_589),
.C(n_586),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_582),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_680),
.B(n_479),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_657),
.B(n_207),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_558),
.B(n_244),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_565),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_557),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_576),
.A2(n_481),
.B(n_209),
.C(n_365),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_646),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_547),
.B(n_187),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_641),
.A2(n_312),
.B1(n_356),
.B2(n_198),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_564),
.Y(n_732)
);

BUFx5_ASAP7_75t_L g733 ( 
.A(n_689),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_554),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_568),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_604),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_682),
.B(n_250),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_603),
.B(n_250),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_569),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_630),
.B(n_264),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_630),
.B(n_266),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_660),
.B(n_267),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_648),
.Y(n_743)
);

INVx5_ASAP7_75t_L g744 ( 
.A(n_561),
.Y(n_744)
);

OAI221xp5_ASAP7_75t_L g745 ( 
.A1(n_660),
.A2(n_325),
.B1(n_328),
.B2(n_329),
.C(n_330),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_569),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_563),
.B(n_189),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_626),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_559),
.B(n_191),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_638),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_579),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_612),
.B(n_250),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_605),
.B(n_268),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_571),
.A2(n_331),
.B1(n_333),
.B2(n_324),
.C(n_323),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_641),
.A2(n_250),
.B1(n_210),
.B2(n_345),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_619),
.B(n_210),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_610),
.B(n_270),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_613),
.B(n_274),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_570),
.B(n_191),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_579),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_614),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_622),
.B(n_281),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_689),
.A2(n_210),
.B1(n_345),
.B2(n_254),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_629),
.B(n_284),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_646),
.B(n_320),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_642),
.B(n_287),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_290),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_649),
.B(n_296),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_671),
.A2(n_345),
.B1(n_210),
.B2(n_194),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_592),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_658),
.B(n_659),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_635),
.B(n_192),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_549),
.B(n_189),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_635),
.B(n_192),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_668),
.B(n_670),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_573),
.B(n_199),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_677),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_648),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_683),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_666),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_687),
.B(n_299),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_578),
.B(n_199),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_544),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_687),
.B(n_301),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_595),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_602),
.B(n_190),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_545),
.B(n_210),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_584),
.B(n_588),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_544),
.B(n_201),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_599),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_599),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_545),
.B(n_210),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_686),
.B(n_201),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_597),
.B(n_314),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_555),
.A2(n_334),
.B1(n_319),
.B2(n_318),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_595),
.B(n_315),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_553),
.A2(n_208),
.B1(n_213),
.B2(n_361),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_657),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_653),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_667),
.B(n_336),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_545),
.B(n_210),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_606),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_618),
.B(n_210),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_618),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_632),
.B(n_316),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_620),
.B(n_194),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_632),
.B(n_634),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_634),
.B(n_317),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_667),
.B(n_539),
.C(n_502),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_640),
.B(n_196),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_639),
.B(n_345),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_633),
.B(n_337),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_633),
.B(n_337),
.Y(n_813)
);

AND2x6_ASAP7_75t_SL g814 ( 
.A(n_685),
.B(n_196),
.Y(n_814)
);

AND2x6_ASAP7_75t_SL g815 ( 
.A(n_562),
.B(n_202),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_666),
.B(n_345),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_671),
.B(n_343),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_666),
.B(n_345),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_581),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_645),
.B(n_343),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_640),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_645),
.B(n_348),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_647),
.B(n_348),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_653),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_681),
.B(n_345),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_202),
.C(n_211),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_640),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_552),
.A2(n_345),
.B1(n_351),
.B2(n_359),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_651),
.B(n_350),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_679),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_666),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_664),
.Y(n_832)
);

BUFx4f_ASAP7_75t_L g833 ( 
.A(n_590),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_669),
.B(n_350),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_553),
.B(n_349),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_679),
.A2(n_361),
.B1(n_539),
.B2(n_285),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_676),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_664),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_643),
.B(n_344),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_654),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_665),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_679),
.B(n_672),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_L g843 ( 
.A1(n_575),
.A2(n_285),
.B(n_539),
.C(n_357),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_596),
.B(n_285),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_676),
.Y(n_845)
);

AND2x2_ASAP7_75t_SL g846 ( 
.A(n_552),
.B(n_82),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_674),
.A2(n_359),
.B1(n_357),
.B2(n_353),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_675),
.B(n_353),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_575),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_662),
.B(n_352),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_662),
.B(n_352),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_665),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_611),
.B(n_351),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_694),
.A2(n_572),
.B(n_623),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_698),
.A2(n_572),
.B(n_585),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_807),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_729),
.B(n_765),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_712),
.B(n_611),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_819),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_701),
.A2(n_585),
.B(n_601),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_702),
.A2(n_601),
.B(n_566),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_788),
.B(n_615),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_716),
.A2(n_763),
.B(n_752),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_783),
.B(n_611),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_788),
.B(n_615),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_738),
.A2(n_621),
.B(n_627),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_715),
.A2(n_688),
.B(n_621),
.C(n_627),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_715),
.B(n_567),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_723),
.A2(n_566),
.B(n_661),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_772),
.A2(n_631),
.B(n_636),
.C(n_655),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_842),
.A2(n_661),
.B(n_636),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_842),
.A2(n_661),
.B(n_631),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_763),
.A2(n_655),
.B(n_661),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_561),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_800),
.B(n_561),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_738),
.A2(n_652),
.B(n_624),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_728),
.A2(n_652),
.B(n_338),
.C(n_339),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_778),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_790),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_791),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_778),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_722),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_709),
.A2(n_594),
.B(n_580),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_800),
.B(n_561),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_772),
.B(n_574),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_774),
.B(n_625),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_750),
.B(n_625),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_721),
.A2(n_625),
.B1(n_587),
.B2(n_583),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_693),
.B(n_673),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_774),
.B(n_574),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_799),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_778),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_840),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_789),
.B(n_340),
.C(n_676),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_744),
.A2(n_574),
.B(n_580),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_789),
.B(n_676),
.C(n_587),
.Y(n_896)
);

AO21x1_ASAP7_75t_L g897 ( 
.A1(n_704),
.A2(n_717),
.B(n_705),
.Y(n_897)
);

NOR2x1_ASAP7_75t_L g898 ( 
.A(n_798),
.B(n_608),
.Y(n_898)
);

INVx11_ASAP7_75t_L g899 ( 
.A(n_693),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_793),
.B(n_829),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_748),
.A2(n_624),
.B1(n_574),
.B2(n_598),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_744),
.A2(n_577),
.B(n_580),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_752),
.A2(n_624),
.B(n_637),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_731),
.B(n_719),
.C(n_839),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_744),
.A2(n_577),
.B(n_616),
.Y(n_905)
);

AO22x1_ASAP7_75t_L g906 ( 
.A1(n_817),
.A2(n_624),
.B1(n_678),
.B2(n_673),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_726),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_793),
.B(n_616),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_691),
.B(n_637),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_829),
.B(n_616),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_730),
.B(n_577),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_693),
.B(n_577),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_733),
.B(n_616),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_730),
.B(n_608),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_849),
.A2(n_624),
.B(n_637),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_744),
.A2(n_608),
.B(n_598),
.Y(n_916)
);

AO22x1_ASAP7_75t_L g917 ( 
.A1(n_817),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_917)
);

AOI21xp33_ASAP7_75t_L g918 ( 
.A1(n_719),
.A2(n_11),
.B(n_13),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_848),
.B(n_598),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_700),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_799),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_848),
.B(n_598),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_776),
.B(n_594),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_776),
.B(n_782),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_737),
.A2(n_176),
.B(n_163),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_737),
.A2(n_161),
.B(n_155),
.Y(n_926)
);

NAND2x1_ASAP7_75t_L g927 ( 
.A(n_722),
.B(n_144),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_833),
.B(n_14),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_743),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_839),
.A2(n_21),
.B(n_23),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_785),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_695),
.B(n_132),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_804),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_749),
.A2(n_759),
.B1(n_830),
.B2(n_703),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_756),
.A2(n_116),
.B(n_112),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_740),
.A2(n_741),
.B(n_771),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_786),
.B(n_26),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_802),
.A2(n_108),
.B(n_102),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_692),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_696),
.B(n_29),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_775),
.A2(n_101),
.B(n_96),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_706),
.B(n_30),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_743),
.A2(n_88),
.B(n_73),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_747),
.B(n_30),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_710),
.B(n_38),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_714),
.B(n_39),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_825),
.A2(n_39),
.B(n_40),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_787),
.A2(n_40),
.B(n_41),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_713),
.B(n_44),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_833),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_727),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_830),
.A2(n_44),
.B(n_45),
.C(n_47),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_781),
.A2(n_784),
.B(n_808),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_755),
.A2(n_59),
.B1(n_51),
.B2(n_53),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_806),
.B(n_48),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_733),
.B(n_51),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_796),
.A2(n_53),
.B(n_56),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_732),
.B(n_57),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_735),
.B(n_58),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_805),
.A2(n_58),
.B(n_803),
.Y(n_960)
);

AOI21xp33_ASAP7_75t_L g961 ( 
.A1(n_754),
.A2(n_773),
.B(n_820),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_736),
.B(n_761),
.Y(n_962)
);

BUFx12f_ASAP7_75t_L g963 ( 
.A(n_814),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_778),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_777),
.A2(n_779),
.B(n_739),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_734),
.Y(n_966)
);

AND2x6_ASAP7_75t_SL g967 ( 
.A(n_844),
.B(n_724),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_733),
.B(n_707),
.Y(n_968)
);

BUFx8_ASAP7_75t_L g969 ( 
.A(n_690),
.Y(n_969)
);

AND2x6_ASAP7_75t_L g970 ( 
.A(n_821),
.B(n_827),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_803),
.A2(n_811),
.B(n_850),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_809),
.B(n_745),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_707),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_746),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_853),
.B(n_742),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_811),
.A2(n_851),
.B(n_812),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_810),
.B(n_847),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_724),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_751),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_733),
.B(n_834),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_813),
.A2(n_822),
.B(n_823),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_794),
.B(n_724),
.Y(n_982)
);

OA21x2_ASAP7_75t_L g983 ( 
.A1(n_755),
.A2(n_841),
.B(n_852),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_753),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_787),
.A2(n_792),
.B(n_801),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_792),
.A2(n_801),
.B(n_770),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_844),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_760),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_720),
.A2(n_769),
.B(n_835),
.C(n_828),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_757),
.A2(n_758),
.B(n_766),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_762),
.A2(n_768),
.B(n_764),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_767),
.A2(n_824),
.B(n_838),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_718),
.B(n_846),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_844),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_780),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_832),
.A2(n_846),
.B(n_699),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_836),
.B(n_795),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_708),
.A2(n_826),
.B1(n_769),
.B2(n_797),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_780),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_843),
.B(n_845),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_780),
.Y(n_1001)
);

AOI21x1_ASAP7_75t_L g1002 ( 
.A1(n_697),
.A2(n_699),
.B(n_725),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_816),
.A2(n_818),
.B1(n_725),
.B2(n_697),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_815),
.B(n_831),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_780),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_845),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_828),
.A2(n_831),
.B1(n_837),
.B2(n_845),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_701),
.A2(n_702),
.B(n_698),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_788),
.B(n_715),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_788),
.B(n_715),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_711),
.A2(n_728),
.B(n_715),
.C(n_729),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_788),
.B(n_715),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_788),
.B(n_715),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_694),
.A2(n_650),
.B(n_698),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_694),
.A2(n_650),
.B(n_698),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_694),
.A2(n_650),
.B(n_698),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_807),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_729),
.B(n_551),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_694),
.A2(n_650),
.B(n_698),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_694),
.A2(n_650),
.B(n_698),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_729),
.B(n_551),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_711),
.A2(n_728),
.B(n_715),
.C(n_729),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_807),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_788),
.B(n_715),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_783),
.B(n_715),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_694),
.A2(n_650),
.B(n_698),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_788),
.B(n_715),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_709),
.A2(n_650),
.B(n_558),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_951),
.Y(n_1029)
);

AO31x2_ASAP7_75t_L g1030 ( 
.A1(n_897),
.A2(n_874),
.A3(n_870),
.B(n_996),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_859),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_1015),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_893),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_900),
.B(n_924),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_1015),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_878),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_920),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_904),
.A2(n_1027),
.B1(n_1024),
.B2(n_1025),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1019),
.A2(n_1026),
.B(n_1020),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1019),
.A2(n_1026),
.B(n_1020),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_857),
.B(n_975),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_878),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_996),
.A2(n_860),
.A3(n_865),
.B(n_862),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_994),
.B(n_912),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_886),
.B(n_949),
.C(n_997),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_SL g1048 ( 
.A1(n_888),
.A2(n_998),
.B(n_977),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_1018),
.B(n_1021),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_SL g1050 ( 
.A1(n_938),
.A2(n_948),
.B(n_947),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_993),
.A2(n_934),
.B1(n_1011),
.B2(n_1022),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_875),
.A2(n_884),
.B(n_885),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_973),
.B(n_858),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_855),
.A2(n_863),
.B(n_860),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_980),
.A2(n_873),
.B(n_1008),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_990),
.B(n_991),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_908),
.A2(n_910),
.B(n_981),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_864),
.A2(n_1004),
.B1(n_950),
.B2(n_987),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_981),
.A2(n_923),
.B(n_890),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_856),
.B(n_1017),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_984),
.B(n_937),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_883),
.A2(n_986),
.B(n_1028),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_855),
.A2(n_854),
.B(n_985),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_861),
.A2(n_976),
.B(n_953),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_867),
.A2(n_854),
.A3(n_960),
.B(n_861),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_1000),
.A2(n_919),
.B(n_922),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_990),
.B(n_991),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_913),
.A2(n_911),
.B(n_914),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_L g1069 ( 
.A1(n_868),
.A2(n_956),
.B(n_960),
.C(n_961),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1023),
.B(n_962),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_878),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_879),
.B(n_880),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_SL g1073 ( 
.A1(n_989),
.A2(n_1007),
.B(n_968),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_871),
.A2(n_872),
.B(n_1002),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_969),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_871),
.A2(n_872),
.B(n_869),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_954),
.B(n_930),
.C(n_952),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_944),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_882),
.A2(n_929),
.B1(n_965),
.B2(n_896),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_894),
.A2(n_1003),
.B(n_915),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_939),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_955),
.B(n_882),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_940),
.B(n_946),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_877),
.A2(n_931),
.B(n_933),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_972),
.B(n_881),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_928),
.B(n_907),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_942),
.B(n_945),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_891),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_969),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_958),
.B(n_959),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_881),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_898),
.B(n_912),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_881),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_895),
.A2(n_916),
.B(n_905),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_966),
.B(n_974),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_979),
.B(n_988),
.Y(n_1096)
);

AND2x2_ASAP7_75t_SL g1097 ( 
.A(n_889),
.B(n_892),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_887),
.B(n_978),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_892),
.A2(n_964),
.B1(n_901),
.B2(n_999),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_892),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_906),
.B(n_1005),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_902),
.A2(n_1001),
.B(n_1006),
.Y(n_1103)
);

AOI22x1_ASAP7_75t_L g1104 ( 
.A1(n_876),
.A2(n_941),
.B1(n_903),
.B2(n_926),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_964),
.B(n_995),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_970),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_964),
.B(n_932),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_927),
.A2(n_943),
.B(n_935),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_957),
.B(n_917),
.Y(n_1109)
);

BUFx12f_ASAP7_75t_L g1110 ( 
.A(n_967),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_970),
.B(n_909),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_925),
.A2(n_970),
.B(n_912),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_970),
.A2(n_909),
.B(n_899),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_970),
.A2(n_963),
.B(n_709),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_893),
.B(n_581),
.Y(n_1115)
);

AOI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_1015),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_969),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1018),
.B(n_1021),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1120)
);

AND3x4_ASAP7_75t_L g1121 ( 
.A(n_972),
.B(n_700),
.C(n_721),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_859),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1009),
.A2(n_1010),
.B(n_1013),
.C(n_1012),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1125)
);

NAND2x1_ASAP7_75t_L g1126 ( 
.A(n_882),
.B(n_722),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_900),
.A2(n_924),
.B(n_1009),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_900),
.A2(n_924),
.B(n_1009),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1009),
.A2(n_1010),
.B1(n_1013),
.B2(n_1012),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1009),
.A2(n_1010),
.B(n_1013),
.C(n_1012),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1009),
.A2(n_1010),
.B(n_1013),
.C(n_1012),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_900),
.A2(n_1027),
.B(n_1010),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_900),
.A2(n_924),
.B(n_1009),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_950),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_900),
.A2(n_924),
.B(n_1009),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_893),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_900),
.B(n_733),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

CKINVDCx8_ASAP7_75t_R g1148 ( 
.A(n_967),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_878),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_900),
.B(n_733),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_973),
.B(n_982),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_983),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_900),
.A2(n_924),
.B(n_1009),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_859),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_904),
.B(n_1025),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1008),
.A2(n_863),
.B(n_897),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_900),
.A2(n_924),
.B(n_1009),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_878),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_878),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_866),
.A2(n_992),
.B(n_971),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_899),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1014),
.A2(n_709),
.B(n_1015),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_1015),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1044),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1162),
.A2(n_1047),
.B(n_1048),
.C(n_1140),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1056),
.A2(n_1067),
.B(n_1131),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1160),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1092),
.B(n_1113),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1029),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1141),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1130),
.B(n_1118),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1154),
.B(n_1174),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1120),
.A2(n_1142),
.B1(n_1139),
.B2(n_1150),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1092),
.B(n_1044),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1141),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1061),
.B(n_1040),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1119),
.B(n_1086),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1044),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1049),
.B(n_1043),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1125),
.B(n_1129),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1156),
.A2(n_1169),
.B1(n_1132),
.B2(n_1136),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1147),
.Y(n_1195)
);

INVx2_ASAP7_75t_R g1196 ( 
.A(n_1106),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1124),
.B(n_1132),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1162),
.B(n_1144),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1033),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1074),
.A2(n_1076),
.B(n_1062),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1160),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_1057),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1123),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1115),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1124),
.B(n_1136),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1174),
.B(n_1053),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1143),
.A2(n_1157),
.B1(n_1167),
.B2(n_1070),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1072),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1064),
.A2(n_1068),
.B(n_1054),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1123),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1095),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1044),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1036),
.B(n_1039),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1134),
.A2(n_1158),
.B(n_1175),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1071),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1038),
.B(n_1031),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1078),
.B(n_1034),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1117),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1105),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1036),
.B(n_1034),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1096),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1117),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1135),
.A2(n_1161),
.B(n_1146),
.Y(n_1224)
);

AOI21xp33_ASAP7_75t_L g1225 ( 
.A1(n_1051),
.A2(n_1077),
.B(n_1109),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_L g1226 ( 
.A(n_1060),
.B(n_1083),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1097),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1075),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1087),
.B(n_1090),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1082),
.B(n_1081),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1097),
.Y(n_1231)
);

INVx8_ASAP7_75t_L g1232 ( 
.A(n_1071),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1137),
.B(n_1077),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1085),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1098),
.B(n_1088),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1163),
.B(n_1073),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1046),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1149),
.A2(n_1168),
.B(n_1164),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1032),
.A2(n_1035),
.B(n_1041),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1058),
.B(n_1099),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1107),
.B(n_1105),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1063),
.A2(n_1042),
.B(n_1069),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1075),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1089),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1172),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1052),
.A2(n_1176),
.B(n_1116),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1121),
.A2(n_1080),
.B1(n_1102),
.B2(n_1085),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1071),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1071),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1172),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1037),
.Y(n_1251)
);

NOR2xp67_ASAP7_75t_L g1252 ( 
.A(n_1114),
.B(n_1107),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1037),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1151),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1091),
.Y(n_1255)
);

INVx5_ASAP7_75t_L g1256 ( 
.A(n_1091),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1089),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1102),
.B(n_1145),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1091),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1093),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1163),
.B(n_1145),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1151),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1046),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_SL g1264 ( 
.A1(n_1084),
.A2(n_1079),
.B(n_1103),
.C(n_1171),
.Y(n_1264)
);

CKINVDCx6p67_ASAP7_75t_R g1265 ( 
.A(n_1046),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1163),
.B(n_1153),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1171),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1155),
.B(n_1045),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1111),
.B(n_1101),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1093),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1066),
.A2(n_1108),
.B(n_1050),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1045),
.B(n_1030),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1100),
.A2(n_1104),
.B1(n_1093),
.B2(n_1101),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1110),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1093),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1101),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1101),
.B(n_1112),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1126),
.A2(n_1148),
.B1(n_1110),
.B2(n_1030),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1045),
.B(n_1030),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1094),
.B(n_1152),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1122),
.A2(n_1159),
.B1(n_1170),
.B2(n_1133),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1030),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1065),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1065),
.B(n_1138),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1165),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1166),
.A2(n_1173),
.B(n_904),
.C(n_1009),
.Y(n_1286)
);

INVx5_ASAP7_75t_L g1287 ( 
.A(n_1044),
.Y(n_1287)
);

BUFx5_ASAP7_75t_L g1288 ( 
.A(n_1106),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1029),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_R g1290 ( 
.A(n_1141),
.B(n_565),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1144),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1162),
.A2(n_904),
.B(n_1010),
.C(n_1009),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1047),
.B(n_1025),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1154),
.B(n_1174),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1118),
.A2(n_1009),
.B1(n_1012),
.B2(n_1010),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1044),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1061),
.B(n_1119),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1160),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1130),
.B(n_1118),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1049),
.B(n_1043),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1044),
.Y(n_1301)
);

AO32x1_ASAP7_75t_L g1302 ( 
.A1(n_1051),
.A2(n_1109),
.A3(n_954),
.B1(n_1079),
.B2(n_1130),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1044),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1174),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1141),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_L g1306 ( 
.A(n_1047),
.B(n_1009),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1047),
.A2(n_904),
.B1(n_900),
.B2(n_1162),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1144),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1029),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1061),
.B(n_1119),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1092),
.B(n_878),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1154),
.B(n_1174),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1029),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1047),
.B(n_1061),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1029),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1047),
.B(n_900),
.C(n_904),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1047),
.B(n_1061),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1154),
.B(n_1174),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1056),
.A2(n_1067),
.B(n_936),
.Y(n_1319)
);

CKINVDCx8_ASAP7_75t_R g1320 ( 
.A(n_1141),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1056),
.A2(n_1067),
.B(n_936),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1293),
.A2(n_1307),
.B1(n_1316),
.B2(n_1306),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1291),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1277),
.Y(n_1324)
);

BUFx2_ASAP7_75t_R g1325 ( 
.A(n_1320),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1220),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1178),
.B(n_1292),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1316),
.A2(n_1247),
.B1(n_1225),
.B2(n_1189),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1183),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1202),
.A2(n_1210),
.B(n_1239),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1289),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1227),
.A2(n_1231),
.B1(n_1198),
.B2(n_1295),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1256),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1291),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1313),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1308),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1315),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1219),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1195),
.Y(n_1339)
);

BUFx4f_ASAP7_75t_SL g1340 ( 
.A(n_1304),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1186),
.B(n_1184),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1243),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1193),
.A2(n_1186),
.B1(n_1299),
.B2(n_1184),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1309),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1319),
.A2(n_1321),
.B(n_1215),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1271),
.A2(n_1246),
.B(n_1200),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1235),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1225),
.A2(n_1317),
.B1(n_1314),
.B2(n_1258),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_1188),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1256),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1179),
.A2(n_1224),
.B(n_1238),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1308),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1230),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1209),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1204),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1226),
.A2(n_1278),
.B1(n_1310),
.B2(n_1297),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1204),
.A2(n_1300),
.B1(n_1192),
.B2(n_1295),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1245),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1221),
.A2(n_1190),
.B1(n_1241),
.B2(n_1299),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1207),
.A2(n_1234),
.B1(n_1278),
.B2(n_1208),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1228),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1252),
.B(n_1283),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1240),
.A2(n_1208),
.B(n_1194),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1234),
.A2(n_1194),
.B1(n_1218),
.B2(n_1214),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1280),
.A2(n_1242),
.B(n_1281),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1212),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1286),
.A2(n_1233),
.B(n_1205),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1222),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1214),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1201),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1206),
.B(n_1211),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1250),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1199),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1284),
.B(n_1282),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1268),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1290),
.Y(n_1376)
);

AO21x1_ASAP7_75t_L g1377 ( 
.A1(n_1233),
.A2(n_1197),
.B(n_1205),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1285),
.B(n_1236),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1305),
.A2(n_1223),
.B1(n_1274),
.B2(n_1244),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1253),
.Y(n_1380)
);

CKINVDCx11_ASAP7_75t_R g1381 ( 
.A(n_1257),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1197),
.A2(n_1263),
.B1(n_1237),
.B2(n_1203),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1206),
.A2(n_1318),
.B1(n_1294),
.B2(n_1185),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1181),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1269),
.B(n_1213),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1236),
.A2(n_1264),
.B(n_1272),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1269),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1273),
.A2(n_1181),
.B(n_1266),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1187),
.B(n_1311),
.Y(n_1389)
);

AO21x1_ASAP7_75t_L g1390 ( 
.A1(n_1273),
.A2(n_1272),
.B(n_1279),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1177),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1261),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1217),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1185),
.B(n_1318),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1187),
.B(n_1311),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1254),
.Y(n_1396)
);

AO21x1_ASAP7_75t_L g1397 ( 
.A1(n_1261),
.A2(n_1266),
.B(n_1302),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1288),
.Y(n_1398)
);

BUFx8_ASAP7_75t_L g1399 ( 
.A(n_1294),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1262),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1267),
.A2(n_1251),
.B(n_1270),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1265),
.A2(n_1312),
.B1(n_1180),
.B2(n_1298),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1216),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1312),
.A2(n_1255),
.B(n_1216),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1259),
.A2(n_1287),
.B1(n_1302),
.B2(n_1248),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1259),
.B(n_1287),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1177),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1301),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1301),
.A2(n_1196),
.B(n_1302),
.Y(n_1409)
);

AO21x1_ASAP7_75t_L g1410 ( 
.A1(n_1260),
.A2(n_1275),
.B(n_1287),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1259),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1260),
.A2(n_1275),
.B(n_1191),
.Y(n_1412)
);

NAND2x1p5_ASAP7_75t_L g1413 ( 
.A(n_1177),
.B(n_1191),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1249),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1232),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1249),
.B(n_1276),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1276),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1232),
.A2(n_1303),
.B1(n_1276),
.B2(n_1296),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1296),
.A2(n_1303),
.B(n_1271),
.Y(n_1419)
);

AOI21xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1296),
.A2(n_466),
.B(n_464),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1303),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1293),
.B(n_370),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1201),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1293),
.A2(n_904),
.B1(n_1047),
.B2(n_900),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1182),
.Y(n_1425)
);

BUFx2_ASAP7_75t_R g1426 ( 
.A(n_1320),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1182),
.Y(n_1427)
);

AOI222xp33_ASAP7_75t_L g1428 ( 
.A1(n_1293),
.A2(n_904),
.B1(n_562),
.B2(n_1162),
.C1(n_817),
.C2(n_928),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1293),
.A2(n_904),
.B1(n_886),
.B2(n_928),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1220),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1182),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1256),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1193),
.B(n_1229),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1293),
.A2(n_904),
.B1(n_1047),
.B2(n_900),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1233),
.B(n_1197),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1277),
.B(n_1252),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1277),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1269),
.B(n_1241),
.Y(n_1438)
);

BUFx2_ASAP7_75t_SL g1439 ( 
.A(n_1256),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1291),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1326),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1330),
.A2(n_1345),
.B(n_1390),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1327),
.B(n_1375),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1362),
.B(n_1388),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1392),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1327),
.B(n_1369),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1355),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1367),
.B(n_1438),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1438),
.B(n_1324),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1438),
.B(n_1324),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1374),
.B(n_1435),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_R g1452 ( 
.A(n_1342),
.B(n_1338),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1343),
.B(n_1435),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1346),
.A2(n_1351),
.B(n_1365),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1378),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1390),
.A2(n_1409),
.B(n_1363),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1341),
.B(n_1433),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1378),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1437),
.B(n_1384),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1388),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1386),
.B(n_1339),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1386),
.B(n_1357),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1377),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1326),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1386),
.B(n_1339),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1377),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1430),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1430),
.Y(n_1468)
);

BUFx12f_ASAP7_75t_L g1469 ( 
.A(n_1338),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1397),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1397),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1344),
.B(n_1364),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1429),
.A2(n_1322),
.B(n_1424),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1419),
.A2(n_1409),
.B(n_1436),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1360),
.A2(n_1328),
.B(n_1348),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1323),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1334),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1336),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1359),
.B(n_1356),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1398),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1398),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1434),
.B(n_1353),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1387),
.B(n_1331),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1354),
.B(n_1347),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1352),
.Y(n_1485)
);

CKINVDCx10_ASAP7_75t_R g1486 ( 
.A(n_1325),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1358),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1362),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

AO21x1_ASAP7_75t_L g1491 ( 
.A1(n_1362),
.A2(n_1401),
.B(n_1372),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1428),
.A2(n_1332),
.B(n_1405),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1436),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1412),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1380),
.A2(n_1400),
.B(n_1396),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1440),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1335),
.B(n_1382),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1393),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1371),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1373),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1404),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1337),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1385),
.B(n_1425),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1389),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1427),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1399),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1412),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1422),
.A2(n_1383),
.B1(n_1376),
.B2(n_1402),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1385),
.B(n_1431),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1451),
.B(n_1417),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1494),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1486),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1492),
.A2(n_1376),
.B1(n_1394),
.B2(n_1350),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1448),
.B(n_1395),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1448),
.B(n_1395),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1461),
.B(n_1408),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1461),
.B(n_1403),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1465),
.B(n_1391),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1465),
.B(n_1391),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1456),
.B(n_1391),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1453),
.B(n_1411),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1453),
.B(n_1412),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1464),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1490),
.B(n_1416),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1456),
.B(n_1470),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1480),
.B(n_1416),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1457),
.B(n_1420),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1473),
.A2(n_1492),
.B1(n_1475),
.B2(n_1479),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1451),
.B(n_1462),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1416),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1457),
.B(n_1414),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1444),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1456),
.B(n_1413),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1456),
.B(n_1421),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1495),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1495),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1495),
.Y(n_1537)
);

INVxp33_ASAP7_75t_L g1538 ( 
.A(n_1452),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1481),
.B(n_1449),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_SL g1540 ( 
.A(n_1452),
.B(n_1426),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1445),
.B(n_1333),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1462),
.B(n_1423),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1490),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1486),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1488),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1493),
.Y(n_1546)
);

INVxp67_ASAP7_75t_SL g1547 ( 
.A(n_1491),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1471),
.B(n_1370),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1488),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1444),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_L g1551 ( 
.A(n_1528),
.B(n_1473),
.C(n_1475),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1521),
.B(n_1499),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1513),
.B(n_1482),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1521),
.B(n_1447),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1527),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1539),
.B(n_1481),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1513),
.A2(n_1508),
.B1(n_1475),
.B2(n_1527),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1464),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1540),
.B(n_1482),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1540),
.B(n_1501),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1538),
.A2(n_1508),
.B1(n_1475),
.B2(n_1479),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1542),
.B(n_1500),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1510),
.B(n_1467),
.Y(n_1563)
);

AND2x2_ASAP7_75t_SL g1564 ( 
.A(n_1532),
.B(n_1442),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1510),
.B(n_1477),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1455),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1542),
.A2(n_1446),
.B(n_1472),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1518),
.B(n_1455),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1547),
.B(n_1497),
.C(n_1463),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1512),
.A2(n_1469),
.B1(n_1500),
.B2(n_1379),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1522),
.A2(n_1446),
.B(n_1472),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1514),
.B(n_1496),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1515),
.B(n_1498),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1531),
.A2(n_1506),
.B1(n_1469),
.B2(n_1497),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1515),
.B(n_1441),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1522),
.B(n_1441),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1531),
.B(n_1469),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1549),
.B(n_1441),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1549),
.B(n_1468),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1478),
.C(n_1476),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1468),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1518),
.B(n_1458),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1548),
.B(n_1505),
.C(n_1502),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1526),
.A2(n_1506),
.B1(n_1443),
.B2(n_1509),
.Y(n_1585)
);

AND2x2_ASAP7_75t_SL g1586 ( 
.A(n_1532),
.B(n_1442),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1535),
.A2(n_1474),
.B(n_1454),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1519),
.B(n_1458),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1534),
.B(n_1543),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1516),
.B(n_1517),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1525),
.A2(n_1484),
.B1(n_1466),
.B2(n_1463),
.C(n_1487),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1548),
.B(n_1506),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1550),
.A2(n_1443),
.B(n_1466),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1524),
.A2(n_1450),
.B1(n_1449),
.B2(n_1489),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1534),
.B(n_1507),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1517),
.B(n_1504),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1517),
.B(n_1504),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1541),
.B(n_1442),
.C(n_1460),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1534),
.B(n_1507),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1526),
.B(n_1483),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1525),
.A2(n_1484),
.B1(n_1487),
.B2(n_1503),
.C(n_1509),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1530),
.B(n_1483),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1524),
.A2(n_1450),
.B1(n_1489),
.B2(n_1459),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_L g1604 ( 
.A(n_1544),
.B(n_1432),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1589),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1595),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1577),
.B(n_1529),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1589),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1551),
.A2(n_1442),
.B(n_1491),
.Y(n_1610)
);

CKINVDCx16_ASAP7_75t_R g1611 ( 
.A(n_1571),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1578),
.B(n_1349),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1599),
.B(n_1533),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1587),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1556),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1533),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1587),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1525),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1566),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1569),
.B(n_1532),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1570),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1555),
.B(n_1535),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1554),
.B(n_1543),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1565),
.B(n_1546),
.Y(n_1627)
);

NAND2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1564),
.B(n_1532),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1572),
.B(n_1536),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1579),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1552),
.B(n_1536),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1571),
.B(n_1559),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1587),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1564),
.B(n_1520),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1586),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1596),
.B(n_1537),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1537),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1584),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1558),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1584),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1600),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1586),
.B(n_1520),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1636),
.B(n_1532),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1629),
.B(n_1574),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1611),
.B(n_1632),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1634),
.B(n_1586),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_SL g1648 ( 
.A(n_1611),
.B(n_1551),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1609),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1634),
.B(n_1532),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1622),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1606),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1635),
.B(n_1532),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1507),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1615),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1640),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1637),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1629),
.B(n_1567),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1638),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1573),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1635),
.B(n_1593),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1643),
.B(n_1568),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1643),
.B(n_1576),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1614),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1640),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1638),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1641),
.B(n_1581),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1606),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1628),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1622),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1621),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1613),
.B(n_1622),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1620),
.B(n_1598),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1621),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1636),
.B(n_1511),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1627),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1620),
.B(n_1580),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1649),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1668),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1649),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1628),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1671),
.B(n_1610),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1651),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1672),
.B(n_1623),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1646),
.A2(n_1557),
.B1(n_1561),
.B2(n_1553),
.C(n_1581),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1647),
.B(n_1628),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1648),
.B(n_1575),
.C(n_1560),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1655),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1665),
.B(n_1622),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1645),
.B(n_1612),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1665),
.B(n_1616),
.Y(n_1698)
);

OAI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1678),
.A2(n_1585),
.B1(n_1630),
.B2(n_1607),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1678),
.B(n_1631),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1681),
.A2(n_1604),
.B1(n_1601),
.B2(n_1562),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1659),
.B(n_1631),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1664),
.B(n_1616),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1659),
.B(n_1625),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.B(n_1624),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1651),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1652),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1677),
.B(n_1650),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1656),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1660),
.B(n_1625),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1657),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1656),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1658),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1669),
.B(n_1618),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1660),
.B(n_1662),
.Y(n_1716)
);

CKINVDCx16_ASAP7_75t_R g1717 ( 
.A(n_1650),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1658),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1662),
.B(n_1607),
.Y(n_1719)
);

OAI32xp33_ASAP7_75t_L g1720 ( 
.A1(n_1655),
.A2(n_1617),
.A3(n_1630),
.B1(n_1619),
.B2(n_1626),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1645),
.B(n_1342),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1677),
.B(n_1624),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1668),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1676),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1676),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1668),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1661),
.B(n_1618),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1709),
.B(n_1652),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1712),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1709),
.B(n_1674),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1696),
.B(n_1675),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1700),
.B(n_1670),
.Y(n_1734)
);

XOR2xp5_ASAP7_75t_L g1735 ( 
.A(n_1694),
.B(n_1702),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1721),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1708),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1675),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1686),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1700),
.B(n_1670),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1689),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1697),
.B(n_1661),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1692),
.A2(n_1644),
.B1(n_1604),
.B2(n_1682),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1727),
.B(n_1682),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1707),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1708),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1690),
.B(n_1329),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1695),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1688),
.A2(n_1644),
.B1(n_1666),
.B2(n_1654),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1687),
.B(n_1654),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1687),
.B(n_1693),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1710),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1693),
.B(n_1644),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1699),
.B(n_1644),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1698),
.B(n_1683),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1715),
.B(n_1329),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1713),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1679),
.Y(n_1759)
);

OAI21xp33_ASAP7_75t_L g1760 ( 
.A1(n_1688),
.A2(n_1655),
.B(n_1585),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1688),
.A2(n_1630),
.B1(n_1619),
.B2(n_1680),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1714),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1730),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1735),
.A2(n_1688),
.B1(n_1716),
.B2(n_1695),
.C(n_1691),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1730),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1752),
.B(n_1704),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1760),
.A2(n_1720),
.B(n_1695),
.C(n_1701),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1735),
.A2(n_1706),
.B1(n_1719),
.B2(n_1722),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1739),
.Y(n_1770)
);

AOI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1736),
.A2(n_1720),
.B(n_1716),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1746),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1743),
.A2(n_1731),
.B1(n_1762),
.B2(n_1749),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1752),
.B(n_1706),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1746),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1729),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1739),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1742),
.A2(n_1755),
.B(n_1728),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1756),
.B(n_1722),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1728),
.A2(n_1724),
.B(n_1718),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1747),
.A2(n_1725),
.B(n_1703),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1737),
.B(n_1703),
.C(n_1705),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1751),
.B(n_1705),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1667),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_SL g1786 ( 
.A1(n_1757),
.A2(n_1594),
.B(n_1711),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1737),
.A2(n_1711),
.B(n_1685),
.Y(n_1788)
);

OAI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1750),
.A2(n_1619),
.B1(n_1608),
.B2(n_1605),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1770),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1778),
.B(n_1744),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1770),
.Y(n_1792)
);

OAI31xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1773),
.A2(n_1732),
.A3(n_1733),
.B(n_1761),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1767),
.B(n_1751),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1768),
.A2(n_1744),
.B1(n_1740),
.B2(n_1734),
.C(n_1758),
.Y(n_1795)
);

AO22x2_ASAP7_75t_L g1796 ( 
.A1(n_1772),
.A2(n_1763),
.B1(n_1745),
.B2(n_1753),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1772),
.B(n_1761),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1765),
.A2(n_1763),
.B1(n_1745),
.B2(n_1753),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1775),
.B(n_1732),
.Y(n_1799)
);

NAND2x1p5_ASAP7_75t_L g1800 ( 
.A(n_1775),
.B(n_1748),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1777),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1769),
.B(n_1754),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1776),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1754),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1776),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1767),
.B(n_1738),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1774),
.B(n_1738),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1774),
.B(n_1733),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1781),
.B(n_1733),
.Y(n_1809)
);

AOI32xp33_ASAP7_75t_L g1810 ( 
.A1(n_1795),
.A2(n_1789),
.A3(n_1784),
.B1(n_1764),
.B2(n_1782),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1798),
.B(n_1768),
.C(n_1771),
.Y(n_1811)
);

AOI322xp5_ASAP7_75t_L g1812 ( 
.A1(n_1791),
.A2(n_1783),
.A3(n_1779),
.B1(n_1785),
.B2(n_1784),
.C1(n_1787),
.C2(n_1766),
.Y(n_1812)
);

OAI21xp33_ASAP7_75t_SL g1813 ( 
.A1(n_1793),
.A2(n_1780),
.B(n_1788),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1791),
.B(n_1777),
.C(n_1748),
.Y(n_1814)
);

AOI211xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1799),
.A2(n_1748),
.B(n_1340),
.C(n_1758),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1796),
.Y(n_1816)
);

AOI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1804),
.A2(n_1734),
.B(n_1740),
.C(n_1733),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1809),
.A2(n_1729),
.B(n_1759),
.Y(n_1818)
);

NAND2x1_ASAP7_75t_L g1819 ( 
.A(n_1808),
.B(n_1729),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1797),
.A2(n_1729),
.B(n_1759),
.C(n_1685),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1798),
.A2(n_1726),
.B(n_1723),
.Y(n_1821)
);

AOI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1802),
.A2(n_1726),
.B1(n_1723),
.B2(n_1617),
.C(n_1633),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1816),
.Y(n_1823)
);

NAND3xp33_ASAP7_75t_SL g1824 ( 
.A(n_1811),
.B(n_1800),
.C(n_1805),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_SL g1825 ( 
.A(n_1814),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1813),
.A2(n_1794),
.B1(n_1806),
.B2(n_1807),
.Y(n_1826)
);

NAND4xp75_ASAP7_75t_L g1827 ( 
.A(n_1818),
.B(n_1801),
.C(n_1790),
.D(n_1792),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1810),
.A2(n_1796),
.B(n_1800),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_L g1829 ( 
.A(n_1817),
.B(n_1803),
.C(n_1381),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_L g1830 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1820),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1821),
.Y(n_1832)
);

NAND4xp25_ASAP7_75t_L g1833 ( 
.A(n_1815),
.B(n_1796),
.C(n_1423),
.D(n_1370),
.Y(n_1833)
);

OAI321xp33_ASAP7_75t_L g1834 ( 
.A1(n_1824),
.A2(n_1828),
.A3(n_1833),
.B1(n_1831),
.B2(n_1826),
.C(n_1832),
.Y(n_1834)
);

OAI211xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1829),
.A2(n_1812),
.B(n_1822),
.C(n_1361),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1823),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1830),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1827),
.Y(n_1838)
);

NOR3xp33_ASAP7_75t_L g1839 ( 
.A(n_1825),
.B(n_1381),
.C(n_1361),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1837),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1836),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1838),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1839),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1834),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1835),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1836),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1842),
.A2(n_1679),
.B1(n_1673),
.B2(n_1653),
.C(n_1627),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_SL g1848 ( 
.A(n_1840),
.B(n_1349),
.C(n_1406),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1841),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1842),
.B(n_1667),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1843),
.B(n_1349),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1846),
.Y(n_1852)
);

XNOR2x1_ASAP7_75t_L g1853 ( 
.A(n_1851),
.B(n_1844),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1850),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1849),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1855),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1856),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1845),
.B1(n_1854),
.B2(n_1855),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1857),
.A2(n_1845),
.B1(n_1853),
.B2(n_1849),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1852),
.B(n_1847),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1858),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1860),
.A2(n_1852),
.B(n_1848),
.Y(n_1862)
);

AOI31xp33_ASAP7_75t_L g1863 ( 
.A1(n_1861),
.A2(n_1406),
.A3(n_1410),
.B(n_1418),
.Y(n_1863)
);

XNOR2xp5_ASAP7_75t_L g1864 ( 
.A(n_1862),
.B(n_1860),
.Y(n_1864)
);

XNOR2xp5_ASAP7_75t_L g1865 ( 
.A(n_1864),
.B(n_1860),
.Y(n_1865)
);

OAI221xp5_ASAP7_75t_R g1866 ( 
.A1(n_1865),
.A2(n_1863),
.B1(n_1603),
.B2(n_1407),
.C(n_1439),
.Y(n_1866)
);

AOI211xp5_ASAP7_75t_L g1867 ( 
.A1(n_1866),
.A2(n_1415),
.B(n_1432),
.C(n_1680),
.Y(n_1867)
);


endmodule