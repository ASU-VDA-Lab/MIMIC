module fake_jpeg_1994_n_455 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_455);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_74),
.Y(n_115)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_76),
.A2(n_93),
.B1(n_7),
.B2(n_8),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_14),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_27),
.C(n_26),
.Y(n_122)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_14),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_3),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_19),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_100),
.Y(n_147)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_19),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_108),
.Y(n_164)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_105),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_110),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_28),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_114),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_22),
.B1(n_48),
.B2(n_37),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_119),
.A2(n_121),
.B1(n_145),
.B2(n_150),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_22),
.B1(n_48),
.B2(n_41),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_122),
.B(n_149),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_109),
.B1(n_112),
.B2(n_111),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_123),
.A2(n_152),
.B1(n_166),
.B2(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_41),
.C(n_28),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_187),
.C(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_57),
.B(n_47),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_131),
.B(n_139),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_144),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_27),
.B1(n_50),
.B2(n_39),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_138),
.A2(n_156),
.B1(n_134),
.B2(n_167),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_83),
.B(n_50),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_39),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_72),
.A2(n_32),
.B1(n_38),
.B2(n_44),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_94),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_78),
.B(n_4),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_151),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_84),
.B(n_7),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_158),
.B(n_174),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_67),
.A2(n_9),
.B1(n_10),
.B2(n_68),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_106),
.B(n_82),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_88),
.A2(n_114),
.B1(n_104),
.B2(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_89),
.B(n_99),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_183),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_86),
.B(n_76),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_70),
.B(n_105),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_188),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_105),
.A2(n_31),
.B1(n_23),
.B2(n_74),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_187),
.A2(n_150),
.B1(n_166),
.B2(n_145),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_61),
.B(n_91),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_126),
.A2(n_147),
.A3(n_128),
.B1(n_127),
.B2(n_157),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_191),
.A2(n_218),
.B(n_214),
.Y(n_284)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_193),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_140),
.B(n_172),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_195),
.B(n_232),
.C(n_250),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_160),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_213),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_204),
.B(n_211),
.Y(n_262)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

BUFx8_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_133),
.B(n_153),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_212),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_141),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_118),
.Y(n_217)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

OR2x4_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_138),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_129),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_220),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_175),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_123),
.A2(n_119),
.B1(n_121),
.B2(n_152),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_201),
.B1(n_218),
.B2(n_234),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_153),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_227),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_115),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_230),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_120),
.B(n_136),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_231),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_186),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_249),
.Y(n_263)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_236),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_116),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_239),
.Y(n_299)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_185),
.B1(n_115),
.B2(n_137),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_241),
.A2(n_252),
.B1(n_199),
.B2(n_242),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_173),
.B(n_124),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_242),
.Y(n_280)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_244),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_163),
.B(n_167),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_177),
.B(n_178),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_134),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_116),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_169),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_142),
.B(n_177),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_224),
.B(n_217),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_261),
.A2(n_285),
.B1(n_269),
.B2(n_268),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_268),
.B(n_222),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_195),
.B(n_192),
.C(n_196),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_286),
.C(n_290),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_198),
.A2(n_214),
.B(n_240),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_247),
.B(n_248),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_214),
.B1(n_240),
.B2(n_223),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_205),
.B1(n_243),
.B2(n_230),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_207),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_233),
.A2(n_215),
.B1(n_253),
.B2(n_203),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_242),
.C(n_202),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_191),
.B(n_231),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_212),
.A2(n_235),
.B1(n_229),
.B2(n_210),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_296),
.B1(n_207),
.B2(n_280),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_303),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_261),
.A2(n_228),
.B1(n_216),
.B2(n_200),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_301),
.A2(n_306),
.B1(n_317),
.B2(n_297),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_302),
.B(n_266),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_318),
.B(n_314),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_310),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_221),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_316),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_321),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_313),
.A2(n_297),
.B1(n_293),
.B2(n_283),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_272),
.B1(n_256),
.B2(n_290),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_315),
.A2(n_327),
.B1(n_332),
.B2(n_308),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_276),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_284),
.A2(n_285),
.B1(n_279),
.B2(n_259),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_259),
.A2(n_265),
.B(n_254),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_320),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_260),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_263),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_326),
.Y(n_359)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_324),
.B(n_331),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_325),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_259),
.A2(n_286),
.B1(n_270),
.B2(n_271),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_266),
.Y(n_328)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_255),
.A2(n_264),
.B(n_257),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_293),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_260),
.A2(n_298),
.B1(n_294),
.B2(n_283),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_257),
.B(n_267),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_289),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_294),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_334),
.B(n_277),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_336),
.A2(n_321),
.B1(n_324),
.B2(n_331),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_354),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_343),
.A2(n_345),
.B(n_307),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_255),
.B(n_277),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_339),
.B(n_350),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_357),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_334),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_355),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_325),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_281),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_357),
.C(n_302),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_273),
.C(n_292),
.Y(n_357)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_315),
.A2(n_273),
.A3(n_291),
.B1(n_292),
.B2(n_319),
.C1(n_323),
.C2(n_326),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_333),
.C(n_303),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_352),
.B1(n_360),
.B2(n_317),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_362),
.A2(n_366),
.B1(n_367),
.B2(n_376),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_359),
.A2(n_312),
.B1(n_311),
.B2(n_327),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_377),
.B1(n_344),
.B2(n_348),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_360),
.A2(n_301),
.B1(n_318),
.B2(n_329),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_360),
.A2(n_320),
.B1(n_332),
.B2(n_316),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_374),
.C(n_353),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_305),
.Y(n_369)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_369),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_378),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_382),
.B1(n_340),
.B2(n_351),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_373),
.A2(n_375),
.B(n_379),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_310),
.C(n_322),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_360),
.A2(n_328),
.B1(n_330),
.B2(n_291),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_359),
.A2(n_330),
.B1(n_345),
.B2(n_343),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_338),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_354),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g381 ( 
.A(n_349),
.B(n_358),
.CI(n_354),
.CON(n_381),
.SN(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_346),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_338),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_364),
.A2(n_348),
.B1(n_340),
.B2(n_351),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_389),
.B1(n_394),
.B2(n_395),
.Y(n_402)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_393),
.Y(n_406)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_390),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_371),
.B(n_342),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_397),
.C(n_382),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_374),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_363),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_396),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_347),
.C(n_355),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_341),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_372),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_392),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_390),
.A2(n_361),
.B(n_373),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_393),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_399),
.A2(n_377),
.B1(n_362),
.B2(n_365),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_404),
.A2(n_410),
.B1(n_414),
.B2(n_389),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_391),
.B(n_361),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_405),
.B(n_398),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_400),
.A2(n_379),
.B(n_370),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_412),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_383),
.A2(n_378),
.B1(n_366),
.B2(n_376),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_399),
.A2(n_372),
.B1(n_381),
.B2(n_347),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_397),
.Y(n_415)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_416),
.B(n_417),
.Y(n_428)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_411),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_418),
.A2(n_411),
.B(n_400),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_402),
.A2(n_387),
.B1(n_413),
.B2(n_395),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_419),
.A2(n_396),
.B1(n_407),
.B2(n_384),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_422),
.B(n_404),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_401),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_423),
.B(n_424),
.C(n_412),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_426),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_414),
.C(n_385),
.Y(n_426)
);

AOI21x1_ASAP7_75t_L g436 ( 
.A1(n_427),
.A2(n_408),
.B(n_388),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_430),
.Y(n_439)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_422),
.Y(n_432)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_432),
.Y(n_438)
);

BUFx24_ASAP7_75t_SL g433 ( 
.A(n_420),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_433),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_432),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_420),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_429),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_442),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_426),
.C(n_425),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_444),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_439),
.A2(n_403),
.B(n_388),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_445),
.A2(n_439),
.B(n_437),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g449 ( 
.A1(n_447),
.A2(n_441),
.B(n_386),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_449),
.B(n_450),
.C(n_446),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_440),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_448),
.B(n_434),
.Y(n_452)
);

OAI21x1_ASAP7_75t_SL g453 ( 
.A1(n_452),
.A2(n_386),
.B(n_381),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_381),
.B1(n_405),
.B2(n_341),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_337),
.Y(n_455)
);


endmodule