module real_jpeg_13460_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_309, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_309;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx10_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_32),
.B1(n_35),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_44),
.B1(n_49),
.B2(n_67),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_133),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_133),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_4),
.A2(n_44),
.B1(n_49),
.B2(n_133),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_44),
.B1(n_49),
.B2(n_59),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_7),
.A2(n_32),
.B1(n_35),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_7),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_170),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_7),
.A2(n_44),
.B1(n_49),
.B2(n_170),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_29),
.B1(n_44),
.B2(n_49),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_91),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_91),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_12),
.A2(n_44),
.B1(n_49),
.B2(n_91),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_13),
.B(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_13),
.A2(n_27),
.B(n_197),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_188),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_48),
.B(n_52),
.C(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_13),
.B(n_68),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_13),
.B(n_84),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_13),
.B(n_42),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_13),
.A2(n_35),
.B(n_60),
.C(n_259),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_38),
.B1(n_44),
.B2(n_49),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_15),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_157),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_15),
.A2(n_44),
.B1(n_49),
.B2(n_157),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_16),
.A2(n_44),
.B1(n_49),
.B2(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_16),
.A2(n_32),
.B1(n_35),
.B2(n_55),
.Y(n_101)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_92),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_22),
.B(n_92),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_70),
.C(n_77),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_70),
.B1(n_71),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_24),
.A2(n_25),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_41),
.C(n_57),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_27),
.A2(n_32),
.A3(n_34),
.B1(n_198),
.B2(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_28),
.B(n_188),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_30),
.A2(n_31),
.B1(n_37),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_30),
.A2(n_31),
.B1(n_90),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_30),
.A2(n_31),
.B1(n_132),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_30),
.A2(n_31),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_30),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_31),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_32),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_32),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_33),
.B(n_35),
.Y(n_212)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_35),
.A2(n_53),
.A3(n_62),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_41),
.A2(n_69),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_50),
.B(n_54),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_50),
.B1(n_54),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_50),
.B1(n_76),
.B2(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_42),
.A2(n_50),
.B1(n_88),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_42),
.A2(n_50),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_50),
.B1(n_151),
.B2(n_182),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_42),
.A2(n_50),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_42),
.A2(n_50),
.B1(n_223),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_43),
.A2(n_128),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_43),
.A2(n_152),
.B1(n_181),
.B2(n_261),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_43)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_44),
.B(n_246),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_47),
.A2(n_49),
.B(n_188),
.Y(n_225)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_50),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_52),
.B(n_63),
.Y(n_189)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_65),
.B2(n_68),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_60),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_60),
.A2(n_68),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_60),
.A2(n_68),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_66),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_74),
.B1(n_100),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_64),
.A2(n_100),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_64),
.A2(n_100),
.B1(n_172),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_64),
.A2(n_169),
.B(n_258),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_89),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_79),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_81),
.B1(n_89),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_82),
.A2(n_84),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_82),
.A2(n_84),
.B1(n_177),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_82),
.A2(n_84),
.B1(n_148),
.B2(n_178),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_82),
.A2(n_84),
.B1(n_191),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_82),
.A2(n_84),
.B1(n_188),
.B2(n_244),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_82),
.A2(n_84),
.B1(n_237),
.B2(n_244),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_124),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_83),
.A2(n_146),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_134),
.B(n_307),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_107),
.B(n_110),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_118),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_131),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_120),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_292)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_160),
.B(n_306),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_158),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_137),
.B(n_158),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_138),
.B(n_141),
.Y(n_304)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_142),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.C(n_155),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_143),
.A2(n_144),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_145),
.B(n_149),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_153),
.B(n_155),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_154),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_156),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_301),
.B(n_305),
.Y(n_160)
);

OAI221xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_288),
.B1(n_299),
.B2(n_300),
.C(n_309),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_272),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_215),
.B(n_271),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_192),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_165),
.B(n_192),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.C(n_183),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_166),
.B(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_174),
.C(n_176),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_175),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_179),
.A2(n_183),
.B1(n_184),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_185),
.A2(n_186),
.B1(n_190),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_206),
.B2(n_214),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_193),
.B(n_207),
.C(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_195),
.B(n_201),
.C(n_205),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_208),
.B(n_211),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_265),
.B(n_270),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_253),
.B(n_264),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_233),
.B(n_252),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_226),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_219),
.B(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_241),
.B(n_251),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_239),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_247),
.B(n_250),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_274),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_283),
.C(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_296),
.B2(n_297),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_292),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_297),
.C(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);


endmodule