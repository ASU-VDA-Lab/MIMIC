module fake_jpeg_16890_n_145 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_22),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_47),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_28),
.B1(n_22),
.B2(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_24),
.B1(n_68),
.B2(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_0),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_32),
.C(n_43),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_42),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_43),
.A3(n_29),
.B1(n_53),
.B2(n_19),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_0),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_61),
.B(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_60),
.B1(n_67),
.B2(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_12),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_96),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_102),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_76),
.B(n_87),
.C(n_73),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_100),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_88),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_111),
.B(n_98),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_81),
.B1(n_77),
.B2(n_82),
.C(n_29),
.Y(n_106)
);

OAI321xp33_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_91),
.A3(n_101),
.B1(n_98),
.B2(n_15),
.C(n_20),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_76),
.B(n_23),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_5),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_117),
.B1(n_119),
.B2(n_122),
.Y(n_128)
);

OAI322xp33_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_108),
.A3(n_15),
.B1(n_23),
.B2(n_18),
.C1(n_20),
.C2(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_121),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_91),
.C(n_85),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.C(n_114),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_96),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_113),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_126),
.C(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_119),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_129),
.A2(n_133),
.B(n_128),
.C(n_124),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_127),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_108),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_123),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_136),
.B(n_130),
.C(n_131),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_139),
.B(n_10),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_110),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_6),
.B(n_7),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_12),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_142),
.B(n_85),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_50),
.C(n_69),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_70),
.Y(n_145)
);


endmodule