module fake_jpeg_2787_n_524 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_524);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_524;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_12),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_60),
.Y(n_151)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_64),
.Y(n_132)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_66),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx2_ASAP7_75t_R g133 ( 
.A(n_80),
.Y(n_133)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_11),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_88),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_87),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_15),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_19),
.B(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_91),
.B(n_93),
.Y(n_170)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_15),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_52),
.Y(n_171)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

BUFx4f_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_105),
.Y(n_201)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_118),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_31),
.Y(n_114)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_119),
.B(n_51),
.Y(n_159)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_34),
.B1(n_40),
.B2(n_36),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_124),
.A2(n_147),
.B1(n_156),
.B2(n_9),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_93),
.B(n_19),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_129),
.B(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_153),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_76),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_72),
.A2(n_18),
.B1(n_66),
.B2(n_105),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_150),
.A2(n_175),
.B1(n_181),
.B2(n_194),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_46),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_46),
.B1(n_45),
.B2(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_159),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_45),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_56),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_177),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_60),
.A2(n_56),
.B1(n_29),
.B2(n_37),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_87),
.B(n_52),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_108),
.A2(n_37),
.B1(n_29),
.B2(n_35),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_96),
.A2(n_35),
.B(n_33),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_183),
.A2(n_142),
.B(n_125),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_59),
.A2(n_33),
.B1(n_28),
.B2(n_51),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_187),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_65),
.B(n_28),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_78),
.B(n_15),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_61),
.B(n_0),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_193),
.B(n_185),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_114),
.A2(n_92),
.B1(n_99),
.B2(n_110),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_107),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_R g211 ( 
.A(n_196),
.B(n_51),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_62),
.A2(n_51),
.B1(n_1),
.B2(n_3),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_198),
.A2(n_69),
.B1(n_104),
.B2(n_83),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_204),
.A2(n_217),
.B1(n_240),
.B2(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_106),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_205),
.B(n_216),
.Y(n_275)
);

OR2x2_ASAP7_75t_SL g206 ( 
.A(n_128),
.B(n_80),
.Y(n_206)
);

NOR2x1_ASAP7_75t_R g284 ( 
.A(n_206),
.B(n_224),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_132),
.B(n_146),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_211),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_77),
.B1(n_74),
.B2(n_67),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_126),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_210),
.B(n_212),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_170),
.B(n_102),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_214),
.B(n_256),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_0),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_5),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_220),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_140),
.Y(n_219)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_5),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_137),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

NAND2x1_ASAP7_75t_L g228 ( 
.A(n_158),
.B(n_6),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_248),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_231),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_303)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_132),
.B(n_6),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_128),
.A2(n_8),
.B1(n_9),
.B2(n_177),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_163),
.A2(n_8),
.B1(n_138),
.B2(n_179),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_192),
.A2(n_190),
.B1(n_180),
.B2(n_176),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_242),
.A2(n_245),
.B1(n_265),
.B2(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

INVx11_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g248 ( 
.A(n_133),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_171),
.A2(n_144),
.B1(n_154),
.B2(n_143),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_258),
.Y(n_288)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_138),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_250),
.B(n_251),
.Y(n_307)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_255),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g254 ( 
.A(n_151),
.Y(n_254)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_170),
.B(n_135),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_155),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_259),
.Y(n_294)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_127),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_260),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_194),
.A2(n_198),
.B1(n_181),
.B2(n_175),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_157),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_262),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_166),
.A2(n_150),
.B1(n_188),
.B2(n_134),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_122),
.A2(n_188),
.B1(n_169),
.B2(n_134),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_136),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_186),
.A2(n_135),
.B1(n_197),
.B2(n_123),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_122),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_125),
.A2(n_18),
.B1(n_124),
.B2(n_55),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_169),
.B(n_184),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_264),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_184),
.B(n_230),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_289),
.A2(n_254),
.B(n_223),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_291),
.B(n_293),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_217),
.A2(n_253),
.B1(n_213),
.B2(n_211),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_292),
.A2(n_299),
.B1(n_305),
.B2(n_311),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_253),
.A2(n_221),
.B(n_230),
.C(n_261),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_241),
.B(n_257),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_229),
.A2(n_207),
.B1(n_249),
.B2(n_240),
.Y(n_299)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_224),
.A2(n_208),
.B1(n_221),
.B2(n_206),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_224),
.B(n_234),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_320),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_208),
.A2(n_221),
.B1(n_263),
.B2(n_231),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_215),
.B(n_228),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_314),
.B(n_248),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_234),
.B(n_227),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_221),
.B1(n_259),
.B2(n_252),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_321),
.A2(n_326),
.B1(n_329),
.B2(n_294),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_323),
.A2(n_336),
.B(n_350),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_296),
.A2(n_241),
.B(n_245),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_324),
.A2(n_300),
.B(n_308),
.Y(n_374)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_303),
.A2(n_250),
.B1(n_238),
.B2(n_226),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_296),
.A2(n_288),
.B1(n_271),
.B2(n_289),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_343),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_225),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_337),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_338),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_235),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_342),
.Y(n_361)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

BUFx24_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_273),
.B(n_236),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_232),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_347),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_237),
.B1(n_260),
.B2(n_265),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_345),
.A2(n_348),
.B1(n_349),
.B2(n_301),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_295),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_271),
.B1(n_291),
.B2(n_292),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_286),
.A2(n_312),
.B1(n_288),
.B2(n_298),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_312),
.B(n_283),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_278),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_354),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_297),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_283),
.A2(n_309),
.B1(n_282),
.B2(n_284),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_353),
.A2(n_316),
.B1(n_279),
.B2(n_276),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_312),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_294),
.A2(n_276),
.B1(n_308),
.B2(n_274),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_279),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_339),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_359),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_384),
.B1(n_389),
.B2(n_336),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_317),
.C(n_310),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_369),
.C(n_373),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_331),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_317),
.C(n_310),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_374),
.A2(n_344),
.B(n_351),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_359),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_378),
.Y(n_393)
);

OA22x2_ASAP7_75t_L g379 ( 
.A1(n_349),
.A2(n_345),
.B1(n_348),
.B2(n_322),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_380),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_346),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_381),
.B(n_358),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_321),
.B1(n_326),
.B2(n_342),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_322),
.A2(n_281),
.B1(n_301),
.B2(n_285),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_392),
.A2(n_361),
.B1(n_385),
.B2(n_377),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_384),
.A2(n_323),
.B1(n_347),
.B2(n_324),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_395),
.B1(n_386),
.B2(n_389),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_382),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_376),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_367),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_405),
.Y(n_428)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_367),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_399),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_350),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_408),
.Y(n_421)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_371),
.A2(n_329),
.B(n_337),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_330),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_343),
.C(n_340),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_418),
.C(n_391),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_325),
.B(n_328),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_412),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_379),
.A2(n_358),
.B1(n_338),
.B2(n_281),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_378),
.B1(n_363),
.B2(n_388),
.Y(n_442)
);

OAI31xp33_ASAP7_75t_SL g414 ( 
.A1(n_379),
.A2(n_341),
.A3(n_319),
.B(n_318),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_390),
.Y(n_441)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_364),
.A2(n_290),
.B(n_313),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_373),
.Y(n_426)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_417),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_381),
.B(n_290),
.C(n_313),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_419),
.A2(n_424),
.B1(n_425),
.B2(n_436),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_420),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_402),
.A2(n_364),
.B1(n_379),
.B2(n_360),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_402),
.A2(n_379),
.B1(n_361),
.B2(n_385),
.Y(n_425)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_442),
.B1(n_410),
.B2(n_416),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_437),
.C(n_406),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_366),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_404),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_413),
.A2(n_372),
.B1(n_383),
.B2(n_366),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_380),
.C(n_363),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_393),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_439),
.B(n_411),
.Y(n_446)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_445),
.A2(n_458),
.B1(n_424),
.B2(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_454),
.C(n_459),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_433),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_451),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_456),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_433),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_453),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_409),
.C(n_408),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_455),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_405),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_457),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_419),
.A2(n_394),
.B1(n_397),
.B2(n_392),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_418),
.C(n_398),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_417),
.C(n_403),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_460),
.B(n_461),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_428),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_399),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_428),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_450),
.A2(n_453),
.B1(n_425),
.B2(n_445),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_463),
.A2(n_458),
.B1(n_452),
.B2(n_440),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_426),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_447),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_422),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_468),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_452),
.B1(n_441),
.B2(n_436),
.Y(n_482)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_476),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_477),
.B(n_456),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_481),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_479),
.A2(n_483),
.B1(n_470),
.B2(n_422),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_438),
.Y(n_480)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_480),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_482),
.A2(n_449),
.B1(n_469),
.B2(n_457),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_463),
.A2(n_442),
.B1(n_422),
.B2(n_444),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_487),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_472),
.B(n_468),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_486),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_459),
.C(n_444),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_464),
.C(n_477),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_478),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_388),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_497),
.Y(n_503)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

OAI321xp33_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_465),
.A3(n_474),
.B1(n_473),
.B2(n_431),
.C(n_475),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_498),
.B(n_414),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_469),
.B(n_462),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_499),
.B(n_429),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_479),
.C(n_483),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_502),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_493),
.A2(n_482),
.B(n_485),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_505),
.B(n_507),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_481),
.C(n_432),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_494),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_512),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_510),
.C(n_434),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_375),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_495),
.Y(n_513)
);

OAI21x1_ASAP7_75t_SL g517 ( 
.A1(n_513),
.A2(n_407),
.B(n_390),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_509),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_514),
.A2(n_515),
.B(n_517),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_387),
.C(n_375),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_387),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_518),
.C(n_370),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_375),
.C(n_341),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_341),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_319),
.B(n_272),
.Y(n_524)
);


endmodule