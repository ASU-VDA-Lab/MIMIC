module fake_jpeg_141_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_8),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_17),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_70),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_77),
.B1(n_68),
.B2(n_79),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_94),
.B1(n_62),
.B2(n_61),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_59),
.B1(n_68),
.B2(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_54),
.B1(n_65),
.B2(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_70),
.B1(n_60),
.B2(n_54),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_104),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_65),
.B1(n_50),
.B2(n_55),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_86),
.A3(n_63),
.B1(n_57),
.B2(n_90),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_0),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_50),
.B(n_55),
.C(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_72),
.B1(n_71),
.B2(n_66),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_110),
.Y(n_116)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_3),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_61),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_100),
.B(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_67),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_125),
.B1(n_119),
.B2(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_0),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_124),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_128),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_7),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_8),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_24),
.C(n_48),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_97),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_138),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_140),
.Y(n_170)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_142),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_9),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_11),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_12),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_28),
.B1(n_47),
.B2(n_16),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_150),
.A2(n_152),
.B(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_155),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_13),
.B(n_15),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_15),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_49),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_150),
.B1(n_146),
.B2(n_137),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_134),
.C(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_131),
.C(n_20),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

AO221x1_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_168),
.B1(n_160),
.B2(n_163),
.C(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_18),
.C(n_21),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_46),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_181),
.B1(n_182),
.B2(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_179),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_22),
.C(n_23),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_25),
.C(n_27),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_165),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_30),
.B(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_35),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_178),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_189),
.B1(n_182),
.B2(n_172),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_157),
.B1(n_168),
.B2(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_192),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_183),
.B(n_189),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_186),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_196),
.C(n_192),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_39),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_42),
.Y(n_201)
);


endmodule