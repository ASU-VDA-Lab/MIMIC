module real_aes_4612_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_1004;
wire n_580;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_994;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_992;
wire n_774;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_1025;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_973;
wire n_310;
wire n_725;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_1017;
wire n_1013;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_997;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_649;
wire n_293;
wire n_397;
wire n_358;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_968;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_0), .A2(n_154), .B1(n_433), .B2(n_465), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_1), .A2(n_145), .B1(n_501), .B2(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g416 ( .A(n_2), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_3), .A2(n_97), .B1(n_327), .B2(n_334), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_4), .A2(n_7), .B1(n_442), .B2(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g679 ( .A(n_5), .Y(n_679) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_6), .Y(n_741) );
AND2x4_ASAP7_75t_L g753 ( .A(n_6), .B(n_274), .Y(n_753) );
AND2x4_ASAP7_75t_L g758 ( .A(n_6), .B(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_8), .A2(n_54), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_9), .A2(n_184), .B1(n_430), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_10), .A2(n_163), .B1(n_316), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_11), .A2(n_257), .B1(n_495), .B2(n_501), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_12), .A2(n_68), .B1(n_461), .B2(n_462), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_13), .A2(n_141), .B1(n_462), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_14), .A2(n_106), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_15), .A2(n_117), .B1(n_750), .B2(n_754), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_16), .A2(n_36), .B1(n_497), .B2(n_498), .Y(n_631) );
INVx1_ASAP7_75t_L g587 ( .A(n_17), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_18), .A2(n_101), .B1(n_337), .B2(n_341), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_19), .A2(n_20), .B1(n_369), .B2(n_529), .Y(n_561) );
AO22x1_ASAP7_75t_L g456 ( .A1(n_21), .A2(n_128), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_22), .A2(n_103), .B1(n_430), .B2(n_431), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_23), .A2(n_200), .B1(n_327), .B2(n_334), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_24), .A2(n_120), .B1(n_576), .B2(n_613), .Y(n_612) );
XNOR2x1_ASAP7_75t_L g694 ( .A(n_25), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g1015 ( .A(n_26), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_27), .A2(n_90), .B1(n_488), .B2(n_509), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_28), .A2(n_253), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI211x1_ASAP7_75t_L g1008 ( .A1(n_29), .A2(n_1009), .B(n_1011), .C(n_1018), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_30), .A2(n_86), .B1(n_437), .B2(n_439), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_31), .A2(n_192), .B1(n_411), .B2(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g733 ( .A(n_32), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_33), .A2(n_150), .B1(n_408), .B2(n_981), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_34), .A2(n_135), .B1(n_470), .B2(n_1017), .Y(n_1016) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_35), .A2(n_240), .B1(n_418), .B2(n_642), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_37), .A2(n_254), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_38), .A2(n_278), .B1(n_576), .B2(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_39), .B(n_477), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_40), .B(n_582), .Y(n_730) );
INVx1_ASAP7_75t_SL g289 ( .A(n_41), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_42), .A2(n_111), .B1(n_773), .B2(n_775), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_43), .A2(n_183), .B1(n_411), .B2(n_643), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_44), .A2(n_175), .B1(n_348), .B2(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_45), .B(n_477), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_46), .A2(n_88), .B1(n_442), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_47), .A2(n_279), .B1(n_411), .B2(n_470), .Y(n_727) );
INVx1_ASAP7_75t_L g313 ( .A(n_48), .Y(n_313) );
INVxp67_ASAP7_75t_L g388 ( .A(n_48), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_48), .B(n_218), .Y(n_394) );
INVx1_ASAP7_75t_L g420 ( .A(n_49), .Y(n_420) );
INVx1_ASAP7_75t_L g474 ( .A(n_50), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_51), .A2(n_83), .B1(n_457), .B2(n_464), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_52), .A2(n_204), .B1(n_777), .B2(n_778), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_52), .A2(n_973), .B1(n_987), .B2(n_988), .Y(n_972) );
INVxp67_ASAP7_75t_L g988 ( .A(n_52), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_52), .A2(n_995), .B1(n_997), .B2(n_1023), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_53), .A2(n_263), .B1(n_784), .B2(n_805), .Y(n_852) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_55), .B(n_298), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_56), .A2(n_148), .B1(n_488), .B2(n_489), .Y(n_708) );
INVx1_ASAP7_75t_L g406 ( .A(n_57), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_58), .A2(n_114), .B1(n_604), .B2(n_605), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_59), .A2(n_167), .B1(n_494), .B2(n_551), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_60), .A2(n_65), .B1(n_293), .B2(n_316), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_61), .A2(n_261), .B1(n_389), .B2(n_506), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_62), .A2(n_170), .B1(n_455), .B2(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_63), .A2(n_186), .B1(n_442), .B2(n_443), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_64), .A2(n_130), .B1(n_750), .B2(n_754), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_66), .A2(n_277), .B1(n_346), .B2(n_348), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_67), .A2(n_168), .B1(n_458), .B2(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g559 ( .A(n_69), .Y(n_559) );
INVx2_ASAP7_75t_L g739 ( .A(n_70), .Y(n_739) );
INVx1_ASAP7_75t_L g752 ( .A(n_71), .Y(n_752) );
AND2x4_ASAP7_75t_L g755 ( .A(n_71), .B(n_739), .Y(n_755) );
INVx1_ASAP7_75t_SL g774 ( .A(n_71), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_72), .A2(n_207), .B1(n_418), .B2(n_729), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_73), .A2(n_266), .B1(n_430), .B2(n_431), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_74), .A2(n_133), .B1(n_491), .B2(n_492), .Y(n_629) );
INVx1_ASAP7_75t_L g1022 ( .A(n_75), .Y(n_1022) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_76), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g699 ( .A(n_77), .Y(n_699) );
INVx1_ASAP7_75t_L g413 ( .A(n_78), .Y(n_413) );
OAI22xp33_ASAP7_75t_SL g997 ( .A1(n_79), .A2(n_998), .B1(n_999), .B2(n_1000), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_79), .Y(n_998) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_80), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_81), .A2(n_109), .B1(n_433), .B2(n_465), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_82), .A2(n_179), .B1(n_777), .B2(n_778), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_84), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g802 ( .A(n_85), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_87), .A2(n_157), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_89), .A2(n_524), .B(n_526), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_91), .A2(n_276), .B1(n_773), .B2(n_775), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_92), .A2(n_199), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_93), .A2(n_181), .B1(n_506), .B2(n_509), .C(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_94), .A2(n_275), .B1(n_379), .B2(n_411), .Y(n_560) );
INVx1_ASAP7_75t_L g299 ( .A(n_95), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_95), .B(n_216), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_96), .A2(n_260), .B1(n_379), .B2(n_389), .Y(n_378) );
INVx1_ASAP7_75t_L g409 ( .A(n_98), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_99), .A2(n_245), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_100), .A2(n_107), .B1(n_773), .B2(n_775), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_102), .A2(n_208), .B1(n_461), .B2(n_462), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_104), .A2(n_152), .B1(n_431), .B2(n_455), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_105), .A2(n_172), .B1(n_379), .B2(n_411), .Y(n_531) );
XOR2xp5_ASAP7_75t_L g591 ( .A(n_108), .B(n_592), .Y(n_591) );
XNOR2x2_ASAP7_75t_L g615 ( .A(n_108), .B(n_592), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_110), .A2(n_224), .B1(n_430), .B2(n_431), .Y(n_725) );
INVx1_ASAP7_75t_L g546 ( .A(n_112), .Y(n_546) );
INVx1_ASAP7_75t_L g364 ( .A(n_113), .Y(n_364) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_115), .A2(n_506), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g511 ( .A(n_116), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_118), .A2(n_144), .B1(n_346), .B2(n_1004), .Y(n_1003) );
AOI21xp33_ASAP7_75t_L g508 ( .A1(n_119), .A2(n_509), .B(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_121), .A2(n_269), .B1(n_494), .B2(n_495), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_122), .A2(n_195), .B1(n_554), .B2(n_555), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_123), .A2(n_235), .B1(n_431), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_124), .A2(n_147), .B1(n_346), .B2(n_465), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_125), .A2(n_221), .B1(n_777), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_126), .A2(n_169), .B1(n_408), .B2(n_418), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_127), .A2(n_220), .B1(n_461), .B2(n_462), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_129), .A2(n_252), .B1(n_293), .B2(n_316), .Y(n_292) );
INVxp33_ASAP7_75t_SL g808 ( .A(n_131), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_132), .A2(n_203), .B1(n_369), .B2(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_134), .A2(n_206), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_136), .A2(n_143), .B1(n_337), .B2(n_341), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_137), .A2(n_191), .B1(n_431), .B2(n_455), .Y(n_985) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_138), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_138), .A2(n_190), .B1(n_757), .B2(n_760), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_139), .A2(n_162), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g527 ( .A(n_140), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_142), .A2(n_153), .B1(n_554), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_146), .A2(n_165), .B1(n_355), .B2(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_149), .A2(n_265), .B1(n_337), .B2(n_341), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_151), .B(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_155), .A2(n_231), .B1(n_430), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_156), .A2(n_237), .B1(n_379), .B2(n_411), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_158), .A2(n_188), .B1(n_433), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_159), .A2(n_273), .B1(n_433), .B2(n_537), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_160), .A2(n_264), .B1(n_489), .B2(n_494), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_161), .A2(n_250), .B1(n_684), .B2(n_686), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_164), .A2(n_202), .B1(n_491), .B2(n_492), .Y(n_709) );
XOR2xp5_ASAP7_75t_L g620 ( .A(n_166), .B(n_621), .Y(n_620) );
XOR2xp5_ASAP7_75t_L g662 ( .A(n_166), .B(n_621), .Y(n_662) );
INVx1_ASAP7_75t_L g806 ( .A(n_171), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_173), .A2(n_258), .B1(n_369), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_174), .A2(n_213), .B1(n_422), .B2(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_176), .B(n_605), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_177), .A2(n_255), .B1(n_316), .B2(n_574), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_178), .A2(n_242), .B1(n_461), .B2(n_462), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_180), .A2(n_229), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_182), .A2(n_194), .B1(n_424), .B2(n_507), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_185), .A2(n_355), .B(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_187), .A2(n_234), .B1(n_293), .B2(n_316), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_189), .A2(n_236), .B1(n_504), .B2(n_509), .C(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_193), .A2(n_198), .B1(n_415), .B2(n_418), .Y(n_468) );
INVx1_ASAP7_75t_L g655 ( .A(n_196), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_197), .A2(n_267), .B1(n_461), .B2(n_462), .Y(n_460) );
OA22x2_ASAP7_75t_L g303 ( .A1(n_201), .A2(n_218), .B1(n_298), .B2(n_302), .Y(n_303) );
INVx1_ASAP7_75t_L g322 ( .A(n_201), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_205), .A2(n_271), .B1(n_757), .B2(n_760), .Y(n_767) );
AO22x2_ASAP7_75t_L g400 ( .A1(n_209), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_209), .Y(n_401) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_210), .B(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_211), .A2(n_249), .B1(n_316), .B2(n_457), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_212), .A2(n_226), .B1(n_327), .B2(n_334), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_214), .A2(n_259), .B1(n_530), .B2(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g367 ( .A(n_215), .Y(n_367) );
INVx1_ASAP7_75t_L g315 ( .A(n_216), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_216), .B(n_320), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_217), .A2(n_243), .B1(n_506), .B2(n_507), .Y(n_505) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_218), .A2(n_239), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g851 ( .A(n_219), .Y(n_851) );
XNOR2x2_ASAP7_75t_SL g484 ( .A(n_222), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g668 ( .A(n_223), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_225), .B(n_415), .Y(n_623) );
INVx1_ASAP7_75t_L g717 ( .A(n_227), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_227), .A2(n_244), .B1(n_773), .B2(n_775), .Y(n_780) );
AOI21xp33_ASAP7_75t_L g977 ( .A1(n_228), .A2(n_529), .B(n_978), .Y(n_977) );
OAI21x1_ASAP7_75t_L g450 ( .A1(n_230), .A2(n_451), .B(n_478), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_230), .B(n_454), .Y(n_481) );
INVx1_ASAP7_75t_L g1012 ( .A(n_232), .Y(n_1012) );
INVx1_ASAP7_75t_L g353 ( .A(n_233), .Y(n_353) );
INVx1_ASAP7_75t_L g1020 ( .A(n_238), .Y(n_1020) );
INVx1_ASAP7_75t_L g301 ( .A(n_239), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_239), .B(n_268), .Y(n_395) );
INVx1_ASAP7_75t_L g358 ( .A(n_241), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_246), .A2(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g373 ( .A(n_247), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_248), .A2(n_262), .B1(n_701), .B2(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g979 ( .A(n_251), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_256), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_268), .B(n_308), .Y(n_307) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_270), .A2(n_355), .B(n_473), .Y(n_472) );
INVxp33_ASAP7_75t_L g800 ( .A(n_272), .Y(n_800) );
INVx1_ASAP7_75t_L g759 ( .A(n_274), .Y(n_759) );
INVx1_ASAP7_75t_L g519 ( .A(n_280), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_280), .B(n_538), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_742), .B(n_743), .Y(n_281) );
AOI21xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_616), .B(n_734), .Y(n_282) );
OR2x2_ASAP7_75t_L g742 ( .A(n_283), .B(n_616), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_514), .B2(n_515), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B1(n_448), .B2(n_513), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_398), .B1(n_445), .B2(n_446), .Y(n_287) );
INVx2_ASAP7_75t_L g445 ( .A(n_288), .Y(n_445) );
XNOR2x1_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_351), .Y(n_290) );
AND4x1_ASAP7_75t_L g291 ( .A(n_292), .B(n_326), .C(n_336), .D(n_345), .Y(n_291) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_294), .Y(n_442) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_294), .Y(n_457) );
BUFx12f_ASAP7_75t_L g574 ( .A(n_294), .Y(n_574) );
BUFx3_ASAP7_75t_L g688 ( .A(n_294), .Y(n_688) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_304), .Y(n_294) );
AND2x2_ASAP7_75t_L g347 ( .A(n_295), .B(n_332), .Y(n_347) );
AND2x2_ASAP7_75t_L g362 ( .A(n_295), .B(n_339), .Y(n_362) );
AND2x2_ASAP7_75t_L g377 ( .A(n_295), .B(n_343), .Y(n_377) );
AND2x2_ASAP7_75t_L g434 ( .A(n_295), .B(n_332), .Y(n_434) );
AND2x4_ASAP7_75t_L g488 ( .A(n_295), .B(n_332), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_295), .B(n_325), .Y(n_489) );
AND2x4_ASAP7_75t_L g501 ( .A(n_295), .B(n_339), .Y(n_501) );
AND2x2_ASAP7_75t_L g506 ( .A(n_295), .B(n_343), .Y(n_506) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_303), .Y(n_295) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
NAND2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g302 ( .A(n_298), .Y(n_302) );
INVx3_ASAP7_75t_L g308 ( .A(n_298), .Y(n_308) );
NAND2xp33_ASAP7_75t_L g314 ( .A(n_298), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_298), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_299), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g387 ( .A1(n_301), .A2(n_324), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
AND2x2_ASAP7_75t_L g357 ( .A(n_303), .B(n_330), .Y(n_357) );
AND2x2_ASAP7_75t_L g386 ( .A(n_303), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g495 ( .A(n_304), .B(n_329), .Y(n_495) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g325 ( .A(n_305), .Y(n_325) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_310), .Y(n_305) );
AND2x4_ASAP7_75t_L g332 ( .A(n_306), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g339 ( .A(n_306), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
AND2x2_ASAP7_75t_L g382 ( .A(n_306), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_308), .B(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g320 ( .A(n_308), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_309), .B(n_319), .C(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g340 ( .A(n_311), .Y(n_340) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
BUFx12f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx6_ASAP7_75t_L g444 ( .A(n_317), .Y(n_444) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_325), .Y(n_317) );
AND2x4_ASAP7_75t_L g350 ( .A(n_318), .B(n_332), .Y(n_350) );
AND2x4_ASAP7_75t_L g371 ( .A(n_318), .B(n_343), .Y(n_371) );
AND2x4_ASAP7_75t_L g497 ( .A(n_318), .B(n_332), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_318), .B(n_325), .Y(n_498) );
AND2x4_ASAP7_75t_L g507 ( .A(n_318), .B(n_343), .Y(n_507) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x4_ASAP7_75t_L g335 ( .A(n_325), .B(n_329), .Y(n_335) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_328), .Y(n_430) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_328), .Y(n_455) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AND2x4_ASAP7_75t_L g338 ( .A(n_329), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g342 ( .A(n_329), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g491 ( .A(n_329), .B(n_339), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_329), .B(n_343), .Y(n_492) );
AND2x4_ASAP7_75t_L g494 ( .A(n_329), .B(n_332), .Y(n_494) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_335), .Y(n_431) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_335), .Y(n_551) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_335), .Y(n_571) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g438 ( .A(n_338), .Y(n_438) );
BUFx12f_ASAP7_75t_L g461 ( .A(n_338), .Y(n_461) );
AND2x4_ASAP7_75t_L g356 ( .A(n_339), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g509 ( .A(n_339), .B(n_357), .Y(n_509) );
AND2x4_ASAP7_75t_L g343 ( .A(n_340), .B(n_344), .Y(n_343) );
BUFx5_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g440 ( .A(n_342), .Y(n_440) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_342), .Y(n_462) );
BUFx3_ASAP7_75t_L g555 ( .A(n_342), .Y(n_555) );
AND2x4_ASAP7_75t_L g366 ( .A(n_343), .B(n_357), .Y(n_366) );
AND2x2_ASAP7_75t_L g504 ( .A(n_343), .B(n_357), .Y(n_504) );
BUFx8_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_347), .Y(n_576) );
INVx4_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx4_ASAP7_75t_L g465 ( .A(n_349), .Y(n_465) );
INVx1_ASAP7_75t_L g537 ( .A(n_349), .Y(n_537) );
INVx2_ASAP7_75t_L g577 ( .A(n_349), .Y(n_577) );
INVx4_ASAP7_75t_L g613 ( .A(n_349), .Y(n_613) );
INVx2_ASAP7_75t_SL g723 ( .A(n_349), .Y(n_723) );
INVx1_ASAP7_75t_L g1004 ( .A(n_349), .Y(n_1004) );
INVx8_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_363), .C(n_372), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_358), .B2(n_359), .Y(n_352) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g408 ( .A(n_356), .Y(n_408) );
INVx1_ASAP7_75t_L g525 ( .A(n_356), .Y(n_525) );
BUFx3_ASAP7_75t_L g729 ( .A(n_356), .Y(n_729) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_361), .Y(n_600) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
BUFx3_ASAP7_75t_L g642 ( .A(n_362), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_367), .B2(n_368), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g1014 ( .A1(n_365), .A2(n_1015), .B(n_1016), .Y(n_1014) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_366), .Y(n_529) );
BUFx3_ASAP7_75t_L g582 ( .A(n_366), .Y(n_582) );
BUFx8_ASAP7_75t_SL g602 ( .A(n_366), .Y(n_602) );
INVx2_ASAP7_75t_L g646 ( .A(n_366), .Y(n_646) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g530 ( .A(n_370), .Y(n_530) );
INVx2_ASAP7_75t_L g702 ( .A(n_370), .Y(n_702) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g677 ( .A(n_374), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g1011 ( .A1(n_374), .A2(n_1012), .B(n_1013), .Y(n_1011) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g477 ( .A(n_376), .Y(n_477) );
INVx3_ASAP7_75t_SL g580 ( .A(n_376), .Y(n_580) );
INVx2_ASAP7_75t_L g701 ( .A(n_376), .Y(n_701) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
INVx2_ASAP7_75t_L g597 ( .A(n_377), .Y(n_597) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g604 ( .A(n_380), .Y(n_604) );
INVx5_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_381), .Y(n_470) );
BUFx2_ASAP7_75t_L g643 ( .A(n_381), .Y(n_643) );
BUFx2_ASAP7_75t_L g981 ( .A(n_381), .Y(n_981) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
AND2x2_ASAP7_75t_L g424 ( .A(n_382), .B(n_386), .Y(n_424) );
AND2x4_ASAP7_75t_L g502 ( .A(n_382), .B(n_386), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g392 ( .A(n_384), .Y(n_392) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_390), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_390), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g589 ( .A(n_390), .Y(n_589) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g607 ( .A(n_391), .Y(n_607) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_396), .Y(n_391) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_393), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_427), .Y(n_403) );
NOR3xp33_ASAP7_75t_SL g404 ( .A(n_405), .B(n_412), .C(n_419), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_409), .B2(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g674 ( .A(n_408), .Y(n_674) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx3_ASAP7_75t_L g675 ( .A(n_411), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_416), .B2(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g672 ( .A(n_414), .Y(n_672) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_423), .Y(n_419) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_435), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g685 ( .A(n_430), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_431), .Y(n_686) );
BUFx4f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_434), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_441), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g554 ( .A(n_438), .Y(n_554) );
INVx1_ASAP7_75t_L g569 ( .A(n_438), .Y(n_569) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx5_ASAP7_75t_L g458 ( .A(n_444), .Y(n_458) );
INVx2_ASAP7_75t_L g535 ( .A(n_444), .Y(n_535) );
INVx2_ASAP7_75t_L g721 ( .A(n_444), .Y(n_721) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
OA22x2_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_482), .B1(n_483), .B2(n_512), .Y(n_448) );
INVx2_ASAP7_75t_L g512 ( .A(n_449), .Y(n_512) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_466), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .C(n_459), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_456), .B(n_471), .C(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_459), .B(n_467), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_463), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_SL g680 ( .A(n_470), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_475), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_475), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g649 ( .A(n_475), .Y(n_649) );
NOR2xp67_ASAP7_75t_SL g698 ( .A(n_475), .B(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_475), .B(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_475), .B(n_979), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_499), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .C(n_493), .D(n_496), .Y(n_486) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_497), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .C(n_505), .D(n_508), .Y(n_499) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
XOR2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_562), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_544), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI21x1_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_541), .Y(n_518) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_521), .B(n_542), .C(n_543), .Y(n_541) );
AND4x1_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .C(n_528), .D(n_531), .Y(n_521) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g1019 ( .A(n_530), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_538), .Y(n_532) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_533), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
BUFx2_ASAP7_75t_L g689 ( .A(n_535), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
XNOR2x1_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_548), .B(n_556), .Y(n_547) );
NAND4xp25_ASAP7_75t_SL g548 ( .A(n_549), .B(n_550), .C(n_552), .D(n_553), .Y(n_548) );
BUFx2_ASAP7_75t_L g691 ( .A(n_555), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .C(n_561), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_591), .B1(n_614), .B2(n_615), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_564), .Y(n_614) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g565 ( .A(n_566), .B(n_590), .Y(n_565) );
NAND4xp75_ASAP7_75t_L g566 ( .A(n_567), .B(n_572), .C(n_578), .D(n_583), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_608), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_598), .C(n_601), .D(n_603), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx4_ASAP7_75t_L g1017 ( .A(n_606), .Y(n_1017) );
INVx4_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .C(n_611), .D(n_612), .Y(n_608) );
XNOR2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_664), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_632), .B1(n_656), .B2(n_663), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_627), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .C(n_625), .D(n_626), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .C(n_630), .D(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g663 ( .A(n_632), .Y(n_663) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
XOR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_655), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_650), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .C(n_647), .D(n_648), .Y(n_640) );
INVx2_ASAP7_75t_L g1021 ( .A(n_642), .Y(n_1021) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .C(n_653), .D(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
XOR2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_711), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_693), .B2(n_710), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
XNOR2x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_668), .A2(n_799), .B1(n_801), .B2(n_851), .C(n_852), .Y(n_850) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_682), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g670 ( .A(n_671), .B(n_673), .C(n_676), .Y(n_670) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B(n_681), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g682 ( .A(n_683), .B(n_687), .C(n_690), .D(n_692), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g710 ( .A(n_693), .Y(n_710) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_704), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .C(n_703), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .C(n_708), .D(n_709), .Y(n_704) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
XNOR2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_726), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .C(n_724), .D(n_725), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .C(n_730), .D(n_731), .Y(n_726) );
INVx2_ASAP7_75t_L g1010 ( .A(n_729), .Y(n_1010) );
BUFx10_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .C(n_741), .Y(n_736) );
AND2x2_ASAP7_75t_L g991 ( .A(n_737), .B(n_992), .Y(n_991) );
AND2x2_ASAP7_75t_L g996 ( .A(n_737), .B(n_993), .Y(n_996) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OA21x2_ASAP7_75t_L g1024 ( .A1(n_738), .A2(n_774), .B(n_1025), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g751 ( .A(n_739), .B(n_752), .Y(n_751) );
AND3x4_ASAP7_75t_L g773 ( .A(n_739), .B(n_758), .C(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_740), .B(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_741), .Y(n_993) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_969), .B1(n_971), .B2(n_989), .C(n_994), .Y(n_743) );
AOI211xp5_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_761), .B(n_838), .C(n_927), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g958 ( .A(n_745), .B(n_959), .C(n_960), .Y(n_958) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_746), .A2(n_869), .B1(n_875), .B2(n_894), .Y(n_868) );
AOI21xp33_ASAP7_75t_SL g911 ( .A1(n_746), .A2(n_875), .B(n_912), .Y(n_911) );
AND2x2_ASAP7_75t_L g916 ( .A(n_746), .B(n_917), .Y(n_916) );
BUFx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g867 ( .A(n_747), .Y(n_867) );
AND2x2_ASAP7_75t_L g914 ( .A(n_747), .B(n_796), .Y(n_914) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g874 ( .A(n_748), .Y(n_874) );
OR2x2_ASAP7_75t_L g921 ( .A(n_748), .B(n_812), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_756), .Y(n_748) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .Y(n_750) );
AND2x4_ASAP7_75t_L g757 ( .A(n_751), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g777 ( .A(n_751), .B(n_753), .Y(n_777) );
AND2x4_ASAP7_75t_L g805 ( .A(n_751), .B(n_753), .Y(n_805) );
AND2x2_ASAP7_75t_L g754 ( .A(n_753), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g778 ( .A(n_753), .B(n_755), .Y(n_778) );
AND2x4_ASAP7_75t_L g784 ( .A(n_753), .B(n_755), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_753), .Y(n_1025) );
AND2x4_ASAP7_75t_L g760 ( .A(n_755), .B(n_758), .Y(n_760) );
AND2x4_ASAP7_75t_L g775 ( .A(n_755), .B(n_758), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_755), .B(n_758), .Y(n_801) );
INVx3_ASAP7_75t_L g799 ( .A(n_757), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_786), .B(n_809), .C(n_815), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_763), .A2(n_794), .B1(n_811), .B2(n_843), .C(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_782), .Y(n_763) );
AND2x2_ASAP7_75t_L g816 ( .A(n_764), .B(n_817), .Y(n_816) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_769), .Y(n_764) );
INVx2_ASAP7_75t_L g789 ( .A(n_765), .Y(n_789) );
INVx2_ASAP7_75t_L g827 ( .A(n_765), .Y(n_827) );
INVx1_ASAP7_75t_L g832 ( .A(n_765), .Y(n_832) );
AND2x2_ASAP7_75t_L g835 ( .A(n_765), .B(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_765), .B(n_842), .Y(n_841) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_765), .Y(n_845) );
AND2x2_ASAP7_75t_L g877 ( .A(n_765), .B(n_793), .Y(n_877) );
AND2x2_ASAP7_75t_L g884 ( .A(n_765), .B(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_SL g893 ( .A(n_765), .B(n_857), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_765), .B(n_905), .Y(n_904) );
NAND2xp5_ASAP7_75t_SL g934 ( .A(n_765), .B(n_892), .Y(n_934) );
NAND2xp5_ASAP7_75t_SL g937 ( .A(n_765), .B(n_938), .Y(n_937) );
AND2x2_ASAP7_75t_L g961 ( .A(n_765), .B(n_797), .Y(n_961) );
INVx4_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g864 ( .A(n_766), .B(n_791), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_766), .B(n_796), .Y(n_949) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AOI21xp33_ASAP7_75t_L g887 ( .A1(n_769), .A2(n_888), .B(n_889), .Y(n_887) );
INVx3_ASAP7_75t_SL g892 ( .A(n_769), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_769), .B(n_791), .Y(n_897) );
OR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_779), .Y(n_769) );
AND2x2_ASAP7_75t_L g793 ( .A(n_770), .B(n_779), .Y(n_793) );
AND2x2_ASAP7_75t_L g842 ( .A(n_770), .B(n_817), .Y(n_842) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_L g820 ( .A(n_771), .B(n_779), .Y(n_820) );
AND2x2_ASAP7_75t_L g847 ( .A(n_771), .B(n_779), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_771), .B(n_782), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_771), .B(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_771), .B(n_817), .Y(n_939) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_776), .Y(n_771) );
AND2x2_ASAP7_75t_L g830 ( .A(n_779), .B(n_791), .Y(n_830) );
INVx1_ASAP7_75t_L g886 ( .A(n_779), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_779), .B(n_817), .Y(n_888) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_SL g792 ( .A(n_782), .Y(n_792) );
INVx1_ASAP7_75t_L g817 ( .A(n_782), .Y(n_817) );
OR2x2_ASAP7_75t_L g828 ( .A(n_782), .B(n_820), .Y(n_828) );
AND2x2_ASAP7_75t_L g885 ( .A(n_782), .B(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_782), .B(n_892), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_782), .B(n_877), .Y(n_901) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_785), .Y(n_782) );
INVx2_ASAP7_75t_L g807 ( .A(n_784), .Y(n_807) );
BUFx2_ASAP7_75t_L g970 ( .A(n_784), .Y(n_970) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AOI211xp5_ASAP7_75t_SL g839 ( .A1(n_787), .A2(n_794), .B(n_840), .C(n_843), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_794), .Y(n_787) );
NAND2xp67_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_789), .B(n_883), .Y(n_889) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_790), .A2(n_849), .B1(n_920), .B2(n_922), .C(n_924), .Y(n_919) );
O2A1O1Ixp33_ASAP7_75t_L g928 ( .A1(n_790), .A2(n_816), .B(n_916), .C(n_929), .Y(n_928) );
AND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
AND2x4_ASAP7_75t_L g818 ( .A(n_791), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g863 ( .A(n_793), .Y(n_863) );
AND2x2_ASAP7_75t_L g941 ( .A(n_793), .B(n_817), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_793), .B(n_968), .Y(n_967) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_794), .A2(n_891), .B(n_893), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_794), .B(n_921), .Y(n_935) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g822 ( .A(n_796), .B(n_812), .Y(n_822) );
AND2x2_ASAP7_75t_L g881 ( .A(n_796), .B(n_812), .Y(n_881) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OR2x2_ASAP7_75t_L g833 ( .A(n_797), .B(n_812), .Y(n_833) );
INVx1_ASAP7_75t_L g836 ( .A(n_797), .Y(n_836) );
AND2x2_ASAP7_75t_L g883 ( .A(n_797), .B(n_812), .Y(n_883) );
AND2x2_ASAP7_75t_L g954 ( .A(n_797), .B(n_946), .Y(n_954) );
OR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_803), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI322xp33_ASAP7_75t_L g838 ( .A1(n_809), .A2(n_839), .A3(n_848), .B1(n_853), .B2(n_866), .C1(n_868), .C2(n_911), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_809), .A2(n_932), .B1(n_933), .B2(n_935), .C(n_936), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_809), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_945) );
CKINVDCx14_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
CKINVDCx14_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_812), .Y(n_824) );
OR2x2_ASAP7_75t_L g900 ( .A(n_812), .B(n_874), .Y(n_900) );
AND2x2_ASAP7_75t_L g908 ( .A(n_812), .B(n_873), .Y(n_908) );
AND2x2_ASAP7_75t_L g946 ( .A(n_812), .B(n_874), .Y(n_946) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
O2A1O1Ixp33_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_818), .B(n_821), .C(n_823), .Y(n_815) );
AND2x2_ASAP7_75t_L g846 ( .A(n_817), .B(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g905 ( .A(n_817), .B(n_886), .Y(n_905) );
NOR2x1_ASAP7_75t_R g933 ( .A(n_817), .B(n_934), .Y(n_933) );
AND2x2_ASAP7_75t_L g879 ( .A(n_818), .B(n_827), .Y(n_879) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_820), .B(n_827), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_821), .B(n_846), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_821), .B(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AOI211xp5_ASAP7_75t_L g929 ( .A1(n_822), .A2(n_825), .B(n_871), .C(n_930), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_822), .B(n_832), .Y(n_968) );
OAI211xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B(n_829), .C(n_834), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_824), .B(n_832), .Y(n_855) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g898 ( .A(n_827), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_827), .B(n_885), .Y(n_930) );
A2O1A1Ixp33_ASAP7_75t_L g951 ( .A1(n_827), .A2(n_914), .B(n_941), .C(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g837 ( .A(n_828), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g918 ( .A(n_830), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g917 ( .A(n_833), .Y(n_917) );
OAI221xp5_ASAP7_75t_L g962 ( .A1(n_833), .A2(n_963), .B1(n_964), .B2(n_965), .C(n_967), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_837), .Y(n_834) );
A2O1A1Ixp33_ASAP7_75t_L g895 ( .A1(n_835), .A2(n_847), .B(n_896), .C(n_899), .Y(n_895) );
INVx2_ASAP7_75t_L g860 ( .A(n_836), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_836), .B(n_867), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_837), .B(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g950 ( .A(n_842), .Y(n_950) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_846), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_845), .B(n_881), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_847), .B(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g959 ( .A(n_847), .Y(n_959) );
AOI22xp5_ASAP7_75t_SL g943 ( .A1(n_848), .A2(n_870), .B1(n_944), .B2(n_962), .Y(n_943) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
O2A1O1Ixp33_ASAP7_75t_L g936 ( .A1(n_849), .A2(n_880), .B(n_937), .C(n_940), .Y(n_936) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_850), .B(n_867), .Y(n_866) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_850), .Y(n_871) );
OAI211xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B(n_859), .C(n_865), .Y(n_854) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
OR2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_863), .A2(n_897), .B(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g926 ( .A(n_864), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_872), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_SL g923 ( .A(n_872), .Y(n_923) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_878), .B(n_880), .C(n_882), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g912 ( .A1(n_878), .A2(n_913), .B1(n_915), .B2(n_918), .C(n_919), .Y(n_912) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
AOI211xp5_ASAP7_75t_SL g882 ( .A1(n_883), .A2(n_884), .B(n_887), .C(n_890), .Y(n_882) );
INVx1_ASAP7_75t_L g964 ( .A(n_883), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_884), .B(n_947), .Y(n_963) );
INVx1_ASAP7_75t_L g952 ( .A(n_888), .Y(n_952) );
INVx1_ASAP7_75t_L g942 ( .A(n_889), .Y(n_942) );
INVx1_ASAP7_75t_L g956 ( .A(n_891), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_892), .B(n_926), .Y(n_925) );
OAI21xp5_ASAP7_75t_SL g940 ( .A1(n_892), .A2(n_941), .B(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g947 ( .A(n_893), .Y(n_947) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_901), .C(n_902), .Y(n_894) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g932 ( .A(n_901), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_906), .B1(n_908), .B2(n_909), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_920), .B(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_931), .C(n_943), .Y(n_927) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NAND5xp2_ASAP7_75t_L g944 ( .A(n_945), .B(n_951), .C(n_953), .D(n_955), .E(n_957), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
INVxp67_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g969 ( .A(n_970), .Y(n_969) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g987 ( .A(n_973), .Y(n_987) );
NOR2xp67_ASAP7_75t_L g973 ( .A(n_974), .B(n_982), .Y(n_973) );
NAND4xp25_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .C(n_977), .D(n_980), .Y(n_974) );
NAND4xp25_ASAP7_75t_L g982 ( .A(n_983), .B(n_984), .C(n_985), .D(n_986), .Y(n_982) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVxp33_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
NAND2x1_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1008), .Y(n_1001) );
AND4x1_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1005), .C(n_1006), .D(n_1007), .Y(n_1002) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1020), .B1(n_1021), .B2(n_1022), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
endmodule