module fake_jpeg_25052_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_59),
.Y(n_86)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_24),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_35),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_40),
.B1(n_28),
.B2(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_43),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_21),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_16),
.B(n_20),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_21),
.B(n_25),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_40),
.B1(n_28),
.B2(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_42),
.B1(n_44),
.B2(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_71),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_75),
.B1(n_87),
.B2(n_105),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_83),
.B1(n_106),
.B2(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_77),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_69),
.B1(n_68),
.B2(n_58),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_44),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_89),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_52),
.C(n_64),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_90),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_85),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_43),
.C(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_54),
.B(n_24),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_27),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_96),
.A2(n_103),
.B(n_34),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_53),
.B(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_18),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_97),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_88),
.B1(n_108),
.B2(n_101),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_81),
.B(n_34),
.CI(n_22),
.CON(n_114),
.SN(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_34),
.B(n_96),
.C(n_33),
.D(n_19),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_22),
.B(n_25),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_34),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_53),
.B1(n_23),
.B2(n_39),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_105),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_23),
.B1(n_39),
.B2(n_38),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_30),
.B1(n_39),
.B2(n_38),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_132),
.B1(n_96),
.B2(n_99),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_43),
.B1(n_18),
.B2(n_33),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_0),
.B(n_1),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_73),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_100),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_141),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_75),
.C(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_135),
.C(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_136),
.B1(n_133),
.B2(n_114),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_155),
.B1(n_164),
.B2(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_163),
.B(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_76),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_73),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_84),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_123),
.B1(n_130),
.B2(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_159),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_85),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_88),
.B1(n_101),
.B2(n_80),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_80),
.B1(n_82),
.B2(n_78),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_78),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_113),
.B(n_109),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_125),
.A2(n_82),
.B1(n_43),
.B2(n_18),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_33),
.B1(n_19),
.B2(n_2),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_186),
.C(n_147),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_111),
.B1(n_120),
.B2(n_127),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_182),
.B1(n_189),
.B2(n_190),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_114),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_153),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_119),
.B1(n_109),
.B2(n_115),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_192),
.B(n_197),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_119),
.C(n_113),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_115),
.B1(n_127),
.B2(n_34),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_149),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_19),
.B1(n_8),
.B2(n_10),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_196),
.B1(n_163),
.B2(n_142),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_145),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_0),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_152),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_217),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_168),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_150),
.B1(n_156),
.B2(n_143),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_204),
.B(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_158),
.C(n_138),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_215),
.C(n_185),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_141),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_178),
.C(n_171),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_177),
.B(n_151),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_191),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_169),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_167),
.B1(n_7),
.B2(n_10),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_195),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_231),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_180),
.C(n_172),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_238),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_172),
.C(n_197),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_197),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_202),
.B1(n_179),
.B2(n_194),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_192),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_238),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_197),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_245),
.Y(n_254)
);

XOR2x2_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_197),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_257),
.B(n_198),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_202),
.B1(n_204),
.B2(n_201),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_248),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_252),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_217),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_240),
.A2(n_212),
.B1(n_219),
.B2(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_179),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_194),
.B1(n_218),
.B2(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_259),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_182),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_210),
.B1(n_184),
.B2(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_198),
.Y(n_262)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_228),
.C(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_265),
.C(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_235),
.C(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_225),
.C(n_233),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_229),
.C(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_200),
.B1(n_6),
.B2(n_11),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_274),
.A2(n_275),
.B1(n_271),
.B2(n_248),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_272),
.B1(n_261),
.B2(n_258),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_247),
.C(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_282),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_258),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_259),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_251),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_265),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_267),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_254),
.B(n_269),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

OAI21x1_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_278),
.B(n_285),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_295),
.B1(n_294),
.B2(n_15),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_280),
.C(n_6),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_15),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_301),
.B(n_2),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_298),
.A2(n_288),
.B(n_286),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_1),
.B(n_2),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_303),
.B(n_3),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_3),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_3),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_3),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_4),
.Y(n_308)
);


endmodule