module fake_jpeg_30271_n_330 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_330);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_19),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_1),
.Y(n_106)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_68),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_34),
.B1(n_38),
.B2(n_31),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_77),
.B1(n_83),
.B2(n_85),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_40),
.B1(n_23),
.B2(n_34),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_71),
.A2(n_86),
.B1(n_90),
.B2(n_15),
.Y(n_150)
);

AND2x4_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_22),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_107),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_34),
.B1(n_31),
.B2(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_40),
.B1(n_23),
.B2(n_42),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_94),
.B1(n_102),
.B2(n_7),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_31),
.B1(n_22),
.B2(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_22),
.B1(n_36),
.B2(n_25),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_39),
.B1(n_37),
.B2(n_42),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_108),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_110),
.B1(n_114),
.B2(n_8),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_29),
.B1(n_26),
.B2(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_26),
.B1(n_39),
.B2(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_1),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_65),
.A2(n_64),
.B1(n_66),
.B2(n_6),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_119),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_66),
.B(n_64),
.C(n_60),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_66),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_134),
.C(n_76),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_123),
.B(n_134),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_131),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_6),
.B(n_7),
.Y(n_126)
);

OR2x6_ASAP7_75t_L g185 ( 
.A(n_126),
.B(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_92),
.B(n_106),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_138),
.B1(n_90),
.B2(n_88),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_145),
.Y(n_158)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_7),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_8),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_91),
.B(n_112),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_8),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_143),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_9),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_9),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_80),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_87),
.B(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_87),
.B(n_17),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_76),
.A2(n_14),
.B1(n_15),
.B2(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_95),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_152),
.B1(n_113),
.B2(n_69),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_71),
.A2(n_15),
.B1(n_88),
.B2(n_73),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_153),
.A2(n_145),
.B1(n_135),
.B2(n_139),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_126),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_161),
.A2(n_162),
.B1(n_172),
.B2(n_187),
.Y(n_218)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_69),
.A3(n_109),
.B1(n_72),
.B2(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_174),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_95),
.B1(n_72),
.B2(n_104),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_136),
.B1(n_147),
.B2(n_120),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_111),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_177),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_122),
.B(n_80),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_118),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_121),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_125),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_125),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_136),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_130),
.B(n_142),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_190),
.B(n_199),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_150),
.B1(n_152),
.B2(n_149),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_191),
.A2(n_200),
.B1(n_203),
.B2(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_158),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_149),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_213),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_151),
.B1(n_115),
.B2(n_132),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_161),
.B1(n_185),
.B2(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_218),
.B1(n_173),
.B2(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_144),
.B1(n_141),
.B2(n_140),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_116),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_119),
.C(n_160),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_169),
.C(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_232),
.C(n_194),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_213),
.A2(n_185),
.B(n_162),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_238),
.B(n_243),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_185),
.B(n_163),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_243),
.B(n_221),
.C(n_224),
.Y(n_247)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_206),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_240),
.B1(n_198),
.B2(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_181),
.C(n_170),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_166),
.B1(n_173),
.B2(n_182),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_235),
.A2(n_228),
.B1(n_207),
.B2(n_224),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_156),
.B(n_171),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_192),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_171),
.B(n_182),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_200),
.B(n_209),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_190),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_248),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_197),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_253),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

OAI31xp33_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_262),
.A3(n_234),
.B(n_236),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_219),
.A2(n_196),
.B1(n_217),
.B2(n_211),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_258),
.B1(n_255),
.B2(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_214),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_264),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_231),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_235),
.C(n_220),
.Y(n_268)
);

AOI211xp5_ASAP7_75t_SL g266 ( 
.A1(n_247),
.A2(n_222),
.B(n_238),
.C(n_229),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_269),
.B1(n_248),
.B2(n_259),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_232),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_257),
.C(n_252),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_231),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_239),
.B1(n_234),
.B2(n_236),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_281),
.B1(n_250),
.B2(n_204),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_279),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_233),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_245),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_233),
.B1(n_225),
.B2(n_216),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_284),
.C(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_263),
.C(n_262),
.Y(n_284)
);

BUFx12f_ASAP7_75t_SL g285 ( 
.A(n_266),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_288),
.B(n_277),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_294),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_276),
.B1(n_273),
.B2(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_295),
.B1(n_275),
.B2(n_189),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_199),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_250),
.B1(n_225),
.B2(n_223),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_242),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_189),
.B1(n_188),
.B2(n_210),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_302),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_179),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_292),
.B(n_288),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_295),
.B(n_286),
.Y(n_307)
);

XOR2x2_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_283),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_294),
.C(n_293),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_284),
.A2(n_267),
.B(n_271),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_155),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_310),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_313),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_293),
.B(n_188),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_314),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_179),
.C(n_155),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_304),
.C(n_298),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_318),
.B(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_300),
.B1(n_297),
.B2(n_296),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_310),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_321),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_299),
.B(n_304),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_319),
.C(n_317),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_324),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_323),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_317),
.Y(n_330)
);


endmodule