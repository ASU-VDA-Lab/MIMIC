module fake_jpeg_91_n_531 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_24),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_53),
.B(n_77),
.Y(n_149)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx2_ASAP7_75t_SL g158 ( 
.A(n_59),
.Y(n_158)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_70),
.Y(n_124)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_19),
.B(n_12),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_32),
.B(n_12),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_89),
.Y(n_137)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_37),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_47),
.B1(n_41),
.B2(n_17),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_103),
.A2(n_110),
.B1(n_112),
.B2(n_115),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_41),
.B1(n_27),
.B2(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_47),
.B1(n_41),
.B2(n_17),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_59),
.A2(n_80),
.B1(n_47),
.B2(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_32),
.B1(n_45),
.B2(n_33),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_139),
.B1(n_148),
.B2(n_150),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_59),
.A2(n_17),
.B1(n_45),
.B2(n_43),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_153),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_21),
.B1(n_43),
.B2(n_38),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_69),
.A2(n_38),
.B1(n_33),
.B2(n_21),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_79),
.A2(n_29),
.B1(n_37),
.B2(n_34),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_71),
.A2(n_34),
.B1(n_42),
.B2(n_44),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_161),
.B1(n_0),
.B2(n_4),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_73),
.B(n_42),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_74),
.B(n_27),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_159),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_98),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_86),
.A2(n_50),
.B1(n_67),
.B2(n_81),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_99),
.B1(n_100),
.B2(n_72),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_168),
.A2(n_204),
.B1(n_209),
.B2(n_104),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_114),
.B(n_34),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_171),
.A2(n_205),
.B(n_210),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx2_ASAP7_75t_SL g213 ( 
.A(n_172),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_114),
.A2(n_96),
.B(n_40),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_178),
.B(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_176),
.B(n_179),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_88),
.B1(n_85),
.B2(n_58),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_177),
.A2(n_162),
.B1(n_118),
.B2(n_133),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_124),
.A2(n_19),
.B1(n_22),
.B2(n_55),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_22),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_185),
.Y(n_226)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_198),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_48),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_140),
.C(n_139),
.Y(n_212)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_90),
.B(n_81),
.C(n_78),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_115),
.B(n_161),
.C(n_112),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_78),
.B(n_68),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_132),
.A2(n_68),
.B1(n_11),
.B2(n_2),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_103),
.B1(n_150),
.B2(n_108),
.Y(n_232)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_200),
.Y(n_239)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_203),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_111),
.B(n_0),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_116),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_206),
.B(n_134),
.Y(n_243)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_116),
.B(n_0),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_120),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_243),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_163),
.B1(n_166),
.B2(n_207),
.Y(n_256)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_202),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_242),
.B1(n_190),
.B2(n_168),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_160),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_186),
.B(n_185),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_171),
.A2(n_151),
.B(n_141),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_247),
.B(n_173),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_196),
.B1(n_204),
.B2(n_169),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_189),
.A2(n_108),
.B1(n_136),
.B2(n_133),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_179),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_176),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_147),
.B(n_160),
.C(n_151),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_223),
.A2(n_178),
.B1(n_195),
.B2(n_208),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_254),
.B(n_219),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_188),
.B(n_194),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_208),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_255),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_165),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_201),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_242),
.B1(n_232),
.B2(n_243),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_270),
.B1(n_275),
.B2(n_246),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_200),
.B1(n_162),
.B2(n_106),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_211),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_277),
.Y(n_299)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_174),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_219),
.A2(n_233),
.B1(n_235),
.B2(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_211),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_211),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_217),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_248),
.A2(n_219),
.B1(n_233),
.B2(n_221),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_281),
.A2(n_295),
.B1(n_300),
.B2(n_301),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_219),
.B1(n_228),
.B2(n_240),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_285),
.B(n_254),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_266),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_252),
.A2(n_221),
.B1(n_240),
.B2(n_226),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_293),
.A2(n_305),
.B1(n_277),
.B2(n_271),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_303),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_251),
.A2(n_247),
.B1(n_226),
.B2(n_230),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_269),
.A2(n_247),
.B1(n_217),
.B2(n_246),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_231),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_231),
.B1(n_220),
.B2(n_239),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_222),
.B1(n_220),
.B2(n_227),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_309),
.B1(n_270),
.B2(n_258),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_256),
.A2(n_239),
.B1(n_106),
.B2(n_175),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_278),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_170),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_244),
.C(n_225),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_270),
.B1(n_250),
.B2(n_267),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_280),
.Y(n_318)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_321),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_314),
.A2(n_323),
.B1(n_337),
.B2(n_302),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_260),
.B1(n_259),
.B2(n_249),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_315),
.A2(n_327),
.B1(n_332),
.B2(n_218),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_318),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_273),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_319),
.B(n_326),
.Y(n_366)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

AO22x1_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_276),
.B1(n_253),
.B2(n_260),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_261),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_301),
.A2(n_254),
.B1(n_253),
.B2(n_264),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g375 ( 
.A1(n_329),
.A2(n_331),
.B(n_334),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_299),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_336),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_309),
.A2(n_255),
.B1(n_259),
.B2(n_268),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_255),
.B1(n_272),
.B2(n_263),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_255),
.B(n_237),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_333),
.A2(n_341),
.B(n_306),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_183),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_282),
.A2(n_289),
.B1(n_293),
.B2(n_305),
.Y(n_337)
);

XOR2x1_ASAP7_75t_L g338 ( 
.A(n_283),
.B(n_203),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_281),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_141),
.C(n_107),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_181),
.C(n_145),
.Y(n_349)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_342),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_283),
.A2(n_288),
.B(n_298),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_307),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_288),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_346),
.B(n_322),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_357),
.C(n_359),
.Y(n_398)
);

XOR2x2_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_337),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_326),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_351),
.B(n_367),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_318),
.B(n_292),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_354),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_292),
.B1(n_298),
.B2(n_302),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_323),
.B1(n_313),
.B2(n_328),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_360),
.B1(n_331),
.B2(n_327),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_356),
.A2(n_358),
.B(n_365),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_333),
.Y(n_357)
);

AO21x2_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_297),
.B(n_290),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_308),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_297),
.B1(n_290),
.B2(n_291),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_362),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_319),
.B(n_215),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_311),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_263),
.Y(n_369)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_107),
.C(n_244),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_372),
.C(n_373),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_311),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_336),
.C(n_340),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_225),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_198),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_182),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_339),
.C(n_215),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_378),
.Y(n_411)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_316),
.Y(n_384)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_386),
.B1(n_396),
.B2(n_402),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_407),
.B1(n_360),
.B2(n_374),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_391),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_357),
.Y(n_409)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_369),
.Y(n_390)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_316),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_393),
.Y(n_430)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_406),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_332),
.B1(n_334),
.B2(n_329),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_238),
.Y(n_431)
);

AOI21xp33_ASAP7_75t_L g399 ( 
.A1(n_345),
.A2(n_338),
.B(n_320),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_399),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_358),
.A2(n_325),
.B1(n_324),
.B2(n_312),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_375),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_215),
.C(n_145),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_363),
.C(n_349),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_238),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_345),
.A2(n_291),
.B1(n_272),
.B2(n_227),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_416),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_385),
.A2(n_358),
.B1(n_375),
.B2(n_356),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_379),
.B1(n_390),
.B2(n_407),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_412),
.B(n_420),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_359),
.C(n_372),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_414),
.B(n_417),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_350),
.C(n_376),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_383),
.A2(n_358),
.B(n_373),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_418),
.A2(n_167),
.B(n_218),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_419),
.A2(n_396),
.B1(n_393),
.B2(n_392),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_377),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_348),
.C(n_344),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_423),
.B(n_427),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_344),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_403),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_187),
.C(n_184),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_383),
.A2(n_238),
.B(n_192),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_428),
.Y(n_438)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_401),
.Y(n_434)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_414),
.C(n_417),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_436),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_389),
.C(n_404),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_382),
.Y(n_439)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_439),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_441),
.A2(n_413),
.B1(n_213),
.B2(n_180),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_402),
.B1(n_384),
.B2(n_379),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_447),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_444),
.A2(n_446),
.B1(n_452),
.B2(n_432),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_422),
.A2(n_391),
.B1(n_403),
.B2(n_397),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_431),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_450),
.Y(n_458)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_451),
.B(n_455),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_410),
.A2(n_213),
.B1(n_218),
.B2(n_183),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_419),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_421),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_453),
.C(n_436),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_459),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_434),
.Y(n_459)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_430),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_466),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_462),
.B(n_463),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_445),
.A2(n_418),
.B(n_428),
.Y(n_463)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_409),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_472),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_416),
.C(n_423),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_469),
.B(n_471),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_449),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_119),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_408),
.C(n_427),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_446),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_442),
.B(n_424),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_454),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_464),
.A2(n_444),
.B(n_460),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_484),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_438),
.C(n_437),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_482),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_461),
.A2(n_451),
.B1(n_447),
.B2(n_437),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_452),
.B1(n_147),
.B2(n_119),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_492),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_472),
.A2(n_128),
.B(n_199),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_487),
.A2(n_475),
.B(n_471),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_491),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_458),
.Y(n_490)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_490),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_119),
.C(n_191),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_481),
.B(n_468),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_496),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_469),
.Y(n_496)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_483),
.B(n_462),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_501),
.Y(n_508)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_479),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_486),
.A2(n_474),
.B(n_467),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_502),
.B(n_484),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_480),
.B(n_6),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_505),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_478),
.B(n_6),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_486),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_506),
.A2(n_487),
.B(n_8),
.C(n_9),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_477),
.C(n_476),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_508),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_509),
.A2(n_511),
.B(n_512),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_476),
.B(n_489),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_SL g512 ( 
.A(n_502),
.B(n_491),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_514),
.A2(n_493),
.B(n_500),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_493),
.A2(n_10),
.B(n_7),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_497),
.B(n_8),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_517),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_500),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_518),
.A2(n_522),
.B(n_516),
.Y(n_523)
);

OAI21xp33_ASAP7_75t_SL g525 ( 
.A1(n_519),
.A2(n_521),
.B(n_515),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_504),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_7),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_525),
.A2(n_526),
.B(n_7),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_7),
.B(n_10),
.Y(n_526)
);

AO21x1_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_528),
.B(n_524),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_7),
.C(n_10),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_10),
.B(n_509),
.Y(n_531)
);


endmodule