module fake_jpeg_3471_n_473 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_46),
.B(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_16),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_56),
.Y(n_116)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_71),
.Y(n_92)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_75),
.Y(n_110)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_0),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_24),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_19),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_38),
.B1(n_26),
.B2(n_27),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_90),
.A2(n_137),
.B1(n_79),
.B2(n_47),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_95),
.B(n_4),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_19),
.B1(n_42),
.B2(n_31),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_97),
.A2(n_99),
.B1(n_121),
.B2(n_135),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_19),
.B1(n_42),
.B2(n_31),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_45),
.B(n_43),
.C(n_27),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_59),
.B(n_61),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_50),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_111),
.B(n_112),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_45),
.B(n_43),
.Y(n_112)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_51),
.A2(n_19),
.B1(n_42),
.B2(n_31),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_44),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_44),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_78),
.A2(n_42),
.B1(n_31),
.B2(n_29),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_70),
.A2(n_38),
.B1(n_44),
.B2(n_22),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_44),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_142),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_84),
.A2(n_42),
.B1(n_31),
.B2(n_54),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_73),
.B1(n_82),
.B2(n_36),
.Y(n_180)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_63),
.B(n_44),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g187 ( 
.A(n_144),
.Y(n_187)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_53),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_148),
.B(n_167),
.Y(n_214)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_152),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_72),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_156),
.A2(n_191),
.B1(n_121),
.B2(n_135),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_157),
.B(n_172),
.Y(n_251)
);

CKINVDCx9p33_ASAP7_75t_R g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_159),
.Y(n_242)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_125),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_169),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_90),
.A2(n_24),
.B1(n_28),
.B2(n_30),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_163),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_252)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_125),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_22),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_91),
.B(n_55),
.C(n_80),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_183),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_128),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_36),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_177),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_52),
.B1(n_38),
.B2(n_77),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_175),
.A2(n_94),
.B1(n_132),
.B2(n_147),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_114),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_249)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_109),
.B(n_1),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_124),
.A2(n_32),
.B1(n_30),
.B2(n_28),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_114),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_192),
.Y(n_233)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_118),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_2),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_2),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_196),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_2),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_97),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_4),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_5),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_203),
.Y(n_244)
);

OAI22x1_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_100),
.B1(n_125),
.B2(n_99),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_204),
.A2(n_8),
.B(n_10),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_153),
.A3(n_171),
.B1(n_149),
.B2(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_205),
.B(n_221),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_226),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_216),
.B(n_150),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_148),
.B(n_153),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_220),
.A2(n_240),
.B(n_216),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_105),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_228),
.B1(n_161),
.B2(n_167),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_156),
.A2(n_96),
.B1(n_126),
.B2(n_106),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_249),
.B1(n_190),
.B2(n_182),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_165),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_175),
.A2(n_145),
.B1(n_108),
.B2(n_134),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_241),
.B1(n_166),
.B2(n_199),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_151),
.A2(n_94),
.B(n_134),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_232),
.A2(n_152),
.B(n_187),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_170),
.A2(n_98),
.B(n_145),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_98),
.B1(n_138),
.B2(n_146),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_138),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_189),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_248),
.B(n_217),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_166),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_206),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_253),
.Y(n_319)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_255),
.B(n_289),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_262),
.Y(n_302)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_258),
.B(n_261),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_214),
.A2(n_194),
.B(n_179),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_259),
.A2(n_294),
.B(n_229),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_229),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_209),
.B(n_150),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_270),
.B1(n_283),
.B2(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_206),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_220),
.A2(n_242),
.B1(n_228),
.B2(n_245),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_282),
.B1(n_241),
.B2(n_250),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_155),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_273),
.B(n_274),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_212),
.B(n_168),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_209),
.B(n_197),
.C(n_188),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_280),
.C(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_158),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_207),
.B(n_173),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_158),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_286),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_224),
.A2(n_181),
.B(n_164),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_279),
.A2(n_280),
.B(n_281),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_214),
.A2(n_160),
.B1(n_176),
.B2(n_203),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_204),
.A2(n_187),
.B1(n_182),
.B2(n_9),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_205),
.B(n_187),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_6),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_288),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_215),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_290),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g293 ( 
.A(n_224),
.B(n_11),
.C(n_12),
.Y(n_293)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_215),
.B(n_13),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_11),
.B(n_12),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_296),
.B(n_246),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_232),
.A2(n_13),
.B(n_249),
.C(n_230),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_208),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_208),
.B1(n_218),
.B2(n_231),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_298),
.A2(n_305),
.B1(n_307),
.B2(n_321),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_265),
.A2(n_244),
.B1(n_249),
.B2(n_247),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_300),
.A2(n_314),
.B1(n_315),
.B2(n_325),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_244),
.B1(n_249),
.B2(n_247),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_313),
.C(n_324),
.Y(n_353)
);

AO22x1_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_211),
.B1(n_237),
.B2(n_219),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_331),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_275),
.C(n_265),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_264),
.A2(n_222),
.B1(n_237),
.B2(n_211),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_278),
.A2(n_246),
.B1(n_231),
.B2(n_219),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_320),
.A2(n_295),
.B(n_284),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_266),
.A2(n_276),
.B1(n_253),
.B2(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_258),
.B(n_218),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_256),
.A2(n_222),
.B1(n_227),
.B2(n_217),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_259),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_262),
.A2(n_13),
.B1(n_227),
.B2(n_273),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_329),
.A2(n_294),
.B1(n_290),
.B2(n_285),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_288),
.A2(n_13),
.B1(n_227),
.B2(n_282),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_334),
.A2(n_283),
.B1(n_263),
.B2(n_274),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_339),
.B1(n_350),
.B2(n_335),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_259),
.B(n_281),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_344),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_331),
.A2(n_296),
.B1(n_277),
.B2(n_269),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_289),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_340),
.B(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_301),
.B(n_287),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_348),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_326),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_345),
.B(n_362),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_347),
.B(n_332),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_268),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_SL g349 ( 
.A(n_306),
.B(n_296),
.C(n_288),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_359),
.C(n_303),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_321),
.A2(n_263),
.B1(n_279),
.B2(n_254),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_304),
.B(n_267),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_357),
.Y(n_373)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_257),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_364),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_367),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_324),
.C(n_311),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_300),
.A2(n_312),
.B1(n_319),
.B2(n_305),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_360),
.A2(n_366),
.B1(n_334),
.B2(n_309),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_295),
.B(n_292),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_363),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_271),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_297),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_312),
.A2(n_308),
.B1(n_314),
.B2(n_298),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_307),
.A2(n_320),
.B(n_333),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_330),
.B(n_303),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_363),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_323),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_377),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_356),
.A2(n_335),
.B1(n_323),
.B2(n_336),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_371),
.A2(n_372),
.B1(n_351),
.B2(n_361),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_374),
.A2(n_378),
.B1(n_350),
.B2(n_346),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_360),
.A2(n_366),
.B1(n_343),
.B2(n_351),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_309),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_381),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_352),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_364),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_318),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_318),
.C(n_328),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_393),
.C(n_338),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_332),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_337),
.Y(n_395)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_339),
.Y(n_397)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_397),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_336),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_411),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_405),
.C(n_410),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_401),
.A2(n_374),
.B1(n_390),
.B2(n_393),
.Y(n_420)
);

AOI21x1_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_367),
.B(n_358),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_402),
.A2(n_407),
.B(n_401),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_403),
.A2(n_382),
.B1(n_387),
.B2(n_378),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_349),
.C(n_365),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_415),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_346),
.Y(n_408)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_408),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_344),
.C(n_383),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_385),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_386),
.Y(n_412)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_392),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_372),
.A2(n_373),
.B1(n_371),
.B2(n_384),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_376),
.B1(n_381),
.B2(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_373),
.Y(n_416)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_417),
.A2(n_429),
.B1(n_418),
.B2(n_419),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_408),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_431),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_420),
.A2(n_424),
.B1(n_406),
.B2(n_413),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_376),
.Y(n_426)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_428),
.A2(n_433),
.B(n_398),
.Y(n_440)
);

INVx13_ASAP7_75t_L g431 ( 
.A(n_412),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_433),
.A2(n_402),
.B(n_403),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_435),
.A2(n_439),
.B(n_432),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_409),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_438),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_410),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_420),
.A2(n_405),
.B(n_400),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_447),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_398),
.C(n_406),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_445),
.C(n_421),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_427),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_444),
.A2(n_425),
.B1(n_434),
.B2(n_430),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_424),
.C(n_426),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_418),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_444),
.A2(n_429),
.B1(n_434),
.B2(n_425),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_449),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_450),
.B(n_453),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_437),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_454),
.A2(n_435),
.B(n_447),
.Y(n_461)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_446),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_455),
.B(n_456),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g458 ( 
.A1(n_451),
.A2(n_439),
.B(n_442),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_460),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_454),
.A2(n_440),
.B(n_446),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_452),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_456),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_465),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_452),
.Y(n_465)
);

OAI21xp33_ASAP7_75t_L g468 ( 
.A1(n_466),
.A2(n_457),
.B(n_450),
.Y(n_468)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g469 ( 
.A1(n_468),
.A2(n_464),
.B(n_466),
.C(n_453),
.D(n_449),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_469),
.B(n_467),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_441),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_471),
.A2(n_445),
.B(n_443),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_472),
.B(n_443),
.Y(n_473)
);


endmodule