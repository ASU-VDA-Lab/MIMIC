module real_jpeg_12920_n_17 (n_5, n_4, n_8, n_0, n_12, n_251, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_251;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_5),
.A2(n_31),
.B1(n_37),
.B2(n_39),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_7),
.A2(n_37),
.B1(n_39),
.B2(n_59),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_59),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_59),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_37),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_8),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_46),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_10),
.B(n_55),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_10),
.A2(n_37),
.B1(n_39),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_26),
.C(n_42),
.Y(n_145)
);

NAND2x1_ASAP7_75t_SL g149 ( 
.A(n_10),
.B(n_64),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_100),
.B(n_156),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_51),
.B(n_65),
.C(n_183),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_10),
.B(n_205),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_12),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_12),
.B(n_52),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_61),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_61),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_37),
.B1(n_39),
.B2(n_70),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_15),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_84)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_20),
.B(n_105),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.C(n_62),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_22),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_23),
.B(n_34),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_24),
.A2(n_29),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_24),
.A2(n_29),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_24),
.B(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_25),
.B(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_29),
.B(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_32),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_37),
.B(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_39),
.A2(n_66),
.B(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_40),
.A2(n_47),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_40),
.A2(n_45),
.B1(n_47),
.B2(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_40),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_40),
.B(n_143),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_40),
.A2(n_47),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_44),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_44),
.B(n_141),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_44),
.A2(n_153),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_47),
.B(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_62),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_60),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_49),
.A2(n_56),
.B(n_141),
.C(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_50),
.A2(n_58),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_50),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_51),
.A2(n_53),
.A3(n_56),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B(n_68),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_67),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_63),
.A2(n_68),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_63),
.A2(n_91),
.B1(n_118),
.B2(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2x1_ASAP7_75t_R g71 ( 
.A(n_64),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_69),
.Y(n_119)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_86),
.B2(n_87),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_85),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_97),
.B2(n_104),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_91),
.A2(n_119),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_95),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_101),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_100),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_100),
.A2(n_101),
.B1(n_126),
.B2(n_185),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_101),
.A2(n_162),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_141),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_101),
.A2(n_170),
.B(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_110),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_106),
.B(n_108),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_110),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_120),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_238)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_120),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_234),
.A3(n_243),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_216),
.B(n_233),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_195),
.B(n_215),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_178),
.B(n_194),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_158),
.B(n_177),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_146),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_142),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_139),
.A2(n_142),
.B(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_151),
.C(n_154),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_166),
.B(n_176),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B(n_175),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_180),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_189),
.C(n_193),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_184),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_208),
.B2(n_209),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_211),
.C(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_203),
.C(n_207),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_229),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_230),
.C(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_228),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_225),
.C(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_241),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_237),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule