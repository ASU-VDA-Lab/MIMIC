module fake_jpeg_851_n_117 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_3),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_50),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_37),
.B1(n_42),
.B2(n_38),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_53),
.B(n_50),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_46),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_35),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_34),
.B1(n_38),
.B2(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_50),
.B1(n_49),
.B2(n_37),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_43),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_72),
.C(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_71),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_69),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_33),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_25),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_71),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.C(n_95),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_1),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_85),
.B(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_1),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_18),
.C(n_17),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_4),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_103),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_90),
.B1(n_87),
.B2(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_105),
.B1(n_89),
.B2(n_8),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_79),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_101),
.B1(n_102),
.B2(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_104),
.C(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_111),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_106),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_6),
.C2(n_11),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_9),
.B(n_10),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_12),
.Y(n_117)
);


endmodule