module fake_jpeg_16297_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_43),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_68),
.B(n_23),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_84),
.B1(n_91),
.B2(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_19),
.B1(n_26),
.B2(n_28),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_70),
.A2(n_72),
.B1(n_77),
.B2(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_26),
.B1(n_29),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_26),
.B1(n_21),
.B2(n_16),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_2),
.B(n_3),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_79),
.A2(n_98),
.B(n_86),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_38),
.A2(n_34),
.B1(n_22),
.B2(n_33),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_29),
.B1(n_32),
.B2(n_37),
.Y(n_84)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_113),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_41),
.A2(n_29),
.B1(n_14),
.B2(n_32),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_37),
.B1(n_32),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_16),
.B1(n_14),
.B2(n_21),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_95),
.B1(n_102),
.B2(n_103),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_34),
.B1(n_22),
.B2(n_33),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_28),
.B1(n_25),
.B2(n_15),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_30),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_42),
.B(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_25),
.B1(n_15),
.B2(n_23),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_109),
.B1(n_34),
.B2(n_22),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_30),
.B1(n_23),
.B2(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_40),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_36),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_36),
.B1(n_31),
.B2(n_30),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_62),
.B1(n_57),
.B2(n_48),
.Y(n_131)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_64),
.B1(n_58),
.B2(n_57),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_120),
.A2(n_116),
.B1(n_99),
.B2(n_112),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_123),
.B(n_132),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_126),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_36),
.Y(n_127)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_129),
.Y(n_201)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_116),
.B1(n_111),
.B2(n_97),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_47),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_96),
.C(n_31),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_2),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_141),
.B1(n_113),
.B2(n_87),
.Y(n_191)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_73),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_72),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_3),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_137),
.B1(n_124),
.B2(n_132),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_4),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_168),
.Y(n_198)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_77),
.B(n_36),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_78),
.B(n_44),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_85),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_89),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_75),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_89),
.B(n_36),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_4),
.Y(n_168)
);

OR2x2_ASAP7_75t_SL g169 ( 
.A(n_104),
.B(n_5),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_99),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_171),
.A2(n_137),
.B(n_124),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_120),
.B1(n_165),
.B2(n_144),
.Y(n_218)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_191),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_112),
.B1(n_111),
.B2(n_110),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_192),
.B1(n_197),
.B2(n_207),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_202),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_208),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_188),
.A2(n_169),
.B1(n_121),
.B2(n_147),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_122),
.Y(n_238)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_128),
.A2(n_118),
.B1(n_114),
.B2(n_97),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_133),
.B(n_96),
.C(n_92),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_119),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_142),
.A2(n_36),
.B1(n_31),
.B2(n_8),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_5),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_148),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_141),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_124),
.B(n_5),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_214),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_120),
.A2(n_31),
.B1(n_8),
.B2(n_9),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_178),
.B1(n_202),
.B2(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_120),
.A2(n_31),
.B1(n_8),
.B2(n_9),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_186),
.B(n_145),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_217),
.B(n_257),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_218),
.A2(n_223),
.B1(n_224),
.B2(n_230),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_222),
.B(n_242),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_119),
.B1(n_168),
.B2(n_152),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_205),
.B1(n_212),
.B2(n_193),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_176),
.Y(n_261)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_234),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_132),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_241),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_141),
.B1(n_147),
.B2(n_160),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_237),
.B1(n_240),
.B2(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_143),
.B1(n_139),
.B2(n_155),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_245),
.C(n_223),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_177),
.A2(n_122),
.B(n_143),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_242),
.B(n_245),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_163),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_180),
.A2(n_151),
.B(n_146),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_187),
.A2(n_135),
.B1(n_9),
.B2(n_10),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_171),
.B(n_31),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_187),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_249),
.B1(n_181),
.B2(n_175),
.Y(n_269)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_149),
.B1(n_11),
.B2(n_13),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_10),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_254),
.B(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_211),
.B(n_10),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_11),
.B(n_13),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_208),
.B(n_13),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_194),
.B1(n_172),
.B2(n_209),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_291),
.B(n_234),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_268),
.C(n_279),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_264),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_253),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_203),
.C(n_182),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_269),
.B(n_288),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_226),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_274),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_175),
.B1(n_181),
.B2(n_214),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_277),
.B1(n_252),
.B2(n_255),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_174),
.B1(n_179),
.B2(n_189),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_190),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_190),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_282),
.C(n_284),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_204),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_227),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_189),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_226),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_227),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_251),
.A2(n_170),
.B1(n_174),
.B2(n_196),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_251),
.B(n_239),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_299),
.B(n_316),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_298),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_307),
.B1(n_318),
.B2(n_269),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_259),
.A2(n_218),
.B(n_233),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_305),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_258),
.A2(n_231),
.B1(n_237),
.B2(n_219),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_306),
.B1(n_291),
.B2(n_290),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_243),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_278),
.A2(n_231),
.B1(n_254),
.B2(n_248),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_247),
.B1(n_249),
.B2(n_246),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_314),
.C(n_304),
.Y(n_341)
);

BUFx2_ASAP7_75t_SL g312 ( 
.A(n_263),
.Y(n_312)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_254),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_317),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_275),
.A2(n_220),
.B(n_252),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_283),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_267),
.A2(n_170),
.B1(n_220),
.B2(n_256),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_275),
.B(n_195),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_276),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_322),
.B(n_311),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_282),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_325),
.C(n_326),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_261),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_279),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_280),
.C(n_271),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_328),
.C(n_337),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_271),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_331),
.A2(n_319),
.B1(n_318),
.B2(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_277),
.B(n_273),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_297),
.B(n_299),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_284),
.C(n_260),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_268),
.C(n_236),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_341),
.C(n_337),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_302),
.A2(n_236),
.B1(n_272),
.B2(n_303),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_339),
.A2(n_302),
.B1(n_296),
.B2(n_305),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_294),
.Y(n_340)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_340),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_324),
.B(n_321),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_345),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_331),
.A2(n_336),
.B1(n_334),
.B2(n_333),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_346),
.A2(n_353),
.B1(n_343),
.B2(n_352),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_317),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_347),
.B(n_355),
.C(n_359),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_292),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_351),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_352),
.B1(n_354),
.B2(n_356),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_336),
.A2(n_310),
.B1(n_295),
.B2(n_313),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_333),
.A2(n_295),
.B1(n_315),
.B2(n_293),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_293),
.B1(n_311),
.B2(n_308),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_330),
.A2(n_342),
.B1(n_341),
.B2(n_322),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_342),
.B1(n_329),
.B2(n_339),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_357),
.B(n_327),
.Y(n_365)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_326),
.C(n_325),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_350),
.A2(n_324),
.B(n_328),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_367),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_359),
.Y(n_363)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_363),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_364),
.A2(n_365),
.B(n_356),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_350),
.A2(n_321),
.B(n_323),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_371),
.C(n_373),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_372),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_346),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_377),
.A2(n_367),
.B(n_362),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_360),
.C(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_368),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_382),
.B(n_376),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_374),
.A2(n_364),
.B(n_366),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_383),
.B(n_384),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_387),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_382),
.Y(n_387)
);

OAI31xp33_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_378),
.A3(n_363),
.B(n_361),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_388),
.Y(n_390)
);

OAI211xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_389),
.B(n_372),
.C(n_376),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_361),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_370),
.C(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_393),
.B(n_345),
.Y(n_394)
);

OAI321xp33_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_378),
.A3(n_375),
.B1(n_355),
.B2(n_348),
.C(n_358),
.Y(n_395)
);


endmodule