module real_aes_7226_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_725;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g473 ( .A1(n_0), .A2(n_163), .B(n_474), .C(n_477), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_1), .B(n_468), .Y(n_478) );
INVx1_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
INVx1_ASAP7_75t_L g161 ( .A(n_3), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_4), .B(n_164), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_5), .A2(n_463), .B(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_6), .A2(n_78), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_6), .Y(n_122) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_6), .A2(n_186), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_7), .A2(n_40), .B1(n_151), .B2(n_209), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_8), .A2(n_9), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_8), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_9), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_10), .B(n_186), .Y(n_194) );
AND2x6_ASAP7_75t_L g166 ( .A(n_11), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_12), .A2(n_166), .B(n_454), .C(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_13), .B(n_41), .Y(n_119) );
INVx1_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
INVx1_ASAP7_75t_L g142 ( .A(n_15), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_16), .B(n_147), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_17), .B(n_164), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_18), .B(n_138), .Y(n_196) );
AO32x2_ASAP7_75t_L g247 ( .A1(n_19), .A2(n_137), .A3(n_180), .B1(n_186), .B2(n_248), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_20), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_20), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_21), .A2(n_32), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_21), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_22), .B(n_151), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_23), .B(n_138), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_24), .A2(n_57), .B1(n_151), .B2(n_209), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g211 ( .A1(n_25), .A2(n_83), .B1(n_147), .B2(n_151), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_26), .B(n_151), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_27), .A2(n_180), .B(n_454), .C(n_485), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_28), .A2(n_180), .B(n_454), .C(n_547), .Y(n_546) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_29), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_30), .A2(n_729), .B1(n_730), .B2(n_733), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_30), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_31), .B(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_32), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_32), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_33), .A2(n_463), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_34), .B(n_182), .Y(n_224) );
INVx2_ASAP7_75t_L g149 ( .A(n_35), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_36), .A2(n_460), .B(n_503), .C(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_37), .B(n_151), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_38), .B(n_182), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_39), .B(n_231), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_42), .B(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_43), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_44), .B(n_164), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_45), .B(n_463), .Y(n_545) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_46), .A2(n_438), .B1(n_724), .B2(n_725), .C1(n_734), .C2(n_737), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_47), .A2(n_460), .B(n_503), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_48), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_49), .B(n_151), .Y(n_189) );
INVx1_ASAP7_75t_L g475 ( .A(n_50), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_51), .A2(n_92), .B1(n_209), .B2(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g528 ( .A(n_52), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_53), .B(n_151), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_54), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_55), .B(n_463), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_56), .B(n_159), .Y(n_193) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_58), .A2(n_62), .B1(n_147), .B2(n_151), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_59), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_60), .B(n_151), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_61), .B(n_151), .Y(n_228) );
INVx1_ASAP7_75t_L g167 ( .A(n_63), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_64), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_65), .B(n_468), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_66), .A2(n_153), .B(n_159), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_67), .B(n_151), .Y(n_162) );
INVx1_ASAP7_75t_L g141 ( .A(n_68), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_69), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_70), .B(n_164), .Y(n_506) );
AO32x2_ASAP7_75t_L g206 ( .A1(n_71), .A2(n_180), .A3(n_186), .B1(n_207), .B2(n_212), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_72), .B(n_165), .Y(n_519) );
INVx1_ASAP7_75t_L g176 ( .A(n_73), .Y(n_176) );
INVx1_ASAP7_75t_L g219 ( .A(n_74), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_75), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_76), .B(n_487), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_77), .A2(n_454), .B(n_456), .C(n_460), .Y(n_453) );
INVx1_ASAP7_75t_L g123 ( .A(n_78), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_79), .B(n_147), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_80), .Y(n_537) );
INVx1_ASAP7_75t_L g746 ( .A(n_81), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_82), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_84), .B(n_209), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_85), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_86), .B(n_147), .Y(n_223) );
INVx2_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_88), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_89), .B(n_179), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_90), .B(n_147), .Y(n_190) );
OR2x2_ASAP7_75t_L g115 ( .A(n_91), .B(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g441 ( .A(n_91), .B(n_117), .Y(n_441) );
INVx2_ASAP7_75t_L g445 ( .A(n_91), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_93), .A2(n_104), .B1(n_147), .B2(n_148), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_94), .B(n_463), .Y(n_501) );
INVx1_ASAP7_75t_L g505 ( .A(n_95), .Y(n_505) );
AOI22xp5_ASAP7_75t_SL g105 ( .A1(n_96), .A2(n_106), .B1(n_742), .B2(n_748), .Y(n_105) );
INVxp67_ASAP7_75t_L g540 ( .A(n_97), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_98), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_99), .B(n_147), .Y(n_174) );
INVx1_ASAP7_75t_L g457 ( .A(n_100), .Y(n_457) );
INVx1_ASAP7_75t_L g515 ( .A(n_101), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_102), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g530 ( .A(n_103), .B(n_182), .Y(n_530) );
OA21x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_111), .B(n_436), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g741 ( .A(n_109), .Y(n_741) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_120), .B(n_434), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g435 ( .A(n_115), .Y(n_435) );
INVx1_ASAP7_75t_SL g747 ( .A(n_115), .Y(n_747) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_116), .B(n_445), .Y(n_739) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g444 ( .A(n_117), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_130), .B2(n_433), .Y(n_125) );
INVx1_ASAP7_75t_L g433 ( .A(n_126), .Y(n_433) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR5x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_324), .C(n_382), .D(n_418), .E(n_425), .Y(n_130) );
NAND3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_270), .C(n_294), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_202), .B1(n_236), .B2(n_241), .C(n_251), .Y(n_132) );
OAI21xp5_ASAP7_75t_SL g404 ( .A1(n_133), .A2(n_405), .B(n_407), .Y(n_404) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_183), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_134), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
INVx2_ASAP7_75t_L g240 ( .A(n_135), .Y(n_240) );
AND2x2_ASAP7_75t_L g253 ( .A(n_135), .B(n_185), .Y(n_253) );
AND2x2_ASAP7_75t_L g307 ( .A(n_135), .B(n_184), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_135), .B(n_170), .Y(n_322) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_168), .Y(n_135) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_136), .A2(n_171), .B(n_181), .Y(n_170) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_137), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_139), .B(n_140), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_157), .B(n_166), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_150), .C(n_153), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_146), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_146), .A2(n_548), .B(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx3_ASAP7_75t_L g218 ( .A(n_151), .Y(n_218) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_151), .Y(n_459) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g209 ( .A(n_152), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_152), .Y(n_210) );
AND2x6_ASAP7_75t_L g454 ( .A(n_152), .B(n_455), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_153), .A2(n_457), .B(n_458), .C(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_154), .A2(n_222), .B(n_223), .Y(n_221) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g487 ( .A(n_155), .Y(n_487) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g165 ( .A(n_156), .Y(n_165) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
INVx1_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
INVx1_ASAP7_75t_L g455 ( .A(n_156), .Y(n_455) );
AND2x2_ASAP7_75t_L g464 ( .A(n_156), .B(n_160), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_162), .C(n_163), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_158), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_158), .A2(n_486), .B(n_488), .Y(n_485) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_163), .A2(n_192), .B(n_193), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_163), .A2(n_179), .B1(n_199), .B2(n_200), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_163), .A2(n_179), .B1(n_249), .B2(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_164), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_164), .A2(n_189), .B(n_190), .Y(n_188) );
O2A1O1Ixp5_ASAP7_75t_SL g217 ( .A1(n_164), .A2(n_218), .B(n_219), .C(n_220), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_164), .B(n_540), .Y(n_539) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g207 ( .A1(n_165), .A2(n_179), .B1(n_208), .B2(n_211), .Y(n_207) );
BUFx3_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_166), .A2(n_188), .B(n_191), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_166), .A2(n_217), .B(n_221), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_166), .A2(n_227), .B(n_232), .Y(n_226) );
INVx4_ASAP7_75t_SL g461 ( .A(n_166), .Y(n_461) );
AND2x4_ASAP7_75t_L g463 ( .A(n_166), .B(n_464), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_166), .B(n_464), .Y(n_516) );
AND2x2_ASAP7_75t_L g340 ( .A(n_169), .B(n_281), .Y(n_340) );
AND2x2_ASAP7_75t_L g373 ( .A(n_169), .B(n_185), .Y(n_373) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g280 ( .A(n_170), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g293 ( .A(n_170), .B(n_185), .Y(n_293) );
AND2x2_ASAP7_75t_L g300 ( .A(n_170), .B(n_281), .Y(n_300) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_170), .Y(n_309) );
AND2x2_ASAP7_75t_L g316 ( .A(n_170), .B(n_184), .Y(n_316) );
INVx1_ASAP7_75t_L g347 ( .A(n_170), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_180), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_178), .A2(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g476 ( .A(n_179), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g197 ( .A(n_180), .B(n_198), .C(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g212 ( .A(n_182), .Y(n_212) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_182), .A2(n_216), .B(n_224), .Y(n_215) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_182), .A2(n_226), .B(n_235), .Y(n_225) );
INVx1_ASAP7_75t_L g493 ( .A(n_182), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_182), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_182), .A2(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g323 ( .A(n_183), .Y(n_323) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_195), .Y(n_183) );
INVx2_ASAP7_75t_L g279 ( .A(n_184), .Y(n_279) );
AND2x2_ASAP7_75t_L g301 ( .A(n_184), .B(n_240), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_184), .B(n_347), .Y(n_352) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_185), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g424 ( .A(n_185), .B(n_388), .Y(n_424) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_194), .Y(n_185) );
INVx4_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_186), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_186), .A2(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
INVx3_ASAP7_75t_L g339 ( .A(n_195), .Y(n_339) );
OR2x2_ASAP7_75t_L g369 ( .A(n_195), .B(n_370), .Y(n_369) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_195), .B(n_279), .Y(n_395) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
AO21x1_ASAP7_75t_L g281 ( .A1(n_198), .A2(n_201), .B(n_282), .Y(n_281) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_201), .A2(n_452), .B(n_465), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_201), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g468 ( .A(n_201), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_201), .B(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_201), .A2(n_514), .B(n_521), .Y(n_513) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_202), .A2(n_253), .A3(n_267), .B1(n_339), .B2(n_416), .B3(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
OR2x2_ASAP7_75t_L g268 ( .A(n_204), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_204), .B(n_265), .Y(n_327) );
OR2x2_ASAP7_75t_L g380 ( .A(n_204), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g306 ( .A(n_205), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g331 ( .A(n_205), .B(n_213), .Y(n_331) );
AND2x2_ASAP7_75t_L g398 ( .A(n_205), .B(n_243), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_205), .A2(n_298), .B(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
INVx1_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
AND2x2_ASAP7_75t_L g277 ( .A(n_206), .B(n_247), .Y(n_277) );
AND2x2_ASAP7_75t_L g326 ( .A(n_206), .B(n_246), .Y(n_326) );
INVx2_ASAP7_75t_L g477 ( .A(n_210), .Y(n_477) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_210), .Y(n_507) );
INVx1_ASAP7_75t_L g490 ( .A(n_212), .Y(n_490) );
INVx2_ASAP7_75t_SL g368 ( .A(n_213), .Y(n_368) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
INVx2_ASAP7_75t_L g288 ( .A(n_214), .Y(n_288) );
INVx1_ASAP7_75t_L g419 ( .A(n_214), .Y(n_419) );
AND2x2_ASAP7_75t_L g432 ( .A(n_214), .B(n_313), .Y(n_432) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g259 ( .A(n_215), .Y(n_259) );
OR2x2_ASAP7_75t_L g265 ( .A(n_215), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_215), .Y(n_276) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_225), .Y(n_243) );
AND2x2_ASAP7_75t_L g260 ( .A(n_225), .B(n_246), .Y(n_260) );
INVx1_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
INVx1_ASAP7_75t_L g273 ( .A(n_225), .Y(n_273) );
AND2x2_ASAP7_75t_L g298 ( .A(n_225), .B(n_247), .Y(n_298) );
INVx2_ASAP7_75t_L g314 ( .A(n_225), .Y(n_314) );
AND2x2_ASAP7_75t_L g407 ( .A(n_225), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_225), .B(n_288), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g262 ( .A(n_238), .Y(n_262) );
INVx1_ASAP7_75t_L g291 ( .A(n_238), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_238), .B(n_322), .Y(n_388) );
INVx1_ASAP7_75t_SL g348 ( .A(n_239), .Y(n_348) );
INVx2_ASAP7_75t_L g269 ( .A(n_240), .Y(n_269) );
AND2x2_ASAP7_75t_L g338 ( .A(n_240), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g354 ( .A(n_240), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx1_ASAP7_75t_L g416 ( .A(n_242), .Y(n_416) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g271 ( .A(n_244), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g374 ( .A(n_244), .B(n_364), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_244), .A2(n_385), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g287 ( .A(n_245), .B(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g312 ( .A(n_245), .Y(n_312) );
INVx1_ASAP7_75t_L g336 ( .A(n_245), .Y(n_336) );
OR2x2_ASAP7_75t_L g400 ( .A(n_246), .B(n_259), .Y(n_400) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_246), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g313 ( .A(n_247), .B(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_254), .B1(n_261), .B2(n_263), .Y(n_251) );
OR2x2_ASAP7_75t_L g330 ( .A(n_252), .B(n_280), .Y(n_330) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_253), .A2(n_372), .B1(n_374), .B2(n_375), .C1(n_376), .C2(n_379), .Y(n_371) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_260), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g318 ( .A(n_257), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_259), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_259), .Y(n_343) );
AND2x2_ASAP7_75t_L g391 ( .A(n_259), .B(n_260), .Y(n_391) );
INVx1_ASAP7_75t_L g409 ( .A(n_259), .Y(n_409) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g375 ( .A(n_262), .B(n_301), .Y(n_375) );
AND2x2_ASAP7_75t_L g417 ( .A(n_262), .B(n_293), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_264), .B(n_312), .Y(n_399) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_265), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g292 ( .A(n_269), .B(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g360 ( .A(n_269), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B(n_278), .C(n_283), .Y(n_270) );
INVxp67_ASAP7_75t_L g284 ( .A(n_271), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_272), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_272), .B(n_319), .Y(n_414) );
BUFx3_ASAP7_75t_L g378 ( .A(n_273), .Y(n_378) );
INVx1_ASAP7_75t_L g285 ( .A(n_274), .Y(n_285) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g304 ( .A(n_276), .B(n_298), .Y(n_304) );
INVx1_ASAP7_75t_SL g344 ( .A(n_277), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g334 ( .A(n_279), .Y(n_334) );
AND2x2_ASAP7_75t_L g357 ( .A(n_279), .B(n_340), .Y(n_357) );
INVx1_ASAP7_75t_SL g328 ( .A(n_280), .Y(n_328) );
INVx1_ASAP7_75t_L g355 ( .A(n_281), .Y(n_355) );
AOI31xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .A3(n_286), .B(n_289), .Y(n_283) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g376 ( .A(n_287), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g350 ( .A(n_288), .Y(n_350) );
BUFx2_ASAP7_75t_L g364 ( .A(n_288), .Y(n_364) );
AND2x2_ASAP7_75t_L g392 ( .A(n_288), .B(n_313), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g365 ( .A(n_292), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_293), .B(n_360), .Y(n_406) );
AND2x2_ASAP7_75t_L g413 ( .A(n_293), .B(n_339), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_299), .B(n_302), .C(n_317), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_299), .A2(n_326), .B1(n_327), .B2(n_328), .C(n_329), .Y(n_325) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g333 ( .A(n_300), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g370 ( .A(n_301), .Y(n_370) );
OAI32xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .A3(n_308), .B1(n_310), .B2(n_315), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_304), .A2(n_357), .B(n_358), .C(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
OAI21xp5_ASAP7_75t_SL g420 ( .A1(n_312), .A2(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g381 ( .A(n_313), .Y(n_381) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_319), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NAND4xp25_ASAP7_75t_SL g324 ( .A(n_325), .B(n_337), .C(n_356), .D(n_371), .Y(n_324) );
AND2x2_ASAP7_75t_L g363 ( .A(n_326), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g385 ( .A(n_326), .B(n_378), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_328), .B(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_332), .B2(n_335), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_330), .A2(n_381), .B1(n_412), .B2(n_414), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_330), .A2(n_419), .B(n_420), .C(n_423), .Y(n_418) );
INVx2_ASAP7_75t_L g389 ( .A(n_331), .Y(n_389) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_333), .A2(n_367), .B1(n_384), .B2(n_385), .C1(n_386), .C2(n_389), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_341), .C(n_345), .Y(n_337) );
INVx1_ASAP7_75t_L g403 ( .A(n_338), .Y(n_403) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_342), .A2(n_346), .B1(n_349), .B2(n_351), .Y(n_345) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g372 ( .A(n_354), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g430 ( .A(n_357), .Y(n_430) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_366), .B2(n_369), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_364), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g421 ( .A(n_369), .Y(n_421) );
INVx1_ASAP7_75t_L g402 ( .A(n_373), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_375), .Y(n_429) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND5xp2_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .C(n_404), .D(n_410), .E(n_415), .Y(n_382) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_393), .C(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI31xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .A3(n_400), .B(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g422 ( .A(n_398), .Y(n_422) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI222xp33_ASAP7_75t_L g425 ( .A1(n_412), .A2(n_414), .B1(n_426), .B2(n_429), .C1(n_430), .C2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_434), .B(n_437), .C(n_740), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_443), .B2(n_446), .Y(n_439) );
INVx2_ASAP7_75t_L g735 ( .A(n_440), .Y(n_735) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_442), .A2(n_446), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g736 ( .A(n_443), .Y(n_736) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR3x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_632), .C(n_681), .Y(n_446) );
NAND5xp2_ASAP7_75t_L g447 ( .A(n_448), .B(n_566), .C(n_595), .D(n_603), .E(n_618), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_494), .B(n_510), .C(n_550), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_479), .Y(n_449) );
AND2x2_ASAP7_75t_L g561 ( .A(n_450), .B(n_558), .Y(n_561) );
AND2x2_ASAP7_75t_L g594 ( .A(n_450), .B(n_480), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_450), .B(n_498), .Y(n_687) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_467), .Y(n_450) );
INVx2_ASAP7_75t_L g497 ( .A(n_451), .Y(n_497) );
BUFx2_ASAP7_75t_L g661 ( .A(n_451), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
INVx5_ASAP7_75t_L g472 ( .A(n_454), .Y(n_472) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g470 ( .A1(n_461), .A2(n_471), .B(n_472), .C(n_473), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_461), .A2(n_472), .B(n_537), .C(n_538), .Y(n_536) );
BUFx2_ASAP7_75t_L g483 ( .A(n_463), .Y(n_483) );
AND2x2_ASAP7_75t_L g479 ( .A(n_467), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g559 ( .A(n_467), .Y(n_559) );
AND2x2_ASAP7_75t_L g645 ( .A(n_467), .B(n_558), .Y(n_645) );
AND2x2_ASAP7_75t_L g700 ( .A(n_467), .B(n_497), .Y(n_700) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_478), .Y(n_467) );
INVx2_ASAP7_75t_L g503 ( .A(n_472), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g617 ( .A(n_479), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_479), .B(n_498), .Y(n_664) );
INVx5_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
AND2x4_ASAP7_75t_L g579 ( .A(n_480), .B(n_559), .Y(n_579) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_480), .Y(n_601) );
AND2x2_ASAP7_75t_L g676 ( .A(n_480), .B(n_661), .Y(n_676) );
AND2x2_ASAP7_75t_L g679 ( .A(n_480), .B(n_499), .Y(n_679) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
AOI21xp5_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_484), .B(n_490), .Y(n_481) );
INVx2_ASAP7_75t_L g489 ( .A(n_487), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_489), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_489), .A2(n_507), .B(n_528), .C(n_529), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_494), .B(n_559), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_494), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
AND2x2_ASAP7_75t_L g584 ( .A(n_496), .B(n_559), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_496), .B(n_499), .Y(n_602) );
INVx1_ASAP7_75t_L g622 ( .A(n_496), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_496), .B(n_558), .Y(n_667) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_496), .Y(n_709) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_497), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_498), .B(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_498), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_498), .A2(n_554), .B(n_615), .C(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g621 ( .A(n_498), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g630 ( .A(n_498), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g634 ( .A(n_498), .B(n_558), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_498), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g649 ( .A(n_498), .B(n_559), .Y(n_649) );
AND2x2_ASAP7_75t_L g699 ( .A(n_498), .B(n_700), .Y(n_699) );
INVx5_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g563 ( .A(n_499), .Y(n_563) );
AND2x2_ASAP7_75t_L g604 ( .A(n_499), .B(n_557), .Y(n_604) );
AND2x2_ASAP7_75t_L g616 ( .A(n_499), .B(n_591), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_499), .B(n_645), .Y(n_663) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_508), .Y(n_499) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_531), .Y(n_510) );
INVx1_ASAP7_75t_L g552 ( .A(n_511), .Y(n_552) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
OR2x2_ASAP7_75t_L g554 ( .A(n_512), .B(n_523), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_512), .B(n_561), .C(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_512), .B(n_533), .Y(n_571) );
OR2x2_ASAP7_75t_L g586 ( .A(n_512), .B(n_574), .Y(n_586) );
AND2x2_ASAP7_75t_L g592 ( .A(n_512), .B(n_542), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_512), .B(n_723), .Y(n_722) );
INVx5_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_513), .B(n_533), .Y(n_589) );
AND2x2_ASAP7_75t_L g628 ( .A(n_513), .B(n_543), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_513), .B(n_542), .Y(n_656) );
OR2x2_ASAP7_75t_L g659 ( .A(n_513), .B(n_542), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVx5_ASAP7_75t_SL g574 ( .A(n_523), .Y(n_574) );
OR2x2_ASAP7_75t_L g580 ( .A(n_523), .B(n_532), .Y(n_580) );
AND2x2_ASAP7_75t_L g596 ( .A(n_523), .B(n_597), .Y(n_596) );
AOI321xp33_ASAP7_75t_L g603 ( .A1(n_523), .A2(n_604), .A3(n_605), .B1(n_606), .B2(n_612), .C(n_614), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_523), .B(n_531), .Y(n_613) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_523), .Y(n_626) );
OR2x2_ASAP7_75t_L g673 ( .A(n_523), .B(n_571), .Y(n_673) );
AND2x2_ASAP7_75t_L g695 ( .A(n_523), .B(n_592), .Y(n_695) );
AND2x2_ASAP7_75t_L g714 ( .A(n_523), .B(n_533), .Y(n_714) );
OR2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_530), .Y(n_523) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_542), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_533), .B(n_542), .Y(n_555) );
AND2x2_ASAP7_75t_L g564 ( .A(n_533), .B(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g591 ( .A(n_533), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_533), .B(n_592), .Y(n_597) );
INVxp67_ASAP7_75t_L g627 ( .A(n_533), .Y(n_627) );
OR2x2_ASAP7_75t_L g669 ( .A(n_533), .B(n_574), .Y(n_669) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_541), .Y(n_533) );
OR2x2_ASAP7_75t_L g551 ( .A(n_542), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g565 ( .A(n_542), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_542), .B(n_554), .Y(n_598) );
AND2x2_ASAP7_75t_L g647 ( .A(n_542), .B(n_591), .Y(n_647) );
AND2x2_ASAP7_75t_L g685 ( .A(n_542), .B(n_574), .Y(n_685) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_543), .B(n_574), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B(n_556), .C(n_560), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_551), .A2(n_553), .B1(n_678), .B2(n_680), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_553), .A2(n_576), .B1(n_631), .B2(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_SL g705 ( .A(n_554), .Y(n_705) );
INVx1_ASAP7_75t_SL g605 ( .A(n_555), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_557), .B(n_577), .Y(n_607) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_557), .A2(n_598), .B1(n_605), .B2(n_619), .C1(n_623), .C2(n_629), .Y(n_618) );
AND2x2_ASAP7_75t_L g708 ( .A(n_557), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g583 ( .A(n_558), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_558), .B(n_578), .Y(n_653) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_558), .Y(n_690) );
AND2x2_ASAP7_75t_L g693 ( .A(n_558), .B(n_602), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_558), .B(n_709), .Y(n_719) );
INVx1_ASAP7_75t_L g610 ( .A(n_559), .Y(n_610) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_559), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g701 ( .A1(n_561), .A2(n_702), .B(n_703), .C(n_706), .Y(n_701) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_563), .B(n_625), .C(n_628), .Y(n_624) );
OR2x2_ASAP7_75t_L g652 ( .A(n_563), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_563), .B(n_579), .Y(n_680) );
OR2x2_ASAP7_75t_L g585 ( .A(n_565), .B(n_586), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B(n_575), .C(n_587), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_568), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g674 ( .A(n_569), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_570), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g588 ( .A(n_573), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_574), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g642 ( .A(n_574), .B(n_592), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_574), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_574), .B(n_591), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_580), .B1(n_581), .B2(n_585), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_577), .B(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_579), .B(n_621), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_580), .A2(n_644), .B1(n_646), .B2(n_648), .C(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g698 ( .A(n_583), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g711 ( .A(n_583), .B(n_700), .Y(n_711) );
INVx1_ASAP7_75t_L g631 ( .A(n_584), .Y(n_631) );
INVx1_ASAP7_75t_L g702 ( .A(n_585), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_586), .A2(n_669), .B(n_692), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_590), .B(n_593), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_598), .B(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g635 ( .A(n_596), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_597), .A2(n_683), .B1(n_686), .B2(n_688), .C(n_691), .Y(n_682) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_605), .A2(n_695), .B1(n_696), .B2(n_698), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g671 ( .A(n_607), .Y(n_671) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp67_ASAP7_75t_SL g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g675 ( .A(n_611), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g640 ( .A(n_616), .Y(n_640) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_621), .B(n_645), .Y(n_697) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_627), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g713 ( .A(n_628), .B(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g720 ( .A(n_628), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_635), .B(n_636), .C(n_670), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_643), .C(n_662), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g723 ( .A(n_647), .Y(n_723) );
AND2x2_ASAP7_75t_L g660 ( .A(n_649), .B(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_658), .B2(n_660), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
OR2x2_ASAP7_75t_L g668 ( .A(n_656), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g721 ( .A(n_657), .Y(n_721) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI31xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .A3(n_665), .B(n_668), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_674), .C(n_677), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
NAND5xp2_ASAP7_75t_L g681 ( .A(n_682), .B(n_694), .C(n_701), .D(n_715), .E(n_718), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_693), .A2(n_719), .B1(n_720), .B2(n_722), .Y(n_718) );
INVx1_ASAP7_75t_SL g717 ( .A(n_695), .Y(n_717) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B(n_712), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
CKINVDCx14_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
CKINVDCx6p67_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g749 ( .A(n_743), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_747), .Y(n_743) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule