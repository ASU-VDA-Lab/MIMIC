module fake_jpeg_27675_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_2),
.B(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_24),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_13),
.B1(n_15),
.B2(n_22),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_18),
.B1(n_16),
.B2(n_24),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_25),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_60),
.Y(n_65)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_43),
.B1(n_44),
.B2(n_25),
.Y(n_76)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_59),
.B1(n_49),
.B2(n_32),
.Y(n_63)
);

BUFx2_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_15),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_40),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_69),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_44),
.B(n_41),
.C(n_43),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_76),
.B1(n_51),
.B2(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_39),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_60),
.B(n_52),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_42),
.C(n_33),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_44),
.Y(n_77)
);

NOR4xp25_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_73),
.C(n_70),
.D(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_85),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_49),
.B1(n_33),
.B2(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_30),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_66),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_95),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_97),
.B(n_84),
.C(n_14),
.D(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_64),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_66),
.B(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR4xp25_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_16),
.C(n_22),
.D(n_14),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_84),
.C(n_86),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_82),
.C(n_33),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_93),
.B(n_14),
.C(n_17),
.D(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_105),
.C(n_108),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_28),
.C(n_30),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_28),
.C(n_14),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_113),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_89),
.B(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_10),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_100),
.C(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_121),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_1),
.B(n_2),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_9),
.A3(n_12),
.B1(n_8),
.B2(n_14),
.C1(n_6),
.C2(n_7),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_109),
.B1(n_49),
.B2(n_21),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_12),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_115),
.Y(n_124)
);

OAI222xp33_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_116),
.B1(n_5),
.B2(n_6),
.C1(n_3),
.C2(n_20),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_128),
.B(n_21),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_5),
.B(n_20),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_5),
.B(n_20),
.C(n_21),
.D(n_26),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_26),
.B2(n_28),
.Y(n_131)
);


endmodule