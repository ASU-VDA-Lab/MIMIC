module real_jpeg_20407_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_41),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_1),
.A2(n_11),
.B(n_23),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_103),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_1),
.A2(n_30),
.B1(n_113),
.B2(n_114),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_37),
.B1(n_42),
.B2(n_75),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_37),
.B1(n_42),
.B2(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_59),
.Y(n_96)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_8),
.A2(n_37),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_51),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_11),
.A2(n_34),
.B(n_55),
.C(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_34),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_12),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_87)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_89),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_62),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_18),
.B(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.C(n_52),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_19),
.A2(n_20),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_33),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_29),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_22),
.B(n_27),
.Y(n_130)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_25),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_26),
.B(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_26),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_28),
.A2(n_96),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_30),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_30),
.B(n_103),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

AOI32xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.A3(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_39),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_35),
.A2(n_57),
.B(n_103),
.C(n_104),
.Y(n_102)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_42),
.B(n_47),
.C(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_60),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_54),
.A2(n_56),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_103),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_82),
.B2(n_83),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_132),
.B(n_137),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_121),
.B(n_131),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_109),
.B(n_120),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_114),
.B(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_115),
.B(n_119),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_128),
.C(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);


endmodule