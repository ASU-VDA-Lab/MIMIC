module fake_jpeg_17465_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_1),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_36),
.B1(n_5),
.B2(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_44),
.C(n_41),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_76),
.B(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_79),
.B1(n_70),
.B2(n_12),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_71),
.B1(n_7),
.B2(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_73),
.C(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_75),
.C(n_14),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_3),
.B(n_16),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_89),
.C(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_18),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_20),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_25),
.B(n_26),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_27),
.C(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_32),
.Y(n_99)
);


endmodule