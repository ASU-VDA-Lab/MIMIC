module fake_jpeg_26678_n_66 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_66);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_66;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_32),
.B(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_32)
);

OAI221xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_4),
.C(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_45),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_25),
.B1(n_28),
.B2(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_6),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_4),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_28),
.C(n_25),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_39),
.C(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_53),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AOI22x1_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_16),
.B1(n_8),
.B2(n_10),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_60),
.B(n_49),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_52),
.B1(n_51),
.B2(n_56),
.Y(n_61)
);

XNOR2x2_ASAP7_75t_SL g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_58),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_59),
.B(n_50),
.Y(n_65)
);

AOI221xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_66)
);


endmodule