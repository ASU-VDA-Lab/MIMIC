module real_jpeg_6602_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_1),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_1),
.B(n_118),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_2),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_2),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_3),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_3),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_3),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_3),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_4),
.B(n_162),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_4),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_4),
.B(n_406),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_5),
.B(n_40),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_5),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_5),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_6),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_6),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_6),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_6),
.B(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_6),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_6),
.B(n_381),
.Y(n_380)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_7),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_7),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_8),
.B(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_8),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_8),
.B(n_403),
.Y(n_402)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_10),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_10),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_10),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_10),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_10),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_10),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_10),
.B(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_11),
.Y(n_293)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_13),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_13),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_13),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_13),
.B(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_13),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_14),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_14),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_14),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_15),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_16),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_16),
.B(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_16),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_16),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_16),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_17),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_17),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_17),
.B(n_88),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_17),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_17),
.B(n_95),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_364),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_314),
.B(n_363),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_267),
.B(n_313),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_227),
.B(n_266),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_150),
.B(n_226),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_133),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_25),
.B(n_133),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_74),
.B2(n_132),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_26),
.B(n_75),
.C(n_115),
.Y(n_265)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_50),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_28),
.B(n_51),
.C(n_73),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.C(n_47),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_29),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_138)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_39),
.Y(n_143)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_42),
.B(n_47),
.Y(n_149)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_46),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_49),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_59),
.B1(n_72),
.B2(n_73),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B(n_58),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_54),
.Y(n_58)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_58),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_58),
.B(n_232),
.C(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_59),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.CI(n_68),
.CON(n_59),
.SN(n_59)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_60),
.B(n_63),
.C(n_68),
.Y(n_264)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_115),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_91),
.C(n_107),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_83),
.C(n_87),
.Y(n_131)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_81),
.Y(n_338)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_82),
.Y(n_252)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_86),
.Y(n_395)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_92),
.B1(n_107),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_103),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_93),
.A2(n_94),
.B1(n_103),
.B2(n_104),
.Y(n_219)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_95),
.Y(n_390)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_96),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_97),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_102),
.Y(n_291)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_102),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_102),
.Y(n_406)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_109),
.B(n_400),
.Y(n_399)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_129),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_116),
.B(n_130),
.C(n_131),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_117),
.B(n_125),
.C(n_127),
.Y(n_243)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_120),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_121)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_148),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_134),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_137),
.B(n_148),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.C(n_141),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_139),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_141),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_144),
.Y(n_190)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_146),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_221),
.B(n_225),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_206),
.B(n_220),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_187),
.B(n_205),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_175),
.B(n_186),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_163),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_158),
.Y(n_304)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_158),
.Y(n_330)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_167),
.C(n_170),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_173),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_181),
.B(n_185),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_179),
.Y(n_346)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_204),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_204),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_191),
.C(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_199),
.C(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_216),
.C(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_265),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_265),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_245),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_231),
.C(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_242),
.B2(n_244),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_248),
.C(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_252),
.Y(n_296)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g400 ( 
.A(n_256),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_261),
.C(n_264),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_269),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_270),
.B(n_286),
.C(n_311),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_286),
.B1(n_311),
.B2(n_312),
.Y(n_271)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_285),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_316)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_279),
.B(n_280),
.C(n_284),
.Y(n_352)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_297),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_298),
.C(n_299),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_287),
.Y(n_412)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_292),
.CI(n_294),
.CON(n_287),
.SN(n_287)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_288),
.B(n_292),
.C(n_294),
.Y(n_360)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_308),
.B2(n_309),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_307),
.C(n_308),
.Y(n_332)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_307),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_321),
.C(n_326),
.Y(n_378)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_362),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_362),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_316),
.B(n_318),
.C(n_348),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_348),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_331),
.B2(n_347),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_319),
.B(n_332),
.C(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_325),
.A2(n_326),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_344),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_339),
.C(n_344),
.Y(n_397)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_361),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_352),
.C(n_353),
.Y(n_368)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_351),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_360),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_354)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_355),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_357),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_358),
.C(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_357),
.A2(n_359),
.B1(n_380),
.B2(n_384),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_409),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_408),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_408),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_385),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_380),
.Y(n_384)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_396),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_404),
.B1(n_405),
.B2(n_407),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_402),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_405),
.Y(n_404)
);


endmodule