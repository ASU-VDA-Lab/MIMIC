module fake_netlist_5_1193_n_653 (n_137, n_91, n_82, n_122, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_653);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_653;

wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_483;
wire n_544;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_48),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_10),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_25),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_39),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_5),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_9),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_55),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_110),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_38),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_35),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_20),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_90),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_28),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_49),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_29),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_138),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_84),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_24),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_14),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_80),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_77),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_109),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_67),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_68),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_37),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_54),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_50),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_12),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_103),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_125),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_60),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_0),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_0),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_1),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_1),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_2),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_153),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_144),
.B(n_3),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_153),
.B(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_144),
.B(n_4),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_4),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_159),
.B(n_5),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_6),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_147),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_185),
.B(n_6),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_7),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_163),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_178),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_182),
.B(n_8),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_8),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_142),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_184),
.B(n_9),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_187),
.B(n_11),
.Y(n_256)
);

CKINVDCx6p67_ASAP7_75t_R g257 ( 
.A(n_209),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_209),
.B1(n_186),
.B2(n_143),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_217),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_214),
.A2(n_189),
.B1(n_195),
.B2(n_204),
.Y(n_260)
);

BUFx6f_ASAP7_75t_SL g261 ( 
.A(n_228),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_196),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_150),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_218),
.B1(n_223),
.B2(n_219),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_241),
.B1(n_226),
.B2(n_224),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_199),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_218),
.A2(n_143),
.B1(n_201),
.B2(n_203),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_214),
.A2(n_202),
.B1(n_207),
.B2(n_210),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_211),
.B(n_11),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_198),
.B1(n_197),
.B2(n_194),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_151),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_193),
.B1(n_192),
.B2(n_191),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_13),
.B1(n_14),
.B2(n_190),
.Y(n_276)
);

AO22x2_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_13),
.B1(n_188),
.B2(n_181),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_155),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_175),
.B1(n_174),
.B2(n_173),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_241),
.A2(n_167),
.B1(n_166),
.B2(n_165),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_158),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_170),
.B1(n_162),
.B2(n_161),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_16),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_253),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_226),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_230),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_238),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_212),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_229),
.B(n_46),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_229),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_212),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_291)
);

AO22x2_ASAP7_75t_L g292 ( 
.A1(n_243),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_220),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_R g296 ( 
.A(n_257),
.B(n_72),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_230),
.A2(n_73),
.B1(n_74),
.B2(n_78),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_250),
.A2(n_79),
.B1(n_81),
.B2(n_85),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_R g301 ( 
.A1(n_220),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_231),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_97),
.B1(n_98),
.B2(n_101),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_243),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_256),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_237),
.B(n_117),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

AO22x2_ASAP7_75t_L g308 ( 
.A1(n_244),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_237),
.B(n_123),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_269),
.B(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_293),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_274),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_237),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_266),
.Y(n_319)
);

XNOR2x2_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_231),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_270),
.B(n_127),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_258),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_213),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_213),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_267),
.B(n_128),
.Y(n_341)
);

NAND2x1p5_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_240),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g344 ( 
.A(n_301),
.B(n_249),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_245),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_260),
.B(n_247),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_262),
.B(n_213),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_277),
.B(n_129),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_277),
.B(n_130),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

OR2x2_ASAP7_75t_SL g357 ( 
.A(n_261),
.B(n_225),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_296),
.B(n_222),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_286),
.B(n_247),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_273),
.B(n_235),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_268),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_279),
.B(n_247),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_282),
.B(n_221),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_259),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_259),
.B(n_254),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_259),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_271),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_259),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_259),
.B(n_254),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_259),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_259),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_259),
.B(n_254),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_254),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_373),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_252),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_252),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_330),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_310),
.B(n_252),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_252),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_248),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_359),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_310),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_344),
.B(n_248),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_248),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_349),
.B(n_242),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_313),
.B(n_359),
.Y(n_404)
);

NAND2x1p5_ASAP7_75t_L g405 ( 
.A(n_350),
.B(n_247),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_324),
.B(n_246),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_246),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_321),
.B(n_131),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_246),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_246),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_248),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_313),
.B(n_242),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_242),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_236),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVx3_ASAP7_75t_SL g419 ( 
.A(n_357),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_366),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_365),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_364),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_345),
.B(n_349),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_345),
.B(n_347),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_319),
.B(n_236),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_319),
.B(n_236),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_363),
.B(n_233),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_316),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_342),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_344),
.B(n_333),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_415),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_334),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_439),
.Y(n_444)
);

BUFx8_ASAP7_75t_SL g445 ( 
.A(n_394),
.Y(n_445)
);

NAND2x1p5_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_336),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_433),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_397),
.B(n_360),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_417),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_331),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_326),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_408),
.B(n_335),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_343),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_348),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_348),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_348),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_346),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_432),
.Y(n_463)
);

BUFx12f_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_413),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_408),
.B(n_354),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_320),
.Y(n_467)
);

INVx3_ASAP7_75t_SL g468 ( 
.A(n_419),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_421),
.B(n_356),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_358),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_378),
.B(n_132),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_361),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_391),
.Y(n_476)
);

AO21x2_ASAP7_75t_L g477 ( 
.A1(n_406),
.A2(n_327),
.B(n_353),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_438),
.B(n_352),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_426),
.B(n_361),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_379),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_424),
.B(n_361),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_361),
.Y(n_484)
);

INVx5_ASAP7_75t_SL g485 ( 
.A(n_482),
.Y(n_485)
);

BUFx12f_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_452),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_395),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

NAND2x1p5_ASAP7_75t_L g492 ( 
.A(n_444),
.B(n_383),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_444),
.B(n_383),
.Y(n_493)
);

NAND2x1p5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_378),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_448),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_458),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_481),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_474),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_484),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_445),
.Y(n_503)
);

BUFx2_ASAP7_75t_SL g504 ( 
.A(n_476),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_476),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_464),
.Y(n_506)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_469),
.B(n_395),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_442),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_468),
.Y(n_511)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_483),
.Y(n_513)
);

INVx3_ASAP7_75t_SL g514 ( 
.A(n_468),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_469),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_455),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_508),
.A2(n_397),
.B1(n_449),
.B2(n_455),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_501),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_503),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_501),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_456),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_502),
.A2(n_449),
.B1(n_443),
.B2(n_341),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_503),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_502),
.A2(n_361),
.B1(n_453),
.B2(n_403),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_467),
.B1(n_328),
.B2(n_479),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_510),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_495),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_510),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_513),
.A2(n_480),
.B1(n_475),
.B2(n_454),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_496),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_496),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_456),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_497),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_499),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_489),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_499),
.A2(n_454),
.B1(n_402),
.B2(n_436),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_465),
.Y(n_537)
);

BUFx2_ASAP7_75t_SL g538 ( 
.A(n_506),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_509),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_509),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_494),
.A2(n_466),
.B1(n_456),
.B2(n_446),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_516),
.A2(n_461),
.B(n_459),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_525),
.A2(n_328),
.B1(n_477),
.B2(n_479),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_522),
.A2(n_466),
.B1(n_504),
.B2(n_505),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_531),
.Y(n_546)
);

BUFx12f_ASAP7_75t_L g547 ( 
.A(n_540),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_525),
.A2(n_517),
.B(n_522),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

AOI222xp33_ASAP7_75t_L g550 ( 
.A1(n_515),
.A2(n_462),
.B1(n_440),
.B2(n_466),
.C1(n_393),
.C2(n_454),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_519),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_534),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_517),
.A2(n_477),
.B1(n_479),
.B2(n_529),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_523),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_518),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_520),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_533),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_541),
.A2(n_479),
.B1(n_404),
.B2(n_414),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_540),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_526),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_529),
.A2(n_436),
.B1(n_396),
.B2(n_462),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_536),
.A2(n_485),
.B1(n_377),
.B2(n_398),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_536),
.A2(n_380),
.B(n_511),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_535),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_521),
.A2(n_473),
.B(n_386),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_521),
.A2(n_396),
.B1(n_478),
.B2(n_457),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_524),
.A2(n_485),
.B1(n_377),
.B2(n_500),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_532),
.A2(n_418),
.B1(n_420),
.B2(n_387),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_535),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_532),
.A2(n_418),
.B1(n_420),
.B2(n_387),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_548),
.B(n_537),
.Y(n_573)
);

AOI221xp5_ASAP7_75t_L g574 ( 
.A1(n_544),
.A2(n_399),
.B1(n_457),
.B2(n_412),
.C(n_388),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_544),
.A2(n_396),
.B1(n_499),
.B2(n_500),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_545),
.A2(n_538),
.B1(n_473),
.B2(n_512),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_565),
.A2(n_524),
.B1(n_514),
.B2(n_485),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_564),
.A2(n_512),
.B1(n_507),
.B2(n_486),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_553),
.A2(n_396),
.B1(n_499),
.B2(n_500),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_553),
.A2(n_396),
.B1(n_499),
.B2(n_500),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_559),
.A2(n_396),
.B1(n_500),
.B2(n_491),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_555),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_570),
.A2(n_514),
.B1(n_485),
.B2(n_506),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_572),
.A2(n_472),
.B1(n_507),
.B2(n_486),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_550),
.A2(n_512),
.B1(n_376),
.B2(n_472),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_569),
.A2(n_512),
.B1(n_446),
.B2(n_472),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_546),
.A2(n_382),
.B1(n_392),
.B2(n_400),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_543),
.B(n_534),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_558),
.A2(n_390),
.B1(n_478),
.B2(n_381),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_543),
.A2(n_494),
.B1(n_534),
.B2(n_442),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_556),
.B(n_557),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_567),
.A2(n_539),
.B1(n_401),
.B2(n_450),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_563),
.A2(n_450),
.B1(n_498),
.B2(n_488),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_563),
.A2(n_450),
.B1(n_498),
.B2(n_488),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_549),
.A2(n_460),
.B1(n_534),
.B2(n_405),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_592),
.A2(n_568),
.B1(n_549),
.B2(n_560),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_573),
.A2(n_578),
.B1(n_589),
.B2(n_585),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_584),
.A2(n_576),
.B(n_583),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_577),
.A2(n_547),
.B1(n_542),
.B2(n_568),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_571),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_588),
.B(n_566),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_562),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_575),
.B(n_561),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_581),
.A2(n_405),
.B(n_450),
.Y(n_604)
);

NAND4xp25_ASAP7_75t_L g605 ( 
.A(n_574),
.B(n_437),
.C(n_416),
.D(n_552),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_552),
.C(n_416),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_590),
.B(n_527),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_594),
.C(n_586),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_579),
.B(n_554),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_580),
.A2(n_451),
.B1(n_430),
.B2(n_379),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_598),
.B(n_595),
.C(n_406),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_595),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_602),
.Y(n_613)
);

NOR3xp33_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_407),
.C(n_409),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_600),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_603),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_608),
.B(n_607),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_616),
.B(n_609),
.Y(n_620)
);

NAND4xp75_ASAP7_75t_SL g621 ( 
.A(n_611),
.B(n_599),
.C(n_597),
.D(n_596),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_613),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_615),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_617),
.B(n_606),
.C(n_407),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_617),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_622),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_623),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_612),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_621),
.B(n_551),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_625),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_626),
.Y(n_631)
);

CKINVDCx8_ASAP7_75t_R g632 ( 
.A(n_629),
.Y(n_632)
);

OA22x2_ASAP7_75t_L g633 ( 
.A1(n_626),
.A2(n_619),
.B1(n_621),
.B2(n_624),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_627),
.Y(n_634)
);

OA22x2_ASAP7_75t_L g635 ( 
.A1(n_630),
.A2(n_614),
.B1(n_445),
.B2(n_451),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_634),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_631),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_633),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_637),
.B(n_635),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_638),
.A2(n_628),
.B1(n_632),
.B2(n_610),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_639),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_638),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_642),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_640),
.B1(n_636),
.B2(n_610),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_644),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_429),
.B1(n_493),
.B2(n_492),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_646),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_430),
.B1(n_429),
.B2(n_411),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_648),
.Y(n_649)
);

AO22x2_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_430),
.B1(n_409),
.B2(n_444),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_650),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_L g652 ( 
.A1(n_651),
.A2(n_134),
.B1(n_139),
.B2(n_463),
.C(n_470),
.Y(n_652)
);

AOI211xp5_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_411),
.B(n_463),
.C(n_470),
.Y(n_653)
);


endmodule