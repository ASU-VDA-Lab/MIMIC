module fake_jpeg_5689_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_34),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_29),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_16),
.B1(n_24),
.B2(n_22),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_43),
.B1(n_15),
.B2(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_51),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_24),
.B1(n_16),
.B2(n_27),
.Y(n_41)
);

OA22x2_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_33),
.B1(n_17),
.B2(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_22),
.B1(n_28),
.B2(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_47),
.Y(n_56)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_30),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_60),
.B(n_48),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_57),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_64),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_36),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_66),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_37),
.B(n_33),
.C(n_35),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_71),
.B1(n_73),
.B2(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_15),
.B1(n_17),
.B2(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_95),
.Y(n_98)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_33),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_64),
.C(n_67),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_53),
.B1(n_47),
.B2(n_4),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_42),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_52),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_1),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_71),
.B1(n_54),
.B2(n_72),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_97),
.B1(n_108),
.B2(n_88),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_72),
.B1(n_62),
.B2(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_105),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_87),
.B(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_113),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_47),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_R g122 ( 
.A(n_106),
.B(n_109),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_77),
.B(n_114),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_85),
.B(n_89),
.C(n_109),
.D(n_76),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_110),
.B(n_101),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_81),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_126),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_91),
.B1(n_80),
.B2(n_84),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_103),
.B1(n_111),
.B2(n_106),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_76),
.C(n_78),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_97),
.C(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_98),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_140),
.C(n_143),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_128),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_125),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_2),
.C(n_3),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_120),
.B(n_121),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_143),
.B(n_4),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_127),
.C(n_118),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_153),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2x1_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_160),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_134),
.B(n_139),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_3),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_144),
.C(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_165),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_152),
.B1(n_144),
.B2(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_161),
.B(n_6),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_170),
.B(n_164),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_3),
.B(n_8),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_162),
.C(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_167),
.C(n_170),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);


endmodule