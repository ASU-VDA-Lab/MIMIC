module fake_jpeg_22563_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_40),
.B(n_45),
.Y(n_84)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_61),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_29),
.B1(n_27),
.B2(n_36),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_66),
.A2(n_77),
.B1(n_28),
.B2(n_4),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_36),
.B1(n_30),
.B2(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_28),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_36),
.B1(n_32),
.B2(n_23),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_75),
.B1(n_38),
.B2(n_37),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_32),
.B1(n_23),
.B2(n_20),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_2),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_34),
.B(n_24),
.C(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_32),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_20),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_35),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_104),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_91),
.B(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_106),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_34),
.B1(n_21),
.B2(n_22),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_93),
.A2(n_95),
.B1(n_121),
.B2(n_69),
.Y(n_154)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_38),
.CON(n_94),
.SN(n_94)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_97),
.B(n_3),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_34),
.B1(n_21),
.B2(n_22),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_108),
.Y(n_125)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_34),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_64),
.A3(n_77),
.B1(n_59),
.B2(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_102),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_62),
.A2(n_19),
.B1(n_33),
.B2(n_35),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_33),
.B1(n_18),
.B2(n_25),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_25),
.B1(n_28),
.B2(n_5),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_3),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_134),
.C(n_102),
.Y(n_161)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_123),
.A2(n_136),
.B1(n_138),
.B2(n_76),
.Y(n_181)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_126),
.Y(n_170)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_130),
.Y(n_173)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_132),
.B(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_83),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_71),
.C(n_56),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_85),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_141),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_53),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

CKINVDCx11_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_92),
.B(n_53),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_89),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_103),
.B1(n_95),
.B2(n_93),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_70),
.B1(n_65),
.B2(n_69),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_107),
.B1(n_121),
.B2(n_96),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_61),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_95),
.B1(n_118),
.B2(n_93),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_181),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_101),
.B(n_108),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_158),
.A2(n_160),
.B(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_91),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_159),
.B(n_183),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_99),
.B(n_109),
.C(n_93),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_110),
.B(n_94),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_143),
.B(n_5),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_185),
.B(n_135),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_103),
.C(n_98),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_152),
.C(n_149),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_135),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_171),
.A2(n_177),
.B1(n_179),
.B2(n_8),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_63),
.B1(n_118),
.B2(n_95),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_186),
.B1(n_138),
.B2(n_123),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_113),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_137),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_145),
.B1(n_129),
.B2(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_124),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_125),
.A2(n_113),
.B(n_82),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_127),
.A2(n_76),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_202),
.C(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_157),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_122),
.B1(n_153),
.B2(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_189),
.A2(n_198),
.B1(n_157),
.B2(n_168),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_182),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_196),
.B(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_171),
.B1(n_161),
.B2(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_176),
.B(n_159),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_143),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_128),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_126),
.C(n_130),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_175),
.C(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_169),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_155),
.B(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_168),
.B1(n_163),
.B2(n_10),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_6),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_186),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_160),
.B1(n_172),
.B2(n_162),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_217),
.B(n_231),
.Y(n_243)
);

NOR3xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_176),
.C(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_205),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_156),
.B(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_223),
.C(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_233),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_235),
.B1(n_207),
.B2(n_192),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_160),
.B(n_162),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_213),
.B1(n_189),
.B2(n_200),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_199),
.B1(n_209),
.B2(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_239),
.B1(n_248),
.B2(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_202),
.C(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_244),
.C(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_232),
.C(n_214),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_196),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_250),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_247),
.B(n_253),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_195),
.B1(n_208),
.B2(n_187),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_203),
.C(n_201),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_163),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_262),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_229),
.B(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_268),
.C(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_230),
.C(n_218),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_261),
.C(n_245),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_223),
.C(n_217),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_220),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_265),
.B1(n_241),
.B2(n_249),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_233),
.B(n_212),
.C(n_10),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_266),
.A2(n_255),
.B1(n_264),
.B2(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_265),
.B1(n_11),
.B2(n_12),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_267),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_275),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_243),
.C(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_278),
.C(n_8),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_245),
.C(n_9),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_261),
.B1(n_265),
.B2(n_12),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_284),
.B1(n_13),
.B2(n_14),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_270),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_8),
.B(n_13),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_13),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_14),
.Y(n_293)
);

AOI31xp33_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_275),
.A3(n_272),
.B(n_279),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_290),
.Y(n_297)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_285),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_284),
.C(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_287),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_294),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_290),
.C(n_282),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_297),
.B(n_280),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_302),
.A2(n_303),
.B(n_301),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_296),
.B(n_297),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_286),
.Y(n_306)
);


endmodule