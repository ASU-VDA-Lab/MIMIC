module fake_netlist_5_1520_n_2241 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2241);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2241;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_1070;
wire n_777;
wire n_422;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_832;
wire n_857;
wire n_1319;
wire n_561;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_1138;
wire n_364;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_91),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_61),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_206),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_93),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_89),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_124),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_29),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_36),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_85),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_60),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_61),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_39),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_86),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_66),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_14),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_199),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_168),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_103),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_144),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_113),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_65),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_17),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_202),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_139),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_99),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_170),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_28),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_220),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_90),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_131),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_51),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_92),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_80),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_79),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_108),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_142),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_48),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_159),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_138),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_167),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_218),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_65),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_45),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_201),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_15),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_72),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_7),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_2),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_49),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_122),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_52),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_109),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_143),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_106),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_75),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_47),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_77),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_51),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_78),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_178),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_1),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_7),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_59),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_33),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_39),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_70),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_135),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_105),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_62),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_125),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_79),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_175),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_116),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_76),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_213),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_120),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_47),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_173),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_10),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_211),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_76),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_43),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_69),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_186),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_62),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_34),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_136),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_49),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_190),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_189),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_183),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_31),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_38),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_101),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_171),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_45),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_81),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_179),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_82),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_18),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_191),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_31),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_149),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_25),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_148),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_3),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_214),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_57),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_196),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_204),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_36),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_14),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_57),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_117),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_132),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_182),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_22),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_26),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_70),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_5),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_210),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_37),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_94),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_66),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_12),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_84),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_67),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_165),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_118),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_19),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_153),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_63),
.Y(n_383)
);

BUFx8_ASAP7_75t_SL g384 ( 
.A(n_185),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_133),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_21),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_137),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_46),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_87),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_126),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_19),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_98),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_97),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_27),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_11),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_187),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_1),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_68),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_197),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_188),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_41),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_58),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_44),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_27),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_176),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_75),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_25),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_151),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_88),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_69),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_102),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_29),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_184),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_172),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_41),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_205),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_23),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_194),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_11),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_53),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_83),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_77),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_141),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_110),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_56),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_181),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_64),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_78),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_53),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_163),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_52),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_111),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_34),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_74),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_30),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_154),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_259),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_290),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_384),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_259),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_277),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_324),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_240),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_277),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_296),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_296),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_222),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_225),
.Y(n_450)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_290),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_240),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_228),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_319),
.B(n_0),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_243),
.B(n_0),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_231),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_234),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_226),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_272),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_251),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_308),
.B(n_2),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_252),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_243),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_265),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_307),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_230),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_308),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_230),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_235),
.B(n_3),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_265),
.B(n_4),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_268),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_350),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_268),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_255),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_269),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_269),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_411),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_260),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_262),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_275),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_423),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_275),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_235),
.B(n_253),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_263),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_232),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_288),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_288),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_264),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_229),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_270),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_293),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_274),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_253),
.B(n_4),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_271),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_346),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_293),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_280),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_304),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_304),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_319),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_305),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_305),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_310),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_400),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_310),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_256),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_311),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_311),
.Y(n_510)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_326),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_284),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_285),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_372),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_372),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_286),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_297),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_299),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_326),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_237),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_239),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_300),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_292),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_301),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_336),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_315),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_316),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_336),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_347),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_347),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_318),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_351),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_351),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_348),
.B(n_5),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_320),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_322),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_325),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_329),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_355),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_424),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_348),
.B(n_6),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_292),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_331),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_416),
.B(n_6),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_335),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_340),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_341),
.Y(n_548)
);

INVxp33_ASAP7_75t_SL g549 ( 
.A(n_242),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_342),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_355),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_244),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_352),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_485),
.B(n_416),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_515),
.B(n_358),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_508),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_508),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_466),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_466),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_508),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_508),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_454),
.B(n_408),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_515),
.B(n_436),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_470),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_487),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_514),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_437),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_437),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_454),
.B(n_541),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_440),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_502),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_441),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_523),
.B(n_292),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_536),
.B(n_408),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_444),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_445),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_536),
.B(n_408),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_446),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_495),
.B(n_261),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_521),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_458),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_471),
.B(n_534),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_463),
.B(n_542),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_448),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_443),
.B(n_232),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_545),
.B(n_224),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_520),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_475),
.B(n_360),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_452),
.B(n_236),
.Y(n_604)
);

BUFx8_ASAP7_75t_L g605 ( 
.A(n_521),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_475),
.B(n_477),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_449),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_469),
.B(n_449),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_477),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_460),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_462),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_478),
.B(n_261),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_462),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_478),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_482),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_482),
.Y(n_617)
);

AND2x2_ASAP7_75t_SL g618 ( 
.A(n_455),
.B(n_295),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_484),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_488),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_549),
.B(n_227),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_489),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_489),
.B(n_236),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_493),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_493),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_552),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_498),
.B(n_295),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_472),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_498),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_500),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_500),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_501),
.A2(n_368),
.B(n_363),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_501),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_503),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_503),
.B(n_238),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_505),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_524),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_507),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_438),
.A2(n_451),
.B1(n_472),
.B2(n_233),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_507),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_509),
.B(n_338),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_635),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_585),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_635),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_597),
.B(n_447),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_635),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_635),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_640),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_635),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_635),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_583),
.B(n_491),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_635),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_635),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_558),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_583),
.B(n_523),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_583),
.B(n_543),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_597),
.B(n_450),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_596),
.B(n_442),
.C(n_465),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_634),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_592),
.B(n_338),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_564),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_643),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_622),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_618),
.A2(n_317),
.B1(n_368),
.B2(n_363),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_622),
.B(n_453),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_634),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_591),
.B(n_238),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_600),
.B(n_457),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_634),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_643),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_564),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_600),
.B(n_461),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_585),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_575),
.B(n_464),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_582),
.B(n_476),
.Y(n_680)
);

INVxp33_ASAP7_75t_L g681 ( 
.A(n_579),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_634),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_575),
.B(n_480),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_634),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_575),
.B(n_509),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_616),
.Y(n_686)
);

BUFx4f_ASAP7_75t_L g687 ( 
.A(n_592),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_625),
.B(n_241),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_643),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_592),
.B(n_256),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_643),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_582),
.B(n_481),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_591),
.B(n_486),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_558),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_616),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_643),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_564),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_596),
.B(n_490),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_591),
.B(n_492),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_591),
.B(n_494),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_643),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_643),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_558),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_591),
.B(n_499),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_572),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_616),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_617),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_617),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_617),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_591),
.B(n_512),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_558),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_630),
.B(n_513),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_564),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_619),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_558),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_585),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_630),
.B(n_510),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_589),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_630),
.B(n_516),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_643),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_517),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_630),
.B(n_518),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_619),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_589),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_630),
.B(n_522),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_619),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_564),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_640),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_556),
.B(n_527),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_573),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_579),
.B(n_543),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_573),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_627),
.Y(n_734)
);

AND3x2_ASAP7_75t_L g735 ( 
.A(n_593),
.B(n_245),
.C(n_241),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_593),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_627),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_593),
.Y(n_738)
);

AND2x6_ASAP7_75t_L g739 ( 
.A(n_592),
.B(n_256),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_594),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_628),
.B(n_531),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_627),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_631),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_618),
.A2(n_317),
.B1(n_376),
.B2(n_369),
.Y(n_744)
);

BUFx4f_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_605),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_628),
.B(n_535),
.Y(n_747)
);

BUFx4f_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_631),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_573),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_642),
.B(n_294),
.C(n_223),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_618),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_558),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_632),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_556),
.B(n_537),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_510),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_558),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_618),
.B(n_538),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_564),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_564),
.B(n_554),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_572),
.B(n_544),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_564),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_586),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_568),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_586),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_632),
.Y(n_767)
);

AOI21x1_ASAP7_75t_L g768 ( 
.A1(n_554),
.A2(n_246),
.B(n_245),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_565),
.B(n_547),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_594),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_608),
.B(n_519),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_599),
.A2(n_376),
.B1(n_402),
.B2(n_369),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_586),
.Y(n_773)
);

INVx4_ASAP7_75t_SL g774 ( 
.A(n_564),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_568),
.Y(n_775)
);

BUFx10_ASAP7_75t_L g776 ( 
.A(n_564),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_605),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_632),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_639),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_586),
.Y(n_780)
);

OR2x6_ASAP7_75t_L g781 ( 
.A(n_599),
.B(n_246),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_587),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_608),
.B(n_550),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_564),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_601),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_587),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_608),
.B(n_553),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_565),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_587),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_587),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_605),
.B(n_526),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_568),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_639),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_639),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_642),
.A2(n_370),
.B1(n_371),
.B2(n_254),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_620),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_620),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_588),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_588),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_605),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_646),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_654),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_753),
.B(n_605),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_646),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_698),
.B(n_601),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_677),
.B(n_439),
.C(n_602),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_760),
.B(n_247),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_673),
.B(n_602),
.C(n_599),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_716),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_760),
.B(n_604),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_705),
.B(n_604),
.Y(n_812)
);

AOI221xp5_ASAP7_75t_L g813 ( 
.A1(n_751),
.A2(n_511),
.B1(n_604),
.B2(n_504),
.C(n_525),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_753),
.A2(n_637),
.B1(n_625),
.B2(n_402),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_686),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_651),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_788),
.B(n_620),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_654),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_686),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_716),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_760),
.B(n_247),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_770),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_676),
.B(n_605),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_788),
.B(n_762),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_648),
.B(n_661),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_717),
.B(n_620),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_717),
.B(n_620),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_700),
.B(n_623),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_704),
.B(n_623),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_676),
.B(n_256),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_695),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_722),
.B(n_623),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_738),
.B(n_606),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_676),
.B(n_256),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_716),
.B(n_623),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_695),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_706),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_679),
.B(n_539),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_785),
.B(n_732),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_664),
.B(n_361),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_SL g841 ( 
.A1(n_795),
.A2(n_459),
.B1(n_467),
.B2(n_456),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_759),
.A2(n_548),
.B1(n_546),
.B2(n_497),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_718),
.B(n_623),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_676),
.B(n_432),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_651),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_718),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_718),
.B(n_625),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_724),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_683),
.B(n_496),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_736),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_736),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_676),
.B(n_432),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_724),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_724),
.B(n_637),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_662),
.B(n_559),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_728),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_678),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_706),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_729),
.B(n_637),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_791),
.B(n_659),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_707),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_707),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_662),
.B(n_506),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_678),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_756),
.B(n_769),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_784),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_757),
.B(n_559),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_708),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_757),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_712),
.B(n_584),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_719),
.B(n_584),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_685),
.B(n_771),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_721),
.B(n_584),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_746),
.B(n_560),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_708),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_783),
.B(n_282),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_740),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_709),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_655),
.Y(n_879)
);

INVx8_ASAP7_75t_L g880 ( 
.A(n_672),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_732),
.B(n_606),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_685),
.B(n_474),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_655),
.A2(n_563),
.B(n_576),
.C(n_560),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_709),
.B(n_584),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_714),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_676),
.B(n_432),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_771),
.B(n_681),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_787),
.B(n_399),
.Y(n_888)
);

O2A1O1Ixp5_ASAP7_75t_L g889 ( 
.A1(n_663),
.A2(n_644),
.B(n_629),
.C(n_266),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_714),
.B(n_584),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_723),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_697),
.B(n_432),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_781),
.A2(n_404),
.B1(n_412),
.B2(n_407),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_668),
.B(n_479),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_668),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_668),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_723),
.B(n_598),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_784),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_726),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_670),
.B(n_248),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_741),
.B(n_249),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_L g902 ( 
.A(n_664),
.B(n_365),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_659),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_660),
.B(n_563),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_726),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_734),
.B(n_598),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_734),
.B(n_598),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_L g908 ( 
.A(n_664),
.B(n_697),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_747),
.B(n_250),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_660),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_737),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_737),
.B(n_598),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_742),
.B(n_598),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_668),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_742),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_743),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_743),
.B(n_749),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_749),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_752),
.B(n_609),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_781),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_752),
.B(n_609),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_755),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_755),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_767),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_735),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_784),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_SL g927 ( 
.A(n_746),
.B(n_483),
.Y(n_927)
);

CKINVDCx11_ASAP7_75t_R g928 ( 
.A(n_800),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_776),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_781),
.B(n_404),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_767),
.B(n_609),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_778),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_663),
.A2(n_557),
.B(n_555),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_778),
.B(n_779),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_776),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_779),
.B(n_793),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_671),
.A2(n_407),
.B1(n_417),
.B2(n_412),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_793),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_680),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_697),
.B(n_432),
.Y(n_940)
);

OAI221xp5_ASAP7_75t_L g941 ( 
.A1(n_669),
.A2(n_744),
.B1(n_772),
.B2(n_781),
.C(n_795),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_781),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_671),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_794),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_794),
.B(n_609),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_674),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_674),
.B(n_609),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_796),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_688),
.B(n_576),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_682),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_693),
.B(n_258),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_796),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_697),
.B(n_568),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_688),
.B(n_610),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_777),
.B(n_410),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_682),
.B(n_629),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_684),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_797),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_797),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_684),
.A2(n_417),
.B(n_425),
.C(n_420),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_688),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_761),
.A2(n_710),
.B1(n_725),
.B2(n_699),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_692),
.B(n_610),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_688),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_799),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_672),
.A2(n_374),
.B1(n_380),
.B2(n_367),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_697),
.B(n_568),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_664),
.B(n_385),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_672),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_799),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_687),
.B(n_629),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_687),
.B(n_745),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_687),
.B(n_629),
.Y(n_973)
);

O2A1O1Ixp5_ASAP7_75t_L g974 ( 
.A1(n_825),
.A2(n_748),
.B(n_745),
.C(n_768),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_825),
.A2(n_748),
.B1(n_745),
.B2(n_672),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_929),
.A2(n_748),
.B(n_713),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_824),
.B(n_672),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_866),
.Y(n_978)
);

AO21x1_ASAP7_75t_L g979 ( 
.A1(n_962),
.A2(n_768),
.B(n_266),
.Y(n_979)
);

NOR2x1_ASAP7_75t_L g980 ( 
.A(n_865),
.B(n_435),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_929),
.A2(n_713),
.B(n_665),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_805),
.B(n_777),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_859),
.B(n_664),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_929),
.A2(n_713),
.B(n_665),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_929),
.A2(n_713),
.B(n_665),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_841),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_941),
.A2(n_425),
.B(n_429),
.C(n_420),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_812),
.B(n_664),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_935),
.A2(n_727),
.B(n_665),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_935),
.A2(n_763),
.B(n_727),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_872),
.B(n_664),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_960),
.A2(n_267),
.B(n_276),
.C(n_257),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_822),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_935),
.A2(n_763),
.B(n_727),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_889),
.A2(n_763),
.B(n_727),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_901),
.B(n_658),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_935),
.A2(n_763),
.B(n_697),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_814),
.A2(n_267),
.B1(n_276),
.B2(n_257),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_956),
.A2(n_647),
.B(n_645),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_901),
.B(n_658),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_909),
.B(n_658),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_933),
.A2(n_647),
.B(n_645),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_909),
.A2(n_433),
.B(n_429),
.C(n_278),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_887),
.B(n_624),
.Y(n_1004)
);

OAI21xp33_ASAP7_75t_L g1005 ( 
.A1(n_876),
.A2(n_281),
.B(n_273),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_860),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_815),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_815),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_971),
.A2(n_776),
.B(n_715),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_826),
.A2(n_650),
.B(n_649),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_973),
.A2(n_776),
.B(n_715),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_851),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_827),
.A2(n_650),
.B(n_649),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_972),
.A2(n_715),
.B(n_703),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_908),
.A2(n_715),
.B(n_703),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_866),
.B(n_774),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_937),
.A2(n_739),
.B1(n_690),
.B2(n_433),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_847),
.A2(n_715),
.B(n_703),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_819),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_854),
.A2(n_754),
.B(n_703),
.Y(n_1020)
);

AOI33xp33_ASAP7_75t_L g1021 ( 
.A1(n_813),
.A2(n_540),
.A3(n_519),
.B1(n_528),
.B2(n_529),
.B3(n_530),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_819),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_831),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_831),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_833),
.B(n_624),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_949),
.B(n_666),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_805),
.A2(n_888),
.B(n_876),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_866),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_814),
.A2(n_279),
.B1(n_289),
.B2(n_278),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_838),
.B(n_849),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_866),
.A2(n_289),
.B1(n_321),
.B2(n_279),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_954),
.B(n_666),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_836),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_953),
.A2(n_653),
.B(n_652),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_870),
.A2(n_754),
.B(n_703),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_879),
.B(n_666),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_809),
.B(n_694),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_836),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_888),
.A2(n_327),
.B(n_321),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_855),
.B(n_694),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_839),
.B(n_528),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_871),
.A2(n_758),
.B(n_754),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_873),
.A2(n_758),
.B(n_754),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_817),
.B(n_694),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_856),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_898),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_882),
.B(n_292),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_802),
.B(n_332),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_818),
.B(n_332),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_850),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_937),
.A2(n_345),
.B(n_349),
.C(n_327),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_837),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_881),
.B(n_332),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_946),
.B(n_950),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_946),
.B(n_711),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_835),
.A2(n_843),
.B(n_947),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_858),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_811),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_863),
.B(n_382),
.C(n_349),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_898),
.B(n_775),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_898),
.Y(n_1061)
);

OAI321xp33_ASAP7_75t_L g1062 ( 
.A1(n_893),
.A2(n_383),
.A3(n_405),
.B1(n_379),
.B2(n_414),
.C(n_377),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_828),
.A2(n_758),
.B(n_754),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_829),
.A2(n_758),
.B(n_765),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_858),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_950),
.B(n_711),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_957),
.B(n_711),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_861),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_877),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_904),
.B(n_838),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_816),
.Y(n_1071)
);

CKINVDCx8_ASAP7_75t_R g1072 ( 
.A(n_845),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_920),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_832),
.A2(n_943),
.B(n_934),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_953),
.A2(n_653),
.B(n_652),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_957),
.B(n_690),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_862),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_862),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_875),
.B(n_690),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_867),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_857),
.B(n_774),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_943),
.A2(n_758),
.B(n_765),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_951),
.A2(n_354),
.B(n_366),
.C(n_345),
.Y(n_1083)
);

AOI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_900),
.A2(n_863),
.B(n_951),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_898),
.B(n_774),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_849),
.B(n_332),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_903),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_917),
.A2(n_765),
.B(n_657),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_936),
.A2(n_765),
.B(n_657),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_926),
.A2(n_765),
.B(n_667),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_900),
.A2(n_366),
.B(n_377),
.C(n_354),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_910),
.B(n_283),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_868),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_884),
.A2(n_667),
.B(n_656),
.Y(n_1094)
);

OAI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_869),
.A2(n_291),
.B(n_287),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_891),
.B(n_690),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_926),
.A2(n_675),
.B(n_656),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_905),
.B(n_690),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_864),
.B(n_298),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_426),
.B(n_379),
.C(n_430),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_926),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_915),
.B(n_690),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_926),
.B(n_774),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_840),
.A2(n_689),
.B(n_675),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_918),
.B(n_690),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_969),
.B(n_689),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_811),
.A2(n_739),
.B1(n_702),
.B2(n_691),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_961),
.A2(n_430),
.B1(n_426),
.B2(n_405),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_L g1109 ( 
.A(n_874),
.B(n_691),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_893),
.A2(n_414),
.B(n_702),
.C(n_720),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_902),
.A2(n_701),
.B(n_696),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_968),
.A2(n_701),
.B(n_696),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_922),
.B(n_739),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_890),
.A2(n_720),
.B(n_730),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_964),
.B(n_775),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_927),
.B(n_895),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_924),
.B(n_739),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_811),
.A2(n_739),
.B1(n_629),
.B2(n_644),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_868),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_878),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_967),
.A2(n_792),
.B(n_731),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_878),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_883),
.A2(n_629),
.B(n_644),
.C(n_532),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_867),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_938),
.B(n_739),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_897),
.A2(n_792),
.B(n_731),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_944),
.B(n_739),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_801),
.B(n_730),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_963),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_906),
.A2(n_750),
.B(n_733),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_907),
.A2(n_750),
.B(n_733),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_885),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_885),
.B(n_764),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_804),
.B(n_764),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_811),
.A2(n_387),
.B1(n_389),
.B2(n_390),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_807),
.B(n_766),
.Y(n_1136)
);

CKINVDCx6p67_ASAP7_75t_R g1137 ( 
.A(n_928),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_942),
.A2(n_392),
.B1(n_393),
.B2(n_396),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_899),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_912),
.A2(n_773),
.B(n_766),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_810),
.B(n_773),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_820),
.B(n_780),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_913),
.A2(n_921),
.B(n_919),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_SL g1144 ( 
.A(n_896),
.B(n_356),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_899),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_931),
.A2(n_782),
.B(n_780),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_928),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_911),
.Y(n_1148)
);

AO21x2_ASAP7_75t_L g1149 ( 
.A1(n_803),
.A2(n_786),
.B(n_782),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_846),
.B(n_786),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_894),
.B(n_806),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_848),
.B(n_789),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_945),
.A2(n_790),
.B(n_789),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_842),
.B(n_401),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_853),
.B(n_790),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_911),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_916),
.B(n_923),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_916),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_939),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_811),
.B(n_798),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_880),
.Y(n_1161)
);

OAI321xp33_ASAP7_75t_L g1162 ( 
.A1(n_930),
.A2(n_551),
.A3(n_529),
.B1(n_530),
.B2(n_532),
.C(n_533),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_948),
.A2(n_958),
.B(n_952),
.Y(n_1163)
);

OAI21xp33_ASAP7_75t_L g1164 ( 
.A1(n_955),
.A2(n_303),
.B(n_302),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1027),
.A2(n_803),
.B(n_860),
.C(n_930),
.Y(n_1165)
);

INVx5_ASAP7_75t_L g1166 ( 
.A(n_1046),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1084),
.A2(n_860),
.B(n_930),
.C(n_923),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1030),
.B(n_914),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1030),
.B(n_966),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_983),
.A2(n_823),
.B(n_880),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_988),
.A2(n_823),
.B(n_880),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_1072),
.B(n_925),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1012),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1070),
.B(n_932),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1074),
.A2(n_932),
.B(n_821),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1008),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_976),
.A2(n_1000),
.B(n_996),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1008),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1046),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1039),
.A2(n_959),
.B(n_808),
.C(n_821),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_982),
.B(n_808),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1069),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1025),
.B(n_401),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1004),
.B(n_965),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1046),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1023),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_982),
.B(n_987),
.C(n_1091),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1001),
.A2(n_970),
.B(n_834),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1124),
.B(n_533),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_980),
.A2(n_421),
.B1(n_418),
.B2(n_413),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1059),
.A2(n_940),
.B(n_892),
.C(n_886),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_981),
.A2(n_834),
.B(n_830),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1129),
.B(n_644),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_984),
.A2(n_844),
.B(n_830),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1101),
.B(n_644),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1046),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_985),
.A2(n_852),
.B(n_844),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1061),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_L g1199 ( 
.A(n_1061),
.B(n_852),
.Y(n_1199)
);

OAI21xp33_ASAP7_75t_SL g1200 ( 
.A1(n_975),
.A2(n_892),
.B(n_886),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_977),
.A2(n_940),
.B1(n_409),
.B2(n_798),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1101),
.B(n_644),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1086),
.B(n_615),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1024),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1012),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1038),
.Y(n_1206)
);

NOR2x1_ASAP7_75t_L g1207 ( 
.A(n_1045),
.B(n_540),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_989),
.A2(n_568),
.B(n_570),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1017),
.A2(n_551),
.B(n_574),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1038),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1159),
.B(n_306),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1057),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_L g1213 ( 
.A1(n_979),
.A2(n_581),
.B(n_574),
.C(n_577),
.Y(n_1213)
);

AND2x6_ASAP7_75t_L g1214 ( 
.A(n_1061),
.B(n_615),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1061),
.Y(n_1215)
);

INVxp33_ASAP7_75t_L g1216 ( 
.A(n_1047),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1058),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1021),
.B(n_615),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1124),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1065),
.Y(n_1220)
);

BUFx8_ASAP7_75t_SL g1221 ( 
.A(n_1147),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_987),
.A2(n_574),
.B(n_614),
.C(n_612),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1009),
.A2(n_568),
.B(n_570),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1091),
.A2(n_641),
.B(n_638),
.C(n_636),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_993),
.B(n_356),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_993),
.B(n_1116),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1021),
.B(n_1053),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1011),
.A2(n_568),
.B(n_570),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1087),
.B(n_309),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1077),
.B(n_615),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1083),
.A2(n_1003),
.B(n_1029),
.C(n_998),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1161),
.B(n_577),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1045),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1077),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1122),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1083),
.A2(n_641),
.B(n_638),
.C(n_636),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_SL g1237 ( 
.A(n_1144),
.B(n_313),
.C(n_312),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1122),
.B(n_621),
.Y(n_1238)
);

CKINVDCx14_ASAP7_75t_R g1239 ( 
.A(n_1137),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1161),
.B(n_577),
.Y(n_1240)
);

NOR2x1_ASAP7_75t_L g1241 ( 
.A(n_1071),
.B(n_578),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1132),
.Y(n_1242)
);

BUFx2_ASAP7_75t_SL g1243 ( 
.A(n_1050),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_SL g1244 ( 
.A(n_986),
.B(n_356),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1132),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_995),
.A2(n_570),
.B(n_571),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1151),
.A2(n_356),
.B1(n_569),
.B2(n_567),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1058),
.B(n_570),
.Y(n_1248)
);

AOI22x1_ASAP7_75t_L g1249 ( 
.A1(n_1143),
.A2(n_641),
.B1(n_638),
.B2(n_636),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1080),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1156),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_990),
.A2(n_567),
.B(n_571),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1156),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_994),
.A2(n_567),
.B(n_571),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_974),
.A2(n_566),
.B(n_569),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1056),
.A2(n_566),
.B(n_569),
.Y(n_1256)
);

AO32x1_ASAP7_75t_L g1257 ( 
.A1(n_1108),
.A2(n_614),
.A3(n_580),
.B1(n_578),
.B2(n_612),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1104),
.A2(n_555),
.B(n_557),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1073),
.B(n_314),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1003),
.A2(n_641),
.B(n_638),
.C(n_636),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_991),
.A2(n_566),
.B(n_561),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1064),
.A2(n_557),
.B(n_561),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1073),
.A2(n_395),
.B1(n_328),
.B2(n_330),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1058),
.B(n_578),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1005),
.A2(n_580),
.B(n_581),
.C(n_612),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1154),
.B(n_323),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1058),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1080),
.A2(n_613),
.B1(n_580),
.B2(n_614),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1080),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1007),
.B(n_621),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1019),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1081),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1035),
.A2(n_557),
.B(n_561),
.Y(n_1273)
);

NOR3xp33_ASAP7_75t_L g1274 ( 
.A(n_1164),
.B(n_333),
.C(n_334),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1017),
.A2(n_406),
.B1(n_339),
.B2(n_343),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1042),
.A2(n_561),
.B(n_562),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1043),
.A2(n_562),
.B(n_555),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1063),
.A2(n_562),
.B(n_555),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1041),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1092),
.B(n_337),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1006),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1048),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1022),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1006),
.B(n_401),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1018),
.A2(n_1020),
.B(n_999),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1049),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1033),
.B(n_621),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1157),
.A2(n_562),
.B(n_603),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1037),
.A2(n_633),
.B(n_626),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1092),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1099),
.B(n_401),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1031),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1028),
.B(n_581),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1052),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1028),
.B(n_434),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1068),
.B(n_621),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1054),
.A2(n_633),
.B(n_626),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1118),
.A2(n_403),
.B1(n_353),
.B2(n_357),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_978),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1162),
.B(n_626),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_978),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1081),
.B(n_626),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1099),
.A2(n_415),
.B(n_359),
.C(n_362),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_R g1304 ( 
.A(n_1093),
.B(n_344),
.Y(n_1304)
);

CKINVDCx14_ASAP7_75t_R g1305 ( 
.A(n_1138),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1051),
.A2(n_633),
.B(n_603),
.C(n_595),
.Y(n_1306)
);

CKINVDCx14_ASAP7_75t_R g1307 ( 
.A(n_1135),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1106),
.A2(n_613),
.B1(n_434),
.B2(n_633),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1078),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1095),
.B(n_364),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1118),
.B(n_373),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1139),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1119),
.A2(n_1120),
.B1(n_1145),
.B2(n_1158),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1060),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1148),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1128),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1106),
.B(n_588),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1016),
.B(n_588),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1014),
.A2(n_590),
.B(n_603),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1026),
.B(n_590),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1060),
.Y(n_1321)
);

NOR3xp33_ASAP7_75t_L g1322 ( 
.A(n_1062),
.B(n_375),
.C(n_378),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1157),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1032),
.B(n_590),
.Y(n_1324)
);

OAI21xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1163),
.A2(n_590),
.B(n_595),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1010),
.A2(n_595),
.B(n_603),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1013),
.A2(n_595),
.B(n_611),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1177),
.A2(n_997),
.B(n_1015),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1285),
.A2(n_1123),
.A3(n_1051),
.B(n_1111),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1271),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1200),
.A2(n_1131),
.B(n_1130),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1177),
.A2(n_1112),
.B(n_1160),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1175),
.A2(n_1044),
.B(n_1088),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1188),
.A2(n_1146),
.B(n_1153),
.Y(n_1334)
);

NAND2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1172),
.B(n_1016),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1183),
.B(n_434),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1173),
.Y(n_1337)
);

NOR2x1_ASAP7_75t_L g1338 ( 
.A(n_1226),
.B(n_1040),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1175),
.A2(n_1089),
.B(n_1082),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1285),
.A2(n_1036),
.B(n_1090),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1171),
.A2(n_1002),
.B(n_1149),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1187),
.A2(n_1123),
.B(n_992),
.C(n_1100),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1291),
.B(n_434),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1288),
.A2(n_1075),
.B(n_1034),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_1229),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1168),
.B(n_1134),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_1211),
.Y(n_1348)
);

AO32x2_ASAP7_75t_L g1349 ( 
.A1(n_1313),
.A2(n_1110),
.A3(n_1149),
.B1(n_1094),
.B2(n_1114),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1178),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1258),
.A2(n_1126),
.B(n_1140),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1262),
.A2(n_1097),
.B(n_1121),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1213),
.A2(n_1155),
.B(n_1152),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1171),
.A2(n_1085),
.B(n_1103),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1176),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1255),
.A2(n_1150),
.B(n_1142),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1221),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1255),
.A2(n_1141),
.B(n_1136),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1182),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1327),
.A2(n_1133),
.B(n_1127),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1290),
.B(n_1055),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1170),
.A2(n_1103),
.B(n_1085),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1188),
.A2(n_1133),
.B(n_1067),
.Y(n_1363)
);

INVx3_ASAP7_75t_SL g1364 ( 
.A(n_1233),
.Y(n_1364)
);

AOI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1266),
.A2(n_381),
.B1(n_386),
.B2(n_388),
.C(n_397),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1280),
.B(n_1115),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1170),
.A2(n_1066),
.B(n_1076),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1217),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1279),
.B(n_398),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1186),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1203),
.A2(n_1125),
.B(n_1117),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1269),
.B(n_1109),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1246),
.A2(n_1107),
.B(n_1102),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1214),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1216),
.B(n_419),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1243),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1204),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1189),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1286),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1192),
.A2(n_1113),
.B(n_1079),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1259),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1246),
.A2(n_1105),
.B(n_1098),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1169),
.A2(n_1181),
.B1(n_1227),
.B2(n_1307),
.Y(n_1383)
);

NAND3x1_ASAP7_75t_L g1384 ( 
.A(n_1241),
.B(n_8),
.C(n_9),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1316),
.B(n_1096),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1206),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1327),
.A2(n_1110),
.B(n_431),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1165),
.A2(n_422),
.B(n_427),
.C(n_428),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1210),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1184),
.B(n_607),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1217),
.Y(n_1391)
);

NAND2x2_ASAP7_75t_L g1392 ( 
.A(n_1281),
.B(n_9),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1174),
.B(n_607),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1244),
.B(n_1284),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1315),
.B(n_1292),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1305),
.A2(n_607),
.B1(n_611),
.B2(n_16),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1326),
.A2(n_1289),
.A3(n_1256),
.B(n_1223),
.Y(n_1397)
);

BUFx2_ASAP7_75t_R g1398 ( 
.A(n_1267),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1212),
.B(n_607),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1278),
.A2(n_613),
.B(n_96),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1282),
.B(n_607),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1310),
.B(n_13),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1219),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1278),
.A2(n_613),
.B(n_100),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1166),
.B(n_607),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1303),
.A2(n_1225),
.B(n_1167),
.C(n_1237),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1220),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1219),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1326),
.A2(n_613),
.A3(n_611),
.B(n_607),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1234),
.B(n_611),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1245),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1231),
.A2(n_607),
.B1(n_611),
.B2(n_16),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1322),
.A2(n_613),
.B1(n_611),
.B2(n_17),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1235),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1180),
.A2(n_611),
.B(n_15),
.C(n_18),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1274),
.A2(n_13),
.B(n_20),
.C(n_21),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1194),
.A2(n_611),
.B(n_114),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_L g1418 ( 
.A(n_1272),
.B(n_613),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1166),
.B(n_112),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1197),
.A2(n_107),
.B(n_221),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1289),
.A2(n_1256),
.B(n_1319),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1320),
.A2(n_95),
.B(n_219),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1219),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1242),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1295),
.A2(n_613),
.B1(n_22),
.B2(n_23),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1250),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1250),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1250),
.B(n_115),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1273),
.A2(n_613),
.B(n_121),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1166),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1273),
.A2(n_613),
.B(n_217),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1276),
.A2(n_613),
.B(n_216),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_1239),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1223),
.A2(n_215),
.B(n_212),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1207),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1191),
.A2(n_24),
.B(n_32),
.C(n_33),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1304),
.B(n_35),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1193),
.B(n_35),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1325),
.A2(n_209),
.B(n_208),
.Y(n_1439)
);

INVx3_ASAP7_75t_SL g1440 ( 
.A(n_1272),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_R g1441 ( 
.A(n_1272),
.B(n_207),
.Y(n_1441)
);

INVx8_ASAP7_75t_L g1442 ( 
.A(n_1166),
.Y(n_1442)
);

CKINVDCx16_ASAP7_75t_R g1443 ( 
.A(n_1263),
.Y(n_1443)
);

O2A1O1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1298),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1251),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1253),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1276),
.A2(n_200),
.B(n_177),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1283),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1275),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1277),
.A2(n_169),
.B(n_164),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

O2A1O1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1311),
.A2(n_46),
.B(n_48),
.C(n_50),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1190),
.B(n_50),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1294),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1309),
.B(n_54),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1195),
.A2(n_160),
.B(n_158),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_SL g1457 ( 
.A1(n_1218),
.A2(n_155),
.B(n_150),
.C(n_147),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1314),
.B(n_1247),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1323),
.Y(n_1459)
);

AO32x2_ASAP7_75t_L g1460 ( 
.A1(n_1201),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1277),
.A2(n_140),
.B(n_130),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1249),
.A2(n_128),
.B(n_127),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1261),
.A2(n_123),
.B(n_59),
.Y(n_1463)
);

AO22x2_ASAP7_75t_L g1464 ( 
.A1(n_1300),
.A2(n_73),
.B1(n_60),
.B2(n_63),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1202),
.A2(n_55),
.B(n_64),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1299),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1324),
.A2(n_67),
.B(n_71),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1312),
.B(n_71),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1199),
.A2(n_73),
.B(n_1208),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1301),
.B(n_1240),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1261),
.A2(n_1265),
.B(n_1317),
.C(n_1252),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1270),
.Y(n_1472)
);

AOI221x1_ASAP7_75t_L g1473 ( 
.A1(n_1319),
.A2(n_1228),
.B1(n_1252),
.B2(n_1254),
.C(n_1222),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_SL g1474 ( 
.A(n_1232),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_SL g1475 ( 
.A(n_1321),
.B(n_1240),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1287),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1254),
.A2(n_1228),
.B(n_1230),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1238),
.A2(n_1302),
.B(n_1296),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_SL g1479 ( 
.A(n_1214),
.B(n_1248),
.Y(n_1479)
);

AO32x2_ASAP7_75t_L g1480 ( 
.A1(n_1257),
.A2(n_1209),
.A3(n_1260),
.B1(n_1224),
.B2(n_1236),
.Y(n_1480)
);

AO31x2_ASAP7_75t_L g1481 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1306),
.B(n_1214),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1297),
.A2(n_1293),
.B(n_1264),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1257),
.A2(n_1248),
.B(n_1318),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1179),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1318),
.A2(n_1179),
.B(n_1185),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1214),
.A2(n_1308),
.A3(n_1268),
.B(n_1198),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1185),
.A2(n_1196),
.B(n_1198),
.Y(n_1487)
);

AO31x2_ASAP7_75t_L g1488 ( 
.A1(n_1214),
.A2(n_1196),
.A3(n_1215),
.B(n_979),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1215),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1280),
.B(n_1027),
.C(n_1030),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1288),
.A2(n_1258),
.B(n_1262),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1200),
.A2(n_1084),
.B(n_1027),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1176),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1183),
.B(n_1070),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1183),
.B(n_1070),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1221),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1490),
.A2(n_1402),
.B1(n_1453),
.B2(n_1492),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1443),
.A2(n_1381),
.B1(n_1396),
.B2(n_1347),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1490),
.A2(n_1435),
.B1(n_1364),
.B2(n_1383),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1330),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1492),
.A2(n_1396),
.B1(n_1412),
.B2(n_1394),
.Y(n_1501)
);

INVx5_ASAP7_75t_L g1502 ( 
.A(n_1442),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1359),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1383),
.A2(n_1395),
.B1(n_1366),
.B2(n_1379),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1355),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1445),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1412),
.A2(n_1464),
.B1(n_1435),
.B2(n_1463),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1494),
.B(n_1495),
.Y(n_1508)
);

INVx6_ASAP7_75t_L g1509 ( 
.A(n_1442),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_R g1510 ( 
.A1(n_1379),
.A2(n_1359),
.B1(n_1376),
.B2(n_1365),
.Y(n_1510)
);

CKINVDCx6p67_ASAP7_75t_R g1511 ( 
.A(n_1433),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1425),
.A2(n_1413),
.B(n_1437),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1442),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1464),
.A2(n_1463),
.B1(n_1413),
.B2(n_1425),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1350),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1348),
.A2(n_1467),
.B1(n_1439),
.B2(n_1344),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1348),
.A2(n_1439),
.B1(n_1392),
.B2(n_1346),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1370),
.Y(n_1518)
);

INVx6_ASAP7_75t_L g1519 ( 
.A(n_1423),
.Y(n_1519)
);

BUFx10_ASAP7_75t_L g1520 ( 
.A(n_1496),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1430),
.Y(n_1521)
);

BUFx12f_ASAP7_75t_L g1522 ( 
.A(n_1423),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1346),
.A2(n_1438),
.B1(n_1338),
.B2(n_1336),
.Y(n_1523)
);

CKINVDCx6p67_ASAP7_75t_R g1524 ( 
.A(n_1440),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1430),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1475),
.A2(n_1460),
.B1(n_1474),
.B2(n_1479),
.Y(n_1526)
);

BUFx2_ASAP7_75t_SL g1527 ( 
.A(n_1474),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1361),
.B(n_1378),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1403),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1475),
.A2(n_1460),
.B1(n_1479),
.B2(n_1419),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1423),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1458),
.A2(n_1339),
.B1(n_1337),
.B2(n_1388),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1375),
.A2(n_1335),
.B1(n_1369),
.B2(n_1372),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1372),
.A2(n_1469),
.B1(n_1468),
.B2(n_1455),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1470),
.A2(n_1476),
.B1(n_1472),
.B2(n_1466),
.Y(n_1535)
);

INVx6_ASAP7_75t_L g1536 ( 
.A(n_1430),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1426),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1385),
.A2(n_1398),
.B1(n_1374),
.B2(n_1406),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1428),
.A2(n_1384),
.B1(n_1436),
.B2(n_1408),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1428),
.A2(n_1418),
.B1(n_1427),
.B2(n_1454),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1448),
.A2(n_1415),
.B1(n_1401),
.B2(n_1451),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1451),
.A2(n_1426),
.B1(n_1414),
.B2(n_1424),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1426),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1459),
.A2(n_1377),
.B1(n_1386),
.B2(n_1389),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1407),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1411),
.B(n_1446),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1460),
.A2(n_1419),
.B1(n_1374),
.B2(n_1434),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1489),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1493),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1449),
.A2(n_1444),
.B1(n_1416),
.B2(n_1420),
.Y(n_1550)
);

BUFx4_ASAP7_75t_R g1551 ( 
.A(n_1441),
.Y(n_1551)
);

INVx6_ASAP7_75t_L g1552 ( 
.A(n_1484),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1484),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1399),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1484),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1399),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1487),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1410),
.Y(n_1558)
);

BUFx8_ASAP7_75t_L g1559 ( 
.A(n_1480),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1488),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1374),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1465),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1434),
.A2(n_1373),
.B1(n_1422),
.B2(n_1331),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1373),
.A2(n_1331),
.B1(n_1382),
.B2(n_1390),
.Y(n_1564)
);

AO22x1_ASAP7_75t_L g1565 ( 
.A1(n_1368),
.A2(n_1391),
.B1(n_1393),
.B2(n_1363),
.Y(n_1565)
);

CKINVDCx11_ASAP7_75t_R g1566 ( 
.A(n_1456),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1452),
.B(n_1485),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1405),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1368),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1343),
.A2(n_1471),
.B1(n_1482),
.B2(n_1417),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1447),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1410),
.Y(n_1572)
);

INVx6_ASAP7_75t_L g1573 ( 
.A(n_1354),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1360),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1360),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1342),
.A2(n_1462),
.B1(n_1450),
.B2(n_1461),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1387),
.A2(n_1353),
.B1(n_1363),
.B2(n_1382),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1387),
.A2(n_1334),
.B1(n_1483),
.B2(n_1421),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1353),
.A2(n_1421),
.B1(n_1358),
.B2(n_1356),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1362),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_1356),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1397),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1334),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1358),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1371),
.A2(n_1478),
.B1(n_1367),
.B2(n_1380),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1328),
.A2(n_1340),
.B1(n_1333),
.B2(n_1341),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1486),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1332),
.A2(n_1477),
.B1(n_1431),
.B2(n_1429),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1486),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1457),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1486),
.Y(n_1591)
);

INVx3_ASAP7_75t_SL g1592 ( 
.A(n_1480),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1473),
.A2(n_1349),
.B1(n_1480),
.B2(n_1329),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1397),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1409),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1397),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1329),
.B(n_1409),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1400),
.A2(n_1404),
.B1(n_1432),
.B2(n_1352),
.Y(n_1598)
);

INVx4_ASAP7_75t_L g1599 ( 
.A(n_1409),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1345),
.A2(n_1351),
.B1(n_1491),
.B2(n_1349),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1481),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1481),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1470),
.B(n_1403),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1402),
.A2(n_1084),
.B1(n_1030),
.B2(n_1027),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1490),
.A2(n_982),
.B1(n_1030),
.B2(n_1168),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1412),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1355),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1364),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1442),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1364),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1402),
.A2(n_1030),
.B1(n_640),
.B2(n_1266),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1347),
.B(n_1030),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1442),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1330),
.Y(n_1614)
);

BUFx2_ASAP7_75t_SL g1615 ( 
.A(n_1474),
.Y(n_1615)
);

CKINVDCx11_ASAP7_75t_R g1616 ( 
.A(n_1433),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1357),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1618)
);

INVx5_ASAP7_75t_L g1619 ( 
.A(n_1442),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1490),
.A2(n_982),
.B1(n_1030),
.B2(n_1168),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1402),
.A2(n_582),
.B1(n_1244),
.B2(n_1030),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1490),
.A2(n_982),
.B1(n_1030),
.B2(n_1168),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1623)
);

CKINVDCx6p67_ASAP7_75t_R g1624 ( 
.A(n_1364),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1402),
.A2(n_582),
.B1(n_1244),
.B2(n_1030),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1402),
.A2(n_1030),
.B1(n_640),
.B2(n_1266),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1330),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1330),
.Y(n_1631)
);

BUFx4f_ASAP7_75t_SL g1632 ( 
.A(n_1364),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1364),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_SL g1634 ( 
.A(n_1346),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1635)
);

INVx8_ASAP7_75t_L g1636 ( 
.A(n_1442),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1364),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1347),
.B(n_1030),
.Y(n_1638)
);

INVx4_ASAP7_75t_L g1639 ( 
.A(n_1442),
.Y(n_1639)
);

CKINVDCx11_ASAP7_75t_R g1640 ( 
.A(n_1433),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1355),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1490),
.A2(n_982),
.B1(n_1030),
.B2(n_1168),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1435),
.A2(n_1490),
.B1(n_1027),
.B2(n_1425),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1494),
.B(n_1495),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1359),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1355),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1364),
.Y(n_1648)
);

CKINVDCx11_ASAP7_75t_R g1649 ( 
.A(n_1433),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1330),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1488),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1402),
.A2(n_1084),
.B1(n_1030),
.B2(n_1027),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1402),
.A2(n_582),
.B1(n_1244),
.B2(n_1030),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1359),
.B(n_1395),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1402),
.A2(n_1084),
.B1(n_1030),
.B2(n_1027),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1355),
.Y(n_1657)
);

INVx6_ASAP7_75t_L g1658 ( 
.A(n_1442),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1402),
.A2(n_582),
.B1(n_1244),
.B2(n_1030),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1364),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1490),
.A2(n_1027),
.B1(n_1030),
.B2(n_1402),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1330),
.Y(n_1662)
);

CKINVDCx11_ASAP7_75t_R g1663 ( 
.A(n_1433),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1402),
.A2(n_582),
.B1(n_1244),
.B2(n_1030),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1357),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1490),
.A2(n_982),
.B1(n_1030),
.B2(n_1168),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1402),
.A2(n_582),
.B1(n_1244),
.B2(n_1030),
.Y(n_1667)
);

CKINVDCx6p67_ASAP7_75t_R g1668 ( 
.A(n_1364),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1582),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1596),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1574),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1575),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1515),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1587),
.B(n_1583),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1580),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1651),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1560),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1518),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1591),
.B(n_1597),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1509),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1502),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1573),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1654),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1557),
.B(n_1589),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1586),
.A2(n_1588),
.B(n_1579),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1612),
.B(n_1638),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1594),
.B(n_1504),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1500),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1509),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1589),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1497),
.A2(n_1626),
.B1(n_1653),
.B2(n_1621),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1581),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1522),
.Y(n_1694)
);

INVx5_ASAP7_75t_L g1695 ( 
.A(n_1573),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1621),
.A2(n_1653),
.B1(n_1626),
.B2(n_1664),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1526),
.B(n_1530),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1531),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1503),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1526),
.B(n_1530),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1497),
.A2(n_1667),
.B1(n_1659),
.B2(n_1664),
.Y(n_1701)
);

CKINVDCx14_ASAP7_75t_R g1702 ( 
.A(n_1616),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1548),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1602),
.B(n_1564),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1581),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1592),
.B(n_1564),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1614),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1584),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1579),
.A2(n_1600),
.B(n_1585),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1630),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1601),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1573),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1601),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1631),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1592),
.B(n_1507),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1650),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1598),
.A2(n_1563),
.B(n_1567),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1561),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1606),
.A2(n_1538),
.B(n_1561),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1662),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1645),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1577),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1506),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1545),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1563),
.A2(n_1572),
.B(n_1558),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1549),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1507),
.B(n_1547),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1604),
.B(n_1652),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1528),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1554),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1501),
.B(n_1546),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1553),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1559),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1556),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1640),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1505),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1555),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1656),
.A2(n_1643),
.B1(n_1655),
.B2(n_1623),
.C(n_1618),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1593),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1593),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1514),
.B(n_1644),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1565),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1514),
.B(n_1607),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1559),
.Y(n_1745)
);

NAND2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1502),
.B(n_1619),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1544),
.A2(n_1516),
.B(n_1541),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1659),
.A2(n_1667),
.B1(n_1499),
.B2(n_1618),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1544),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1569),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1623),
.B(n_1625),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1641),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1646),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1657),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1595),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1599),
.Y(n_1756)
);

AOI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1605),
.A2(n_1642),
.B(n_1666),
.Y(n_1757)
);

AO21x2_ASAP7_75t_L g1758 ( 
.A1(n_1643),
.A2(n_1606),
.B(n_1622),
.Y(n_1758)
);

BUFx2_ASAP7_75t_R g1759 ( 
.A(n_1665),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_R g1760 ( 
.A(n_1649),
.B(n_1663),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1542),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1509),
.Y(n_1762)
);

AO21x1_ASAP7_75t_L g1763 ( 
.A1(n_1550),
.A2(n_1620),
.B(n_1512),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1578),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1578),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1516),
.A2(n_1534),
.B(n_1532),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1576),
.Y(n_1767)
);

INVx4_ASAP7_75t_L g1768 ( 
.A(n_1502),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1625),
.B(n_1647),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1561),
.Y(n_1770)
);

AND2x2_ASAP7_75t_SL g1771 ( 
.A(n_1627),
.B(n_1629),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1576),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1590),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1611),
.A2(n_1628),
.B(n_1627),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1629),
.B(n_1647),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1498),
.B(n_1661),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1540),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1635),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1635),
.B(n_1661),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1508),
.B(n_1523),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1655),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1502),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1539),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1523),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1533),
.A2(n_1517),
.B(n_1562),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1535),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1517),
.B(n_1603),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1619),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1603),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1608),
.B(n_1610),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_SL g1791 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1510),
.A2(n_1634),
.B1(n_1632),
.B2(n_1624),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1529),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1521),
.B(n_1525),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1619),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1552),
.Y(n_1796)
);

AOI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1566),
.A2(n_1536),
.B(n_1519),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1636),
.A2(n_1609),
.B(n_1658),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_SL g1799 ( 
.A(n_1633),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1637),
.A2(n_1648),
.B(n_1660),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1609),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1543),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1527),
.B(n_1615),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1513),
.A2(n_1613),
.B(n_1639),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1668),
.B(n_1632),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1658),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1519),
.B(n_1639),
.Y(n_1807)
);

AO21x1_ASAP7_75t_SL g1808 ( 
.A1(n_1551),
.A2(n_1636),
.B(n_1634),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1675),
.B(n_1742),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1675),
.B(n_1511),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1696),
.A2(n_1617),
.B1(n_1524),
.B2(n_1537),
.C(n_1520),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1731),
.B(n_1519),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1684),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1742),
.B(n_1789),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1676),
.B(n_1687),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1674),
.B(n_1679),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1669),
.B(n_1766),
.Y(n_1817)
);

AOI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1797),
.A2(n_1769),
.B(n_1751),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1739),
.A2(n_1763),
.B1(n_1701),
.B2(n_1692),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1771),
.A2(n_1763),
.B1(n_1748),
.B2(n_1774),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1730),
.Y(n_1821)
);

OA21x2_ASAP7_75t_L g1822 ( 
.A1(n_1717),
.A2(n_1686),
.B(n_1767),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1775),
.A2(n_1779),
.B1(n_1729),
.B2(n_1778),
.C(n_1781),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1680),
.B(n_1744),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1771),
.A2(n_1792),
.B1(n_1727),
.B2(n_1728),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1674),
.B(n_1679),
.Y(n_1826)
);

BUFx4f_ASAP7_75t_SL g1827 ( 
.A(n_1703),
.Y(n_1827)
);

OR2x6_ASAP7_75t_L g1828 ( 
.A(n_1669),
.B(n_1766),
.Y(n_1828)
);

AO32x1_ASAP7_75t_L g1829 ( 
.A1(n_1727),
.A2(n_1728),
.A3(n_1700),
.B1(n_1697),
.B2(n_1776),
.Y(n_1829)
);

AO21x2_ASAP7_75t_L g1830 ( 
.A1(n_1757),
.A2(n_1686),
.B(n_1717),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1724),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1757),
.A2(n_1771),
.B(n_1747),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1731),
.B(n_1735),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1732),
.B(n_1676),
.Y(n_1834)
);

NAND2x1p5_ASAP7_75t_L g1835 ( 
.A(n_1695),
.B(n_1798),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1693),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1779),
.A2(n_1778),
.B1(n_1781),
.B2(n_1776),
.C(n_1758),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1735),
.B(n_1758),
.Y(n_1838)
);

OA21x2_ASAP7_75t_L g1839 ( 
.A1(n_1767),
.A2(n_1772),
.B(n_1747),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1733),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1719),
.A2(n_1783),
.B(n_1785),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1719),
.A2(n_1783),
.B(n_1669),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_L g1843 ( 
.A(n_1676),
.B(n_1790),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1724),
.Y(n_1844)
);

AO32x2_ASAP7_75t_L g1845 ( 
.A1(n_1740),
.A2(n_1741),
.A3(n_1690),
.B1(n_1762),
.B2(n_1801),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1743),
.A2(n_1792),
.B(n_1777),
.Y(n_1846)
);

OAI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1777),
.A2(n_1784),
.B(n_1725),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_SL g1848 ( 
.A1(n_1697),
.A2(n_1700),
.B1(n_1758),
.B2(n_1715),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1749),
.B(n_1708),
.Y(n_1849)
);

AO32x1_ASAP7_75t_L g1850 ( 
.A1(n_1772),
.A2(n_1722),
.A3(n_1715),
.B1(n_1713),
.B2(n_1711),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1734),
.B(n_1745),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1693),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1773),
.A2(n_1745),
.B1(n_1786),
.B2(n_1780),
.Y(n_1853)
);

INVx4_ASAP7_75t_L g1854 ( 
.A(n_1718),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1750),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1749),
.B(n_1708),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1726),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1726),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1798),
.A2(n_1725),
.B(n_1683),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1706),
.B(n_1787),
.Y(n_1860)
);

AO32x2_ASAP7_75t_L g1861 ( 
.A1(n_1681),
.A2(n_1762),
.A3(n_1801),
.B1(n_1768),
.B2(n_1682),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1688),
.B(n_1704),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1800),
.B(n_1695),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1706),
.B(n_1787),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1784),
.B(n_1689),
.Y(n_1865)
);

AOI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1786),
.A2(n_1722),
.B(n_1765),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1723),
.B(n_1720),
.Y(n_1867)
);

CKINVDCx6p67_ASAP7_75t_R g1868 ( 
.A(n_1733),
.Y(n_1868)
);

CKINVDCx11_ASAP7_75t_R g1869 ( 
.A(n_1703),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1761),
.A2(n_1765),
.B(n_1764),
.Y(n_1870)
);

NOR2x1_ASAP7_75t_R g1871 ( 
.A(n_1736),
.B(n_1738),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1707),
.Y(n_1872)
);

O2A1O1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1773),
.A2(n_1721),
.B(n_1699),
.C(n_1764),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1710),
.B(n_1714),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1714),
.B(n_1716),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1736),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1695),
.A2(n_1803),
.B(n_1683),
.C(n_1712),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1670),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1746),
.B(n_1797),
.Y(n_1879)
);

OAI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1702),
.A2(n_1803),
.B(n_1793),
.C(n_1805),
.Y(n_1880)
);

OAI21x1_ASAP7_75t_L g1881 ( 
.A1(n_1683),
.A2(n_1712),
.B(n_1755),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1671),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1683),
.A2(n_1712),
.B1(n_1793),
.B2(n_1808),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1738),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1759),
.Y(n_1885)
);

OA21x2_ASAP7_75t_L g1886 ( 
.A1(n_1705),
.A2(n_1671),
.B(n_1756),
.Y(n_1886)
);

AO32x2_ASAP7_75t_L g1887 ( 
.A1(n_1681),
.A2(n_1682),
.A3(n_1768),
.B1(n_1677),
.B2(n_1691),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1794),
.B(n_1802),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1799),
.B(n_1760),
.Y(n_1889)
);

OAI211xp5_ASAP7_75t_L g1890 ( 
.A1(n_1804),
.A2(n_1754),
.B(n_1753),
.C(n_1709),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1823),
.B(n_1806),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1836),
.Y(n_1892)
);

NAND2xp33_ASAP7_75t_R g1893 ( 
.A(n_1885),
.B(n_1807),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1836),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1815),
.B(n_1760),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1821),
.B(n_1813),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1820),
.A2(n_1712),
.B1(n_1808),
.B2(n_1695),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1809),
.B(n_1834),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1852),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1852),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1819),
.A2(n_1695),
.B1(n_1806),
.B2(n_1770),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1860),
.B(n_1691),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1878),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1816),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1841),
.A2(n_1695),
.B1(n_1791),
.B2(n_1782),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1864),
.B(n_1672),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1826),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1859),
.B(n_1685),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1824),
.B(n_1705),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1841),
.A2(n_1791),
.B1(n_1782),
.B2(n_1682),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1862),
.B(n_1709),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1825),
.A2(n_1807),
.B1(n_1788),
.B2(n_1795),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1839),
.B(n_1709),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1839),
.B(n_1709),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1881),
.B(n_1685),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1826),
.B(n_1685),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1855),
.Y(n_1917)
);

NAND3xp33_ASAP7_75t_L g1918 ( 
.A(n_1823),
.B(n_1754),
.C(n_1788),
.Y(n_1918)
);

AND2x2_ASAP7_75t_SL g1919 ( 
.A(n_1837),
.B(n_1782),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1861),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1886),
.Y(n_1921)
);

INVxp67_ASAP7_75t_SL g1922 ( 
.A(n_1838),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1886),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1814),
.B(n_1752),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1838),
.B(n_1673),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1865),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1874),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1817),
.B(n_1828),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1843),
.B(n_1752),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1867),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1875),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1817),
.B(n_1755),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1849),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1861),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1867),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1848),
.B(n_1756),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1861),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1848),
.B(n_1678),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1882),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1882),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1833),
.Y(n_1941)
);

NOR2x1_ASAP7_75t_R g1942 ( 
.A(n_1891),
.B(n_1869),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1927),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1929),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1921),
.Y(n_1945)
);

NAND2x1_ASAP7_75t_L g1946 ( 
.A(n_1928),
.B(n_1879),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1911),
.B(n_1822),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1911),
.B(n_1822),
.Y(n_1948)
);

NAND3xp33_ASAP7_75t_L g1949 ( 
.A(n_1918),
.B(n_1837),
.C(n_1811),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1917),
.B(n_1870),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1896),
.B(n_1847),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1920),
.B(n_1887),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1892),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1934),
.B(n_1887),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1892),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1894),
.Y(n_1956)
);

OAI33xp33_ASAP7_75t_L g1957 ( 
.A1(n_1939),
.A2(n_1825),
.A3(n_1853),
.B1(n_1873),
.B2(n_1849),
.B3(n_1856),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1894),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1899),
.Y(n_1959)
);

NAND3xp33_ASAP7_75t_SL g1960 ( 
.A(n_1910),
.B(n_1811),
.C(n_1880),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1934),
.A2(n_1873),
.B1(n_1866),
.B2(n_1832),
.C(n_1846),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1921),
.Y(n_1962)
);

INVx4_ASAP7_75t_L g1963 ( 
.A(n_1919),
.Y(n_1963)
);

OAI33xp33_ASAP7_75t_L g1964 ( 
.A1(n_1939),
.A2(n_1853),
.A3(n_1856),
.B1(n_1812),
.B2(n_1833),
.B3(n_1872),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1933),
.B(n_1870),
.Y(n_1965)
);

AO21x2_ASAP7_75t_L g1966 ( 
.A1(n_1923),
.A2(n_1832),
.B(n_1830),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_SL g1967 ( 
.A1(n_1919),
.A2(n_1842),
.B1(n_1880),
.B2(n_1828),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1937),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1915),
.Y(n_1969)
);

NAND3xp33_ASAP7_75t_L g1970 ( 
.A(n_1919),
.B(n_1846),
.C(n_1866),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1900),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1903),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1928),
.B(n_1879),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1927),
.B(n_1847),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1931),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1906),
.B(n_1851),
.Y(n_1976)
);

OAI33xp33_ASAP7_75t_L g1977 ( 
.A1(n_1940),
.A2(n_1812),
.A3(n_1872),
.B1(n_1863),
.B2(n_1796),
.B3(n_1844),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1916),
.B(n_1845),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1916),
.B(n_1845),
.Y(n_1979)
);

AOI221xp5_ASAP7_75t_L g1980 ( 
.A1(n_1922),
.A2(n_1936),
.B1(n_1914),
.B2(n_1913),
.C(n_1938),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1916),
.B(n_1845),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1915),
.Y(n_1982)
);

INVxp67_ASAP7_75t_SL g1983 ( 
.A(n_1925),
.Y(n_1983)
);

OAI321xp33_ASAP7_75t_L g1984 ( 
.A1(n_1912),
.A2(n_1842),
.A3(n_1818),
.B1(n_1890),
.B2(n_1877),
.C(n_1835),
.Y(n_1984)
);

AO21x2_ASAP7_75t_L g1985 ( 
.A1(n_1913),
.A2(n_1914),
.B(n_1890),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1902),
.B(n_1888),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1903),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1940),
.Y(n_1988)
);

OAI322xp33_ASAP7_75t_L g1989 ( 
.A1(n_1930),
.A2(n_1889),
.A3(n_1829),
.B1(n_1858),
.B2(n_1857),
.C1(n_1831),
.C2(n_1737),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1932),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1972),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1972),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1967),
.B(n_1963),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1978),
.B(n_1928),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1987),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1978),
.B(n_1936),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1968),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1979),
.B(n_1909),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1983),
.B(n_1930),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1987),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1953),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1944),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1988),
.B(n_1951),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1979),
.B(n_1909),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1981),
.B(n_1926),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1953),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1955),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1974),
.B(n_1925),
.Y(n_2008)
);

INVx4_ASAP7_75t_L g2009 ( 
.A(n_1963),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1955),
.Y(n_2010)
);

NAND2x1_ASAP7_75t_L g2011 ( 
.A(n_1963),
.B(n_1915),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1965),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1945),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1963),
.B(n_1904),
.Y(n_2014)
);

INVx4_ASAP7_75t_L g2015 ( 
.A(n_1990),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1944),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1984),
.A2(n_1829),
.B(n_1850),
.Y(n_2017)
);

INVx4_ASAP7_75t_L g2018 ( 
.A(n_1990),
.Y(n_2018)
);

NAND2xp33_ASAP7_75t_SL g2019 ( 
.A(n_1942),
.B(n_1893),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1988),
.B(n_1935),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1949),
.B(n_1905),
.Y(n_2021)
);

NOR2x1_ASAP7_75t_L g2022 ( 
.A(n_1949),
.B(n_1895),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1973),
.B(n_1908),
.Y(n_2023)
);

INVxp67_ASAP7_75t_SL g2024 ( 
.A(n_1945),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1974),
.B(n_1898),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1968),
.B(n_1907),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_1956),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1951),
.B(n_1935),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1973),
.B(n_1908),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1962),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1944),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1956),
.B(n_1941),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1958),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1952),
.B(n_1954),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1947),
.B(n_1924),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2001),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2013),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1994),
.B(n_2034),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1994),
.B(n_1952),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2012),
.B(n_1950),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2001),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2006),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2012),
.B(n_1980),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_2019),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2006),
.Y(n_2045)
);

AOI33xp33_ASAP7_75t_L g2046 ( 
.A1(n_2002),
.A2(n_1961),
.A3(n_1954),
.B1(n_1938),
.B2(n_1971),
.B3(n_1959),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2034),
.B(n_1969),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2013),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2007),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2013),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2007),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1997),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1996),
.B(n_1969),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2010),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2022),
.B(n_1876),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2010),
.Y(n_2056)
);

XNOR2x1_ASAP7_75t_L g2057 ( 
.A(n_2022),
.B(n_1810),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_2030),
.Y(n_2058)
);

AOI32xp33_ASAP7_75t_L g2059 ( 
.A1(n_2021),
.A2(n_1942),
.A3(n_1960),
.B1(n_1970),
.B2(n_1957),
.Y(n_2059)
);

INVxp67_ASAP7_75t_SL g2060 ( 
.A(n_1997),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1996),
.B(n_1969),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2002),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2023),
.B(n_1969),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2028),
.B(n_2003),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_2030),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2028),
.B(n_1976),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2023),
.B(n_1982),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2033),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2033),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_2009),
.B(n_1973),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2027),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2027),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_2003),
.B(n_1947),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2032),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2023),
.B(n_1982),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2032),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_2008),
.B(n_1948),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2025),
.B(n_1976),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2020),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2020),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1991),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2023),
.B(n_1982),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2008),
.B(n_1948),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2025),
.B(n_1986),
.Y(n_2084)
);

AND3x2_ASAP7_75t_L g2085 ( 
.A(n_2014),
.B(n_1943),
.C(n_1975),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1991),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_2055),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2059),
.B(n_2031),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_2038),
.B(n_2009),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2038),
.B(n_2015),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2064),
.B(n_1999),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_2070),
.B(n_2009),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2036),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2064),
.B(n_1999),
.Y(n_2094)
);

AND2x4_ASAP7_75t_SL g2095 ( 
.A(n_2062),
.B(n_2009),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2084),
.B(n_1993),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2036),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2078),
.B(n_2035),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2039),
.B(n_2015),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2060),
.B(n_2040),
.Y(n_2100)
);

INVxp67_ASAP7_75t_L g2101 ( 
.A(n_2057),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2059),
.B(n_2046),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2041),
.Y(n_2103)
);

NOR2x1_ASAP7_75t_L g2104 ( 
.A(n_2044),
.B(n_2016),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2041),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2047),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2057),
.B(n_2031),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2039),
.B(n_2015),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2042),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2066),
.B(n_2035),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2070),
.B(n_2015),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2043),
.B(n_2017),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_2070),
.B(n_1827),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2042),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_2070),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2052),
.B(n_1985),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2045),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2071),
.B(n_2017),
.Y(n_2118)
);

INVx1_ASAP7_75t_SL g2119 ( 
.A(n_2085),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2063),
.B(n_2018),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2073),
.B(n_1985),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_2053),
.Y(n_2122)
);

AND2x2_ASAP7_75t_SL g2123 ( 
.A(n_2071),
.B(n_1884),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2047),
.Y(n_2124)
);

CKINVDCx16_ASAP7_75t_R g2125 ( 
.A(n_2053),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2061),
.Y(n_2126)
);

NAND3xp33_ASAP7_75t_SL g2127 ( 
.A(n_2102),
.B(n_1970),
.C(n_2011),
.Y(n_2127)
);

AOI322xp5_ASAP7_75t_L g2128 ( 
.A1(n_2101),
.A2(n_2088),
.A3(n_2112),
.B1(n_2107),
.B2(n_2119),
.C1(n_2118),
.C2(n_2104),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2093),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2100),
.B(n_2073),
.Y(n_2130)
);

O2A1O1Ixp33_ASAP7_75t_SL g2131 ( 
.A1(n_2116),
.A2(n_2072),
.B(n_2011),
.C(n_1871),
.Y(n_2131)
);

OAI321xp33_ASAP7_75t_L g2132 ( 
.A1(n_2100),
.A2(n_2072),
.A3(n_2065),
.B1(n_2058),
.B2(n_2076),
.C(n_2080),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_2095),
.Y(n_2133)
);

AOI211xp5_ASAP7_75t_L g2134 ( 
.A1(n_2113),
.A2(n_1989),
.B(n_1964),
.C(n_2074),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2096),
.B(n_2077),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2091),
.B(n_2077),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2099),
.Y(n_2137)
);

OAI21xp33_ASAP7_75t_L g2138 ( 
.A1(n_2115),
.A2(n_2076),
.B(n_2074),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_2087),
.B(n_2113),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2097),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_SL g2141 ( 
.A(n_2116),
.B(n_1884),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_SL g2142 ( 
.A1(n_2087),
.A2(n_2016),
.B1(n_1985),
.B2(n_2061),
.Y(n_2142)
);

AOI322xp5_ASAP7_75t_L g2143 ( 
.A1(n_2123),
.A2(n_2005),
.A3(n_2024),
.B1(n_2079),
.B2(n_2080),
.C1(n_1998),
.C2(n_2004),
.Y(n_2143)
);

OAI221xp5_ASAP7_75t_SL g2144 ( 
.A1(n_2121),
.A2(n_2083),
.B1(n_1897),
.B2(n_1901),
.C(n_2016),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2099),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2095),
.B(n_2079),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2123),
.A2(n_1829),
.B(n_1946),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_2125),
.B(n_1868),
.Y(n_2148)
);

OAI31xp33_ASAP7_75t_L g2149 ( 
.A1(n_2089),
.A2(n_2082),
.A3(n_2075),
.B(n_2067),
.Y(n_2149)
);

AOI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_2092),
.A2(n_1946),
.B(n_1989),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2122),
.B(n_2005),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2103),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2105),
.Y(n_2153)
);

AOI211xp5_ASAP7_75t_SL g2154 ( 
.A1(n_2092),
.A2(n_2063),
.B(n_2082),
.C(n_2075),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2109),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2155),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_2139),
.B(n_2092),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2133),
.B(n_2089),
.Y(n_2158)
);

OAI21xp5_ASAP7_75t_SL g2159 ( 
.A1(n_2127),
.A2(n_2089),
.B(n_2090),
.Y(n_2159)
);

INVxp67_ASAP7_75t_L g2160 ( 
.A(n_2139),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2142),
.A2(n_2124),
.B1(n_2106),
.B2(n_2098),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2129),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_2130),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2140),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_2148),
.A2(n_2090),
.B1(n_2111),
.B2(n_2108),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_2137),
.B(n_2145),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_2136),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2152),
.Y(n_2168)
);

OAI21xp33_ASAP7_75t_L g2169 ( 
.A1(n_2128),
.A2(n_2143),
.B(n_2138),
.Y(n_2169)
);

NAND2xp33_ASAP7_75t_L g2170 ( 
.A(n_2135),
.B(n_2111),
.Y(n_2170)
);

O2A1O1Ixp33_ASAP7_75t_SL g2171 ( 
.A1(n_2148),
.A2(n_2121),
.B(n_2094),
.C(n_2091),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2146),
.B(n_2106),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2153),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2132),
.A2(n_2094),
.B(n_2114),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_2144),
.B(n_2151),
.Y(n_2175)
);

A2O1A1Ixp33_ASAP7_75t_L g2176 ( 
.A1(n_2147),
.A2(n_2108),
.B(n_2124),
.C(n_2126),
.Y(n_2176)
);

AOI322xp5_ASAP7_75t_L g2177 ( 
.A1(n_2142),
.A2(n_2126),
.A3(n_2117),
.B1(n_2120),
.B2(n_2065),
.C1(n_2058),
.C2(n_2024),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2154),
.B(n_2120),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2141),
.Y(n_2179)
);

BUFx2_ASAP7_75t_L g2180 ( 
.A(n_2141),
.Y(n_2180)
);

AOI21x1_ASAP7_75t_L g2181 ( 
.A1(n_2180),
.A2(n_2163),
.B(n_2161),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2167),
.B(n_2098),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2167),
.B(n_2110),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2178),
.B(n_2149),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2163),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2166),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2160),
.B(n_2110),
.Y(n_2187)
);

NAND3x1_ASAP7_75t_L g2188 ( 
.A(n_2157),
.B(n_2150),
.C(n_2131),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2160),
.B(n_2134),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_2171),
.A2(n_2131),
.B(n_2065),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2169),
.A2(n_2018),
.B1(n_1884),
.B2(n_1840),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_2157),
.B(n_2018),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2166),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2156),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2186),
.B(n_2175),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2191),
.A2(n_2175),
.B1(n_2174),
.B2(n_2170),
.Y(n_2196)
);

NAND3xp33_ASAP7_75t_SL g2197 ( 
.A(n_2190),
.B(n_2159),
.C(n_2177),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_2191),
.B(n_2179),
.C(n_2172),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_2187),
.B(n_2165),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2185),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2193),
.B(n_2158),
.Y(n_2201)
);

O2A1O1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2189),
.A2(n_2173),
.B(n_2168),
.C(n_2162),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2182),
.Y(n_2203)
);

O2A1O1Ixp33_ASAP7_75t_L g2204 ( 
.A1(n_2192),
.A2(n_2164),
.B(n_2176),
.C(n_2058),
.Y(n_2204)
);

AOI211xp5_ASAP7_75t_SL g2205 ( 
.A1(n_2184),
.A2(n_2067),
.B(n_2083),
.C(n_2049),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2183),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2203),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_L g2208 ( 
.A(n_2195),
.B(n_2181),
.C(n_2194),
.Y(n_2208)
);

AOI21xp33_ASAP7_75t_SL g2209 ( 
.A1(n_2206),
.A2(n_2188),
.B(n_2049),
.Y(n_2209)
);

NOR2x1_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_1694),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2196),
.A2(n_2018),
.B1(n_2068),
.B2(n_2045),
.Y(n_2211)
);

O2A1O1Ixp5_ASAP7_75t_SL g2212 ( 
.A1(n_2200),
.A2(n_2054),
.B(n_2051),
.C(n_2056),
.Y(n_2212)
);

O2A1O1Ixp33_ASAP7_75t_L g2213 ( 
.A1(n_2202),
.A2(n_1694),
.B(n_1698),
.C(n_2050),
.Y(n_2213)
);

AO211x2_ASAP7_75t_L g2214 ( 
.A1(n_2208),
.A2(n_2198),
.B(n_2201),
.C(n_2205),
.Y(n_2214)
);

AOI211xp5_ASAP7_75t_L g2215 ( 
.A1(n_2209),
.A2(n_2199),
.B(n_2204),
.C(n_2196),
.Y(n_2215)
);

AOI211xp5_ASAP7_75t_L g2216 ( 
.A1(n_2211),
.A2(n_1698),
.B(n_2051),
.C(n_2068),
.Y(n_2216)
);

AOI211xp5_ASAP7_75t_SL g2217 ( 
.A1(n_2207),
.A2(n_2069),
.B(n_2056),
.C(n_2054),
.Y(n_2217)
);

NAND2x1_ASAP7_75t_SL g2218 ( 
.A(n_2210),
.B(n_2069),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2213),
.A2(n_2081),
.B1(n_2037),
.B2(n_2050),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2212),
.A2(n_2048),
.B(n_2050),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2219),
.B(n_2037),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2218),
.Y(n_2222)
);

NOR3xp33_ASAP7_75t_L g2223 ( 
.A(n_2215),
.B(n_2048),
.C(n_2081),
.Y(n_2223)
);

XOR2xp5_ASAP7_75t_L g2224 ( 
.A(n_2214),
.B(n_1883),
.Y(n_2224)
);

NAND4xp75_ASAP7_75t_L g2225 ( 
.A(n_2220),
.B(n_2048),
.C(n_2086),
.D(n_2014),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2222),
.B(n_2216),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_2224),
.A2(n_2086),
.B1(n_2217),
.B2(n_2029),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_2223),
.A2(n_2086),
.B1(n_1966),
.B2(n_1977),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_2226),
.Y(n_2229)
);

CKINVDCx20_ASAP7_75t_R g2230 ( 
.A(n_2229),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2230),
.A2(n_2227),
.B1(n_2221),
.B2(n_2228),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_2230),
.A2(n_2225),
.B(n_2029),
.Y(n_2232)
);

NAND2x1p5_ASAP7_75t_L g2233 ( 
.A(n_2232),
.B(n_1718),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2231),
.Y(n_2234)
);

OA22x2_ASAP7_75t_L g2235 ( 
.A1(n_2234),
.A2(n_2029),
.B1(n_1992),
.B2(n_1995),
.Y(n_2235)
);

OAI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_2233),
.A2(n_2029),
.B(n_2026),
.Y(n_2236)
);

INVx1_ASAP7_75t_SL g2237 ( 
.A(n_2235),
.Y(n_2237)
);

OAI222xp33_ASAP7_75t_SL g2238 ( 
.A1(n_2237),
.A2(n_2236),
.B1(n_1682),
.B2(n_1768),
.C1(n_1854),
.C2(n_2000),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_2238),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2239),
.A2(n_1966),
.B1(n_1992),
.B2(n_2000),
.Y(n_2240)
);

AOI211xp5_ASAP7_75t_L g2241 ( 
.A1(n_2240),
.A2(n_1718),
.B(n_1782),
.C(n_1795),
.Y(n_2241)
);


endmodule