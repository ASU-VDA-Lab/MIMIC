module fake_jpeg_9880_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_22),
.B1(n_34),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_22),
.B1(n_42),
.B2(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_60),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_45),
.B(n_48),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_83),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_38),
.B1(n_47),
.B2(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_62),
.B1(n_22),
.B2(n_18),
.Y(n_126)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_79),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_91),
.B1(n_101),
.B2(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_80),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_87),
.Y(n_120)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_94),
.C(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_26),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_41),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_27),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_28),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_39),
.C(n_46),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_32),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_28),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_28),
.Y(n_116)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_74),
.B1(n_70),
.B2(n_77),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_122),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_42),
.B1(n_47),
.B2(n_22),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_104),
.B1(n_108),
.B2(n_69),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_131),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_99),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_128),
.B1(n_100),
.B2(n_70),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_83),
.A2(n_18),
.B1(n_34),
.B2(n_43),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_137),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_142),
.B1(n_152),
.B2(n_157),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_82),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_30),
.C(n_29),
.Y(n_178)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_139),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_78),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_100),
.B1(n_88),
.B2(n_98),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_82),
.B(n_100),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_153),
.B(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_145),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_72),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_151),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_116),
.B1(n_120),
.B2(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_162),
.B1(n_84),
.B2(n_33),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_161),
.B1(n_119),
.B2(n_125),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_18),
.B1(n_19),
.B2(n_102),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_104),
.A2(n_92),
.B1(n_69),
.B2(n_34),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_119),
.B1(n_106),
.B2(n_23),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_102),
.B1(n_50),
.B2(n_53),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_79),
.B1(n_28),
.B2(n_33),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_123),
.B1(n_53),
.B2(n_28),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_171),
.B1(n_194),
.B2(n_149),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_143),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_166),
.C(n_169),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_103),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_172),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_118),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_103),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_107),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_174),
.A2(n_188),
.B1(n_193),
.B2(n_13),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_24),
.B1(n_32),
.B2(n_14),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_30),
.C(n_16),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_178),
.C(n_181),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_2),
.B(n_3),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_137),
.B(n_35),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_30),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_147),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_186),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_144),
.B(n_17),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_23),
.B1(n_35),
.B2(n_25),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_13),
.B(n_12),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_25),
.B1(n_35),
.B2(n_17),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_192),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_30),
.B(n_32),
.C(n_16),
.D(n_12),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_24),
.B(n_14),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_85),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_149),
.B1(n_153),
.B2(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_2),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_132),
.B(n_32),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_202),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_215),
.B1(n_221),
.B2(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_213),
.Y(n_246)
);

AO21x2_ASAP7_75t_SL g205 ( 
.A1(n_164),
.A2(n_151),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_140),
.B1(n_138),
.B2(n_145),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_211),
.B1(n_216),
.B2(n_188),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_25),
.B1(n_24),
.B2(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_185),
.B(n_2),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_218),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_177),
.B(n_3),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_211),
.Y(n_245)
);

NOR2x1p5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_11),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_181),
.B1(n_178),
.B2(n_166),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_176),
.A2(n_4),
.B(n_5),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_11),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_165),
.C(n_189),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_232),
.C(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_184),
.C(n_168),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_200),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_214),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_169),
.C(n_197),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_163),
.C(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_217),
.C(n_202),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_170),
.B1(n_5),
.B2(n_6),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_12),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_224),
.C(n_227),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_198),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_253),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_11),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_261),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_204),
.C(n_213),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_265),
.C(n_268),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_199),
.C(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_270),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_219),
.C(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_246),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_243),
.B(n_205),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_223),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_201),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_205),
.C(n_222),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_248),
.B1(n_252),
.B2(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_235),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_265),
.A2(n_252),
.B1(n_229),
.B2(n_205),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_288),
.B1(n_4),
.B2(n_5),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_249),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_228),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_286),
.Y(n_298)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_229),
.B1(n_238),
.B2(n_233),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_251),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_10),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_231),
.C(n_250),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_255),
.C(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_244),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_255),
.B(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_210),
.C(n_220),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_218),
.C(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_300),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_4),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_302),
.Y(n_315)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

AO21x2_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_4),
.B(n_5),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_306),
.B(n_6),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_6),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_304),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_6),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_277),
.B1(n_290),
.B2(n_288),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_309),
.B(n_318),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_311),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_287),
.B1(n_291),
.B2(n_285),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_298),
.B1(n_300),
.B2(n_294),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_287),
.B1(n_8),
.B2(n_9),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_306),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_320),
.B(n_296),
.Y(n_331)
);

INVx11_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_318),
.B(n_312),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_7),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_297),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_295),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_308),
.B(n_314),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_332),
.B(n_322),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_331),
.B(n_323),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_328),
.B(n_324),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_334),
.A2(n_335),
.B(n_336),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_329),
.B(n_321),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_323),
.B(n_313),
.C(n_9),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_7),
.B(n_8),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_9),
.Y(n_342)
);


endmodule