module fake_aes_12383_n_720 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_720);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_720;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_2), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_2), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_73), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_76), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_42), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_53), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_34), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_102), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_88), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_46), .Y(n_117) );
BUFx10_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_7), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_106), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_96), .Y(n_122) );
INVx2_ASAP7_75t_SL g123 ( .A(n_98), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_95), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_52), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_59), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_58), .Y(n_127) );
BUFx10_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_65), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_83), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_74), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_48), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_62), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_6), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_9), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_36), .Y(n_138) );
INVx1_ASAP7_75t_SL g139 ( .A(n_57), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_80), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_94), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_0), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_20), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_55), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_33), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_71), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_60), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_15), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_77), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_123), .B(n_0), .Y(n_153) );
AOI22x1_ASAP7_75t_L g154 ( .A1(n_123), .A2(n_40), .B1(n_104), .B2(n_103), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_149), .B(n_1), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_107), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_144), .B(n_3), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_115), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_136), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_107), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_118), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_115), .B(n_4), .Y(n_166) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_117), .A2(n_5), .B(n_6), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_120), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_125), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_156), .A2(n_142), .B1(n_150), .B2(n_109), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_165), .B(n_152), .Y(n_173) );
INVx8_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_165), .B(n_118), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_165), .B(n_109), .Y(n_177) );
INVx5_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_165), .B(n_128), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_165), .B(n_128), .Y(n_180) );
AND3x2_ASAP7_75t_L g181 ( .A(n_162), .B(n_151), .C(n_145), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_165), .B(n_126), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_155), .B(n_127), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_152), .B(n_129), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_152), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_152), .B(n_137), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_156), .A2(n_150), .B1(n_137), .B2(n_142), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_152), .B(n_108), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_153), .B(n_128), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_166), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_162), .B(n_108), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_164), .B(n_168), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_196), .B(n_155), .Y(n_197) );
AOI221xp5_ASAP7_75t_L g198 ( .A1(n_171), .A2(n_164), .B1(n_157), .B2(n_168), .C(n_169), .Y(n_198) );
O2A1O1Ixp5_ASAP7_75t_L g199 ( .A1(n_192), .A2(n_153), .B(n_166), .C(n_168), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_173), .A2(n_153), .B(n_166), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_177), .B(n_155), .Y(n_201) );
INVxp67_ASAP7_75t_L g202 ( .A(n_194), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_188), .B(n_169), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_186), .B(n_153), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_174), .Y(n_205) );
AND2x6_ASAP7_75t_SL g206 ( .A(n_183), .B(n_157), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_176), .B(n_169), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_191), .B(n_166), .Y(n_208) );
INVxp67_ASAP7_75t_L g209 ( .A(n_183), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_174), .A2(n_187), .B(n_193), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_187), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_174), .B(n_110), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_182), .B(n_170), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_179), .B(n_110), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_174), .B(n_186), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_172), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_193), .Y(n_217) );
NOR2x1p5_ASAP7_75t_L g218 ( .A(n_171), .B(n_119), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_183), .B(n_170), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_174), .A2(n_167), .B1(n_159), .B2(n_170), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_113), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_190), .A2(n_167), .B1(n_111), .B2(n_124), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_186), .B(n_113), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_183), .B(n_114), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_190), .A2(n_167), .B1(n_116), .B2(n_133), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_183), .B(n_114), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_185), .B(n_122), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_184), .A2(n_167), .B1(n_146), .B2(n_141), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_202), .B(n_185), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_198), .A2(n_167), .B1(n_178), .B2(n_175), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_209), .A2(n_178), .B1(n_135), .B2(n_141), .Y(n_233) );
NAND3xp33_ASAP7_75t_SL g234 ( .A(n_222), .B(n_225), .C(n_230), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_200), .A2(n_178), .B(n_189), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_230), .A2(n_178), .B1(n_122), .B2(n_135), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_205), .B(n_178), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_204), .A2(n_178), .B(n_195), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_218), .B(n_197), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_189), .B(n_163), .C(n_161), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_195), .B(n_167), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_218), .B(n_181), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_201), .B(n_163), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_208), .A2(n_154), .B(n_138), .Y(n_245) );
OR2x6_ASAP7_75t_SL g246 ( .A(n_224), .B(n_130), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_203), .B(n_158), .Y(n_247) );
AO22x1_ASAP7_75t_L g248 ( .A1(n_227), .A2(n_131), .B1(n_139), .B2(n_140), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_210), .A2(n_154), .B(n_134), .Y(n_249) );
NAND2xp33_ASAP7_75t_L g250 ( .A(n_220), .B(n_154), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_213), .A2(n_148), .B(n_147), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_199), .A2(n_143), .B(n_160), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_219), .B(n_158), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_132), .B(n_160), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_222), .A2(n_161), .B1(n_160), .B2(n_158), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_211), .A2(n_161), .B(n_8), .C(n_9), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_225), .A2(n_7), .B1(n_8), .B2(n_10), .Y(n_257) );
OA22x2_ASAP7_75t_L g258 ( .A1(n_206), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_217), .A2(n_45), .B(n_101), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_211), .A2(n_226), .B(n_223), .C(n_212), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_207), .A2(n_44), .B(n_100), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_257), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_249), .A2(n_226), .B(n_229), .Y(n_263) );
AOI21x1_ASAP7_75t_L g264 ( .A1(n_245), .A2(n_229), .B(n_216), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_239), .B(n_206), .Y(n_265) );
INVx5_ASAP7_75t_L g266 ( .A(n_241), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_241), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_237), .B(n_215), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_246), .Y(n_269) );
BUFx8_ASAP7_75t_L g270 ( .A(n_243), .Y(n_270) );
BUFx10_ASAP7_75t_L g271 ( .A(n_243), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_247), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_261), .A2(n_216), .B(n_228), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
OAI21xp5_ASAP7_75t_SL g276 ( .A1(n_234), .A2(n_221), .B(n_214), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_244), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g278 ( .A1(n_236), .A2(n_11), .B(n_12), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_242), .A2(n_47), .B(n_99), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_233), .Y(n_280) );
AO31x2_ASAP7_75t_L g281 ( .A1(n_256), .A2(n_13), .A3(n_14), .B(n_15), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_240), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_256), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_255), .B(n_13), .Y(n_284) );
BUFx12f_ASAP7_75t_L g285 ( .A(n_258), .Y(n_285) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_279), .A2(n_259), .B(n_254), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_283), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_279), .A2(n_258), .B(n_252), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_282), .A2(n_250), .B(n_232), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_275), .A2(n_232), .B1(n_231), .B2(n_251), .Y(n_291) );
AO31x2_ASAP7_75t_L g292 ( .A1(n_274), .A2(n_238), .A3(n_260), .B(n_248), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_272), .B(n_237), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_273), .A2(n_260), .B(n_50), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_282), .A2(n_14), .B(n_16), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_272), .B(n_16), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_273), .A2(n_51), .B(n_97), .Y(n_299) );
OAI21x1_ASAP7_75t_SL g300 ( .A1(n_276), .A2(n_17), .B(n_18), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_263), .A2(n_17), .B(n_18), .Y(n_301) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_274), .A2(n_54), .B(n_92), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_277), .B(n_19), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_19), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_263), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_275), .B(n_49), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_304), .B(n_265), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_296), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_304), .B(n_281), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_304), .B(n_285), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_305), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_305), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_281), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_298), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_288), .Y(n_319) );
CKINVDCx14_ASAP7_75t_R g320 ( .A(n_297), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_288), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_293), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_298), .B(n_281), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_297), .B(n_281), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_305), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_294), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_306), .B(n_285), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_297), .B(n_281), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_301), .Y(n_333) );
INVx5_ASAP7_75t_L g334 ( .A(n_331), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_320), .B(n_303), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_310), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_322), .B(n_303), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_322), .B(n_295), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_323), .B(n_301), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_312), .A2(n_262), .B1(n_280), .B2(n_269), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_307), .B(n_295), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_323), .B(n_290), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_307), .B(n_327), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_331), .B(n_296), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_311), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_327), .B(n_290), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_313), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_328), .B(n_302), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_328), .B(n_292), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_329), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_331), .B(n_296), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_319), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_332), .B(n_302), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_331), .B(n_296), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_300), .B1(n_278), .B2(n_284), .C(n_291), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_329), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_316), .B(n_292), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_321), .B(n_302), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_315), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_331), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_321), .B(n_302), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_316), .B(n_302), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_324), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_324), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_337), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_376), .B(n_325), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_376), .B(n_325), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_354), .B(n_309), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_353), .B(n_333), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_359), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_344), .B(n_333), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_369), .B(n_334), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_369), .B(n_317), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_345), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_353), .B(n_330), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_361), .B(n_326), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_334), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_342), .B(n_308), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_347), .B(n_308), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_347), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_348), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_348), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_349), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_361), .B(n_326), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_349), .B(n_326), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_350), .B(n_317), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_350), .B(n_317), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_355), .B(n_317), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_355), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_362), .B(n_300), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_362), .B(n_300), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_367), .B(n_370), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_334), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_334), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_340), .B(n_292), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_336), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_335), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_336), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_367), .B(n_302), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_370), .B(n_371), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_351), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_371), .B(n_289), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_375), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_334), .B(n_289), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_340), .B(n_292), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_354), .B(n_289), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_366), .B(n_289), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_338), .B(n_292), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_366), .B(n_292), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_351), .B(n_292), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_351), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_352), .B(n_292), .Y(n_434) );
AND2x4_ASAP7_75t_SL g435 ( .A(n_369), .B(n_271), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_352), .B(n_292), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_338), .B(n_291), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_343), .B(n_20), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_334), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_352), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_356), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_356), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_375), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_378), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_405), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_426), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_378), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_438), .B(n_341), .C(n_364), .D(n_369), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_421), .B(n_356), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_379), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_421), .B(n_365), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_414), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_380), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_380), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_390), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_439), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_390), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_413), .B(n_339), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_384), .B(n_358), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_396), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_413), .B(n_339), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_396), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_384), .B(n_365), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_385), .B(n_365), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_418), .B(n_341), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_386), .B(n_358), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_397), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_385), .B(n_358), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_431), .B(n_374), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_431), .B(n_374), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_397), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_429), .B(n_374), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_405), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_393), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_429), .B(n_372), .Y(n_478) );
AND2x4_ASAP7_75t_SL g479 ( .A(n_414), .B(n_357), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_381), .B(n_372), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_405), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_398), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_402), .B(n_372), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_398), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_399), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_399), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_406), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_402), .B(n_368), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_406), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_387), .B(n_343), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_439), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_414), .B(n_363), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_381), .B(n_368), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_403), .B(n_368), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_407), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_403), .B(n_377), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_391), .B(n_377), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_382), .B(n_363), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_408), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_382), .B(n_363), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_408), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_428), .B(n_363), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_392), .B(n_357), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_391), .B(n_377), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_411), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_383), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_423), .B(n_357), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_411), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_424), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_423), .B(n_357), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_412), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_428), .B(n_346), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_412), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_424), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_395), .Y(n_516) );
NAND2xp33_ASAP7_75t_L g517 ( .A(n_415), .B(n_306), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_394), .B(n_346), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_437), .B(n_346), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_392), .B(n_400), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_430), .B(n_21), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_416), .B(n_21), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_427), .B(n_22), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_404), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_401), .B(n_22), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_417), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_520), .Y(n_527) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_469), .B(n_388), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_468), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_507), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_449), .B(n_400), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_388), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_444), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_490), .B(n_433), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_450), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_508), .B(n_388), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_479), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_469), .B(n_388), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_469), .B(n_389), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_507), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_453), .B(n_389), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_449), .B(n_432), .Y(n_543) );
NOR2x1p5_ASAP7_75t_SL g544 ( .A(n_445), .B(n_443), .Y(n_544) );
NAND2x1_ASAP7_75t_SL g545 ( .A(n_493), .B(n_420), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_452), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_451), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_452), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_511), .B(n_389), .Y(n_549) );
NOR2xp33_ASAP7_75t_SL g550 ( .A(n_455), .B(n_435), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_511), .B(n_389), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_455), .Y(n_552) );
AND3x1_ASAP7_75t_L g553 ( .A(n_467), .B(n_420), .C(n_410), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_490), .B(n_433), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_460), .B(n_432), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_448), .A2(n_409), .B1(n_435), .B2(n_434), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_458), .A2(n_425), .A3(n_306), .B1(n_441), .B2(n_440), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_454), .Y(n_558) );
INVx3_ASAP7_75t_L g559 ( .A(n_479), .Y(n_559) );
OR2x6_ASAP7_75t_L g560 ( .A(n_493), .B(n_425), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_456), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_472), .B(n_425), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_463), .B(n_442), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_461), .B(n_442), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_472), .B(n_473), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_457), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_465), .B(n_441), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_473), .B(n_436), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_458), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_466), .B(n_436), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_493), .B(n_422), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_524), .B(n_422), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_466), .B(n_434), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_471), .B(n_440), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_480), .B(n_417), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_459), .Y(n_577) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_521), .A2(n_23), .B(n_24), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_446), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_492), .B(n_419), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_477), .B(n_443), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_462), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_471), .B(n_419), .Y(n_583) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_467), .A2(n_306), .B(n_24), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_526), .B(n_383), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_498), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_517), .A2(n_306), .B(n_299), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_516), .B(n_443), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_494), .B(n_424), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_464), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_470), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_474), .B(n_435), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_503), .B(n_23), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_475), .B(n_299), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_294), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_505), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_475), .B(n_299), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_482), .B(n_294), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_484), .B(n_294), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_478), .B(n_299), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_522), .A2(n_268), .B1(n_267), .B2(n_270), .C(n_266), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_478), .B(n_286), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_286), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_528), .A2(n_513), .B(n_499), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_559), .B(n_501), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_580), .Y(n_607) );
OAI322xp33_ASAP7_75t_L g608 ( .A1(n_593), .A2(n_554), .A3(n_535), .B1(n_556), .B2(n_555), .C1(n_527), .C2(n_563), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_535), .B(n_497), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_588), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_559), .B(n_497), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_579), .B(n_523), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_554), .B(n_483), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g614 ( .A(n_601), .B(n_525), .C(n_519), .D(n_518), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_553), .A2(n_483), .B1(n_488), .B2(n_495), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_539), .A2(n_538), .B1(n_572), .B2(n_542), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_550), .A2(n_517), .B(n_515), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_563), .B(n_488), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_588), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_580), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_584), .A2(n_506), .B(n_514), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_540), .B(n_489), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_579), .B(n_491), .Y(n_623) );
OAI32xp33_ASAP7_75t_L g624 ( .A1(n_539), .A2(n_485), .A3(n_487), .B1(n_486), .B2(n_496), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_532), .B(n_495), .Y(n_625) );
INVxp33_ASAP7_75t_L g626 ( .A(n_550), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_529), .B(n_500), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_573), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_601), .A2(n_502), .B1(n_512), .B2(n_509), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_603), .A2(n_515), .B1(n_510), .B2(n_481), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_573), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_562), .A2(n_510), .B1(n_481), .B2(n_476), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_578), .A2(n_476), .B(n_445), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_578), .A2(n_286), .B(n_268), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_537), .B(n_270), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_549), .B(n_551), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_571), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_586), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g639 ( .A1(n_572), .A2(n_268), .A3(n_267), .B(n_270), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_542), .A2(n_266), .B1(n_267), .B2(n_270), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_586), .B(n_286), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_565), .B(n_286), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_533), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_534), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_545), .A2(n_267), .B(n_266), .C(n_271), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_546), .B(n_286), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_560), .A2(n_266), .B1(n_264), .B2(n_271), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_530), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_568), .B(n_264), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_570), .B(n_266), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_543), .B(n_25), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_536), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_547), .A2(n_271), .B1(n_27), .B2(n_28), .C(n_29), .Y(n_653) );
OAI21xp33_ASAP7_75t_L g654 ( .A1(n_626), .A2(n_575), .B(n_544), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_605), .A2(n_540), .B1(n_602), .B2(n_560), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_628), .B(n_574), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_615), .A2(n_548), .A3(n_596), .B1(n_575), .B2(n_583), .C1(n_590), .C2(n_582), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_616), .A2(n_560), .B1(n_531), .B2(n_552), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_612), .A2(n_592), .B1(n_569), .B2(n_561), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_616), .A2(n_621), .B1(n_624), .B2(n_635), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_614), .A2(n_592), .B1(n_594), .B2(n_600), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_611), .B(n_583), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_631), .B(n_558), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_610), .Y(n_664) );
INVxp33_ASAP7_75t_L g665 ( .A(n_639), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_629), .A2(n_566), .B1(n_577), .B2(n_591), .Y(n_666) );
AOI211x1_ASAP7_75t_L g667 ( .A1(n_621), .A2(n_557), .B(n_587), .C(n_585), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_608), .A2(n_541), .B1(n_581), .B2(n_597), .C(n_585), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_604), .A2(n_581), .B1(n_587), .B2(n_599), .C1(n_598), .C2(n_595), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_619), .B(n_576), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_640), .A2(n_567), .B(n_564), .C(n_589), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_617), .B(n_645), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_633), .A2(n_599), .B1(n_598), .B2(n_31), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_606), .A2(n_627), .B1(n_622), .B2(n_623), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_637), .B(n_26), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_643), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_644), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_611), .A2(n_30), .B1(n_35), .B2(n_37), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_633), .A2(n_38), .B1(n_39), .B2(n_41), .C(n_43), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_634), .A2(n_56), .B(n_61), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_652), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_657), .B(n_630), .Y(n_682) );
CKINVDCx16_ASAP7_75t_R g683 ( .A(n_658), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_660), .B(n_634), .C(n_640), .D(n_653), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_665), .B(n_622), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_667), .A2(n_638), .B1(n_642), .B2(n_641), .C(n_613), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_672), .A2(n_650), .B(n_647), .Y(n_687) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_668), .A2(n_646), .B1(n_648), .B2(n_606), .C1(n_609), .C2(n_607), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_660), .B(n_651), .C(n_620), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_655), .A2(n_618), .B1(n_632), .B2(n_636), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_661), .A2(n_649), .B1(n_625), .B2(n_66), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_671), .B(n_63), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_663), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_654), .A2(n_64), .B(n_67), .C(n_68), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_659), .B(n_674), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_684), .B(n_679), .C(n_678), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_683), .B(n_673), .C(n_675), .Y(n_697) );
NOR3xp33_ASAP7_75t_SL g698 ( .A(n_685), .B(n_673), .C(n_680), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_689), .A2(n_669), .B1(n_666), .B2(n_664), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_694), .B(n_681), .C(n_677), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_692), .B(n_662), .Y(n_701) );
NAND4xp25_ASAP7_75t_SL g702 ( .A(n_688), .B(n_656), .C(n_670), .D(n_676), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_696), .B(n_682), .C(n_695), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_699), .B(n_693), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_701), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_697), .B(n_687), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_691), .B(n_690), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_705), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_704), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_708), .Y(n_710) );
XOR2x1_ASAP7_75t_L g711 ( .A(n_709), .B(n_703), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_710), .A2(n_707), .B1(n_698), .B2(n_686), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_711), .A2(n_702), .B(n_700), .Y(n_713) );
OAI31xp33_ASAP7_75t_SL g714 ( .A1(n_713), .A2(n_69), .A3(n_70), .B(n_72), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_712), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_75), .B(n_79), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_716), .B(n_714), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g718 ( .A1(n_717), .A2(n_81), .B(n_82), .Y(n_718) );
OR2x6_ASAP7_75t_L g719 ( .A(n_718), .B(n_85), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_86), .B1(n_90), .B2(n_105), .Y(n_720) );
endmodule