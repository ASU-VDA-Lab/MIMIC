module fake_jpeg_16233_n_355 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_31),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_67),
.Y(n_84)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_61),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_31),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_0),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_36),
.B1(n_34),
.B2(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_24),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_22),
.B1(n_19),
.B2(n_45),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_88),
.A2(n_92),
.B1(n_69),
.B2(n_60),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_49),
.B1(n_55),
.B2(n_69),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_45),
.B1(n_24),
.B2(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_23),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_110),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_55),
.B1(n_70),
.B2(n_49),
.Y(n_127)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_42),
.B1(n_51),
.B2(n_38),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_68),
.A3(n_48),
.B1(n_51),
.B2(n_38),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_109),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_77),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_32),
.Y(n_109)
);

CKINVDCx9p33_ASAP7_75t_R g111 ( 
.A(n_54),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_67),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_63),
.B1(n_70),
.B2(n_58),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_114),
.B1(n_97),
.B2(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_102),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_127),
.B1(n_137),
.B2(n_139),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_23),
.B(n_0),
.Y(n_120)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_125),
.CON(n_155),
.SN(n_155)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_32),
.C(n_23),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_80),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_23),
.B(n_0),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_142),
.B1(n_94),
.B2(n_56),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_127),
.B1(n_119),
.B2(n_121),
.Y(n_178)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_152),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_132),
.Y(n_185)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_162),
.Y(n_169)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_102),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_94),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_115),
.B(n_104),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_130),
.B(n_128),
.Y(n_192)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_126),
.B(n_139),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_172),
.B(n_182),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_131),
.B(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_188),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_118),
.B1(n_123),
.B2(n_119),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_185),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_162),
.B1(n_160),
.B2(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_147),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_143),
.A3(n_155),
.B1(n_144),
.B2(n_145),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_136),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_186),
.C(n_194),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_85),
.C(n_50),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_117),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_193),
.B(n_98),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_158),
.A2(n_105),
.B(n_23),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_147),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_18),
.B(n_85),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_52),
.C(n_50),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_199),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_150),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_0),
.B(n_61),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_212),
.Y(n_230)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_200),
.B(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_165),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_202),
.C(n_210),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_164),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_148),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_52),
.C(n_101),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_157),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_192),
.B1(n_193),
.B2(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_148),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_216),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_159),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_101),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_153),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_178),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_51),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_185),
.B1(n_194),
.B2(n_181),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_223),
.A2(n_229),
.B1(n_38),
.B2(n_27),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_226),
.A2(n_235),
.B1(n_247),
.B2(n_48),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_153),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_209),
.A2(n_152),
.B1(n_134),
.B2(n_124),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_246),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_152),
.B1(n_98),
.B2(n_124),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_95),
.Y(n_239)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_198),
.B(n_95),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_202),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_245),
.B(n_196),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_56),
.B1(n_75),
.B2(n_134),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_25),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_201),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_210),
.B1(n_213),
.B2(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_250),
.B(n_267),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_211),
.B1(n_215),
.B2(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_SL g257 ( 
.A(n_224),
.B(n_1),
.C(n_2),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

AOI21x1_ASAP7_75t_SL g259 ( 
.A1(n_234),
.A2(n_105),
.B(n_48),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_259),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_25),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_25),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_266),
.C(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_37),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_1),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_231),
.B1(n_237),
.B2(n_238),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_37),
.Y(n_302)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_232),
.C(n_231),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_287),
.C(n_289),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_243),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_232),
.C(n_222),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_244),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_254),
.B(n_256),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_301),
.C(n_302),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_258),
.B(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_263),
.B1(n_264),
.B2(n_260),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_297),
.A2(n_289),
.B1(n_288),
.B2(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_245),
.Y(n_300)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_266),
.C(n_27),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_275),
.B1(n_279),
.B2(n_40),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_3),
.B(n_4),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_276),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_L g305 ( 
.A1(n_273),
.A2(n_37),
.A3(n_28),
.B1(n_20),
.B2(n_9),
.C(n_10),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_286),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_273),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_311),
.C(n_317),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_314),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_279),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_318),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_316),
.A2(n_28),
.B1(n_20),
.B2(n_10),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_28),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_5),
.Y(n_318)
);

OR2x4_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_5),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_6),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_5),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_6),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_292),
.Y(n_321)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_323),
.B(n_326),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_324),
.B(n_330),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_297),
.CI(n_302),
.CON(n_327),
.SN(n_327)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_331),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_329),
.B(n_8),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_294),
.B(n_296),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_6),
.Y(n_330)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_307),
.C(n_311),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_332),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_20),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_339),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_8),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_346),
.Y(n_349)
);

OAI221xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_328),
.B1(n_331),
.B2(n_12),
.C(n_13),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_9),
.Y(n_344)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_344),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_9),
.Y(n_346)
);

AOI322xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_342),
.A3(n_337),
.B1(n_345),
.B2(n_334),
.C1(n_11),
.C2(n_15),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

OAI221xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_347),
.B1(n_348),
.B2(n_17),
.C(n_12),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_12),
.C(n_13),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_17),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);


endmodule