module fake_jpeg_12976_n_399 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_399);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_399;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_29),
.C(n_26),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_52),
.Y(n_90)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_25),
.A2(n_1),
.B(n_3),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_54),
.B(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_66),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx12f_ASAP7_75t_SL g67 ( 
.A(n_36),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_83),
.Y(n_101)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_5),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_70),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_37),
.B(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_36),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_28),
.B1(n_30),
.B2(n_40),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_42),
.B1(n_38),
.B2(n_21),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_89),
.B1(n_113),
.B2(n_51),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_43),
.B1(n_40),
.B2(n_30),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_87),
.A2(n_102),
.B1(n_120),
.B2(n_130),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_42),
.B1(n_38),
.B2(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_88),
.A2(n_123),
.B1(n_125),
.B2(n_11),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_38),
.B1(n_42),
.B2(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_28),
.B1(n_41),
.B2(n_31),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_104),
.B1(n_109),
.B2(n_118),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_43),
.B1(n_40),
.B2(n_30),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_56),
.B1(n_71),
.B2(n_45),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_48),
.A2(n_16),
.B1(n_41),
.B2(n_31),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_62),
.A2(n_84),
.B1(n_81),
.B2(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_49),
.A2(n_16),
.B1(n_18),
.B2(n_23),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_43),
.B1(n_39),
.B2(n_33),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_49),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_18),
.B1(n_55),
.B2(n_73),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_5),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_26),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_132),
.A2(n_139),
.B1(n_155),
.B2(n_158),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_74),
.B1(n_68),
.B2(n_77),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_154),
.B1(n_166),
.B2(n_100),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_77),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_138),
.Y(n_186)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_65),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_63),
.B1(n_46),
.B2(n_7),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_144),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_121),
.B(n_122),
.Y(n_141)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_92),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_58),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_SL g191 ( 
.A(n_142),
.B(n_116),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_65),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_6),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_157),
.Y(n_198)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_161),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_9),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_127),
.Y(n_160)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_11),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_168),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_86),
.B(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_161),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_170),
.A2(n_154),
.B1(n_146),
.B2(n_168),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_110),
.B(n_100),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_116),
.C(n_103),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_105),
.B1(n_103),
.B2(n_114),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_108),
.B1(n_105),
.B2(n_92),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_94),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_147),
.Y(n_218)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_178),
.A2(n_194),
.B(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_180),
.A2(n_207),
.B1(n_153),
.B2(n_164),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_200),
.B1(n_213),
.B2(n_214),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_160),
.C(n_167),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_170),
.C(n_137),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_98),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_132),
.A2(n_124),
.B1(n_108),
.B2(n_98),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_124),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_138),
.Y(n_230)
);

NOR2x1_ASAP7_75t_R g209 ( 
.A(n_141),
.B(n_142),
.Y(n_209)
);

OR2x2_ASAP7_75t_SL g239 ( 
.A(n_209),
.B(n_137),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_166),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_212),
.Y(n_240)
);

OAI22x1_ASAP7_75t_SL g213 ( 
.A1(n_165),
.A2(n_162),
.B1(n_175),
.B2(n_142),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_162),
.A2(n_148),
.B1(n_133),
.B2(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_147),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_156),
.B1(n_151),
.B2(n_153),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_148),
.B1(n_174),
.B2(n_155),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_226),
.B1(n_236),
.B2(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_221),
.B(n_246),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_160),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_225),
.A2(n_232),
.B(n_238),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_158),
.B1(n_170),
.B2(n_134),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_170),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_135),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_180),
.A2(n_171),
.B1(n_177),
.B2(n_145),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_211),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_153),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_250),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_176),
.B(n_164),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_251),
.B(n_179),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_186),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_209),
.C(n_188),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_218),
.B1(n_214),
.B2(n_182),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_184),
.B1(n_215),
.B2(n_190),
.Y(n_274)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_178),
.B(n_191),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_253),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_200),
.B1(n_183),
.B2(n_202),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_249),
.A2(n_194),
.B1(n_203),
.B2(n_187),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_198),
.B(n_189),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_194),
.A2(n_186),
.B(n_198),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_224),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_257),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_256),
.A2(n_280),
.B1(n_197),
.B2(n_196),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_225),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_247),
.B1(n_231),
.B2(n_243),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_267),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_270),
.C(n_284),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_187),
.B1(n_179),
.B2(n_204),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_260),
.A2(n_274),
.B1(n_237),
.B2(n_228),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_216),
.B(n_204),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_266),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_222),
.A2(n_216),
.B(n_181),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_235),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_231),
.A2(n_190),
.B1(n_206),
.B2(n_199),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_211),
.B(n_181),
.Y(n_281)
);

BUFx12_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_181),
.B(n_211),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_252),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_246),
.C(n_221),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_290),
.C(n_291),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_249),
.B1(n_233),
.B2(n_245),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_295),
.B1(n_297),
.B2(n_255),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_221),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_238),
.C(n_248),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_229),
.C(n_251),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_298),
.C(n_300),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_234),
.B1(n_236),
.B2(n_240),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_229),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_226),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_250),
.A3(n_220),
.B1(n_254),
.B2(n_223),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_278),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_223),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_302),
.B(n_304),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_253),
.C(n_206),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_199),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_199),
.C(n_227),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_227),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_274),
.B1(n_267),
.B2(n_257),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_196),
.B1(n_197),
.B2(n_280),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_309),
.A2(n_281),
.B1(n_260),
.B2(n_266),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_196),
.B1(n_197),
.B2(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_293),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_312),
.A2(n_313),
.B(n_294),
.Y(n_337)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_306),
.B1(n_304),
.B2(n_286),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_319),
.B1(n_330),
.B2(n_285),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_289),
.A2(n_263),
.B(n_270),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_284),
.B(n_289),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_271),
.B1(n_269),
.B2(n_268),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_289),
.A2(n_270),
.B(n_260),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_284),
.B(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_308),
.A2(n_274),
.B1(n_268),
.B2(n_258),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_266),
.B1(n_258),
.B2(n_259),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_291),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_296),
.A2(n_259),
.B1(n_262),
.B2(n_277),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_335),
.A2(n_344),
.B(n_318),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_336),
.B(n_316),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_339),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_300),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_312),
.B(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_287),
.C(n_290),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_343),
.C(n_331),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_323),
.C(n_331),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_322),
.A2(n_294),
.B(n_301),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_345),
.A2(n_347),
.B(n_320),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_348),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_313),
.A2(n_283),
.B(n_264),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_283),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_326),
.B(n_264),
.Y(n_349)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_349),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_350),
.B(n_358),
.Y(n_364)
);

AOI21x1_ASAP7_75t_SL g370 ( 
.A1(n_351),
.A2(n_361),
.B(n_347),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_330),
.C(n_317),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_353),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_328),
.C(n_329),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_333),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_332),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_321),
.C(n_325),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_324),
.C(n_319),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_360),
.B(n_337),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_332),
.A2(n_314),
.B1(n_327),
.B2(n_320),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_338),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

INVx11_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_366),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_371),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_345),
.B(n_359),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_369),
.A2(n_344),
.B(n_352),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_370),
.A2(n_357),
.B(n_362),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_334),
.C(n_335),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_372),
.A2(n_360),
.B(n_273),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_355),
.A2(n_338),
.B1(n_334),
.B2(n_340),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_373),
.A2(n_374),
.B1(n_314),
.B2(n_363),
.Y(n_382)
);

AO21x1_ASAP7_75t_SL g376 ( 
.A1(n_366),
.A2(n_354),
.B(n_340),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_376),
.A2(n_370),
.B(n_362),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_368),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_371),
.B(n_353),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_382),
.Y(n_390)
);

AOI21x1_ASAP7_75t_L g386 ( 
.A1(n_380),
.A2(n_383),
.B(n_369),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_374),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_388),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_381),
.B(n_364),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_385),
.B(n_389),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_387),
.B(n_265),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_381),
.B(n_367),
.Y(n_389)
);

AOI322xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_378),
.A3(n_379),
.B1(n_350),
.B2(n_273),
.C1(n_265),
.C2(n_196),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_391),
.B(n_393),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_394),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_396),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_397),
.A2(n_392),
.B(n_390),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_395),
.Y(n_399)
);


endmodule