module fake_jpeg_21280_n_185 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx10_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_21),
.B1(n_15),
.B2(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_58),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_21),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_14),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_15),
.B1(n_27),
.B2(n_22),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_38),
.B1(n_31),
.B2(n_33),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_28),
.B1(n_25),
.B2(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_51),
.B1(n_42),
.B2(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_42),
.B2(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_17),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_14),
.B(n_2),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_26),
.B(n_20),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_69),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_67),
.Y(n_94)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_44),
.B(n_46),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_73),
.B(n_29),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_75),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_78),
.Y(n_109)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_85),
.Y(n_112)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_14),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_41),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_89),
.B(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_41),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_41),
.C(n_32),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_110),
.B(n_1),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_65),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_74),
.B1(n_80),
.B2(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_120),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_126),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_86),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_77),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_68),
.B(n_3),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_24),
.B(n_4),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_130),
.B1(n_96),
.B2(n_99),
.C(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_122),
.B(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_102),
.B1(n_91),
.B2(n_96),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_127),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_94),
.B1(n_92),
.B2(n_103),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_103),
.B1(n_108),
.B2(n_106),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_126),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_117),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_130),
.A3(n_119),
.B1(n_129),
.B2(n_127),
.C1(n_124),
.C2(n_125),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_150),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_123),
.Y(n_152)
);

OA21x2_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_154),
.B(n_151),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_128),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_144),
.C(n_143),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_160),
.C(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_141),
.C(n_144),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_154),
.B(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_135),
.B1(n_118),
.B2(n_114),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_101),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_167),
.C(n_168),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_170),
.B(n_159),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_145),
.C(n_118),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_142),
.C(n_105),
.Y(n_168)
);

OAI322xp33_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_101),
.A3(n_105),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_1),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_169),
.B1(n_161),
.B2(n_104),
.Y(n_176)
);

NAND4xp25_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_156),
.C(n_158),
.D(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_104),
.Y(n_180)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_173),
.B(n_172),
.C(n_13),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_177),
.B(n_10),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_4),
.B(n_5),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_181),
.A2(n_182),
.B(n_10),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_6),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_6),
.Y(n_185)
);


endmodule