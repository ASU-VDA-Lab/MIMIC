module real_aes_156_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_820, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_819, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_820;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_819;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g529 ( .A(n_0), .B(n_214), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_1), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g142 ( .A(n_2), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_3), .B(n_508), .Y(n_545) );
NAND2xp33_ASAP7_75t_SL g585 ( .A(n_4), .B(n_163), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_5), .B(n_198), .Y(n_205) );
INVx1_ASAP7_75t_L g578 ( .A(n_6), .Y(n_578) );
INVx1_ASAP7_75t_L g185 ( .A(n_7), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g815 ( .A(n_8), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_9), .Y(n_273) );
AND2x2_ASAP7_75t_L g543 ( .A(n_10), .B(n_166), .Y(n_543) );
INVx2_ASAP7_75t_L g134 ( .A(n_11), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g215 ( .A(n_13), .Y(n_215) );
AOI221x1_ASAP7_75t_L g581 ( .A1(n_14), .A2(n_131), .B1(n_510), .B2(n_582), .C(n_584), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_15), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g117 ( .A(n_16), .Y(n_117) );
INVx1_ASAP7_75t_L g212 ( .A(n_17), .Y(n_212) );
INVx1_ASAP7_75t_SL g227 ( .A(n_18), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_19), .B(n_157), .Y(n_201) );
AOI33xp33_ASAP7_75t_L g177 ( .A1(n_20), .A2(n_51), .A3(n_139), .B1(n_150), .B2(n_178), .B3(n_179), .Y(n_177) );
AOI221xp5_ASAP7_75t_SL g519 ( .A1(n_21), .A2(n_42), .B1(n_508), .B2(n_510), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_22), .A2(n_510), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_23), .B(n_214), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_24), .A2(n_103), .B1(n_808), .B2(n_816), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_25), .A2(n_792), .B1(n_793), .B2(n_800), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_25), .Y(n_792) );
INVx1_ASAP7_75t_L g267 ( .A(n_26), .Y(n_267) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_27), .A2(n_90), .B(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g167 ( .A(n_27), .B(n_90), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_28), .B(n_217), .Y(n_513) );
INVxp67_ASAP7_75t_L g580 ( .A(n_29), .Y(n_580) );
AND2x2_ASAP7_75t_L g567 ( .A(n_30), .B(n_165), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_31), .B(n_137), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_32), .A2(n_510), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_33), .B(n_370), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_33), .Y(n_493) );
OAI22x1_ASAP7_75t_R g794 ( .A1(n_33), .A2(n_37), .B1(n_493), .B2(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_34), .B(n_217), .Y(n_521) );
AND2x2_ASAP7_75t_L g144 ( .A(n_35), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g149 ( .A(n_35), .Y(n_149) );
AND2x2_ASAP7_75t_L g163 ( .A(n_35), .B(n_142), .Y(n_163) );
OR2x6_ASAP7_75t_L g115 ( .A(n_36), .B(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_37), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_38), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_39), .B(n_137), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_40), .A2(n_132), .B1(n_194), .B2(n_198), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_41), .B(n_203), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_43), .A2(n_82), .B1(n_147), .B2(n_510), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_44), .B(n_157), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_45), .B(n_214), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_46), .B(n_172), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_47), .B(n_157), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_48), .Y(n_197) );
AND2x2_ASAP7_75t_L g532 ( .A(n_49), .B(n_165), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_50), .B(n_165), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_52), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g140 ( .A(n_53), .Y(n_140) );
INVx1_ASAP7_75t_L g159 ( .A(n_53), .Y(n_159) );
AND2x2_ASAP7_75t_L g164 ( .A(n_54), .B(n_165), .Y(n_164) );
AOI221xp5_ASAP7_75t_L g183 ( .A1(n_55), .A2(n_75), .B1(n_137), .B2(n_147), .C(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_56), .B(n_137), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_57), .B(n_508), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_58), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_59), .B(n_132), .Y(n_275) );
AOI21xp5_ASAP7_75t_SL g235 ( .A1(n_60), .A2(n_147), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g558 ( .A(n_61), .B(n_165), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_62), .B(n_217), .Y(n_530) );
INVx1_ASAP7_75t_L g208 ( .A(n_63), .Y(n_208) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_64), .B(n_166), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_65), .B(n_214), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_66), .A2(n_510), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g154 ( .A(n_67), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_68), .B(n_217), .Y(n_549) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_69), .B(n_172), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_70), .A2(n_147), .B(n_153), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_71), .Y(n_783) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_72), .A2(n_94), .B1(n_109), .B2(n_110), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_72), .Y(n_109) );
INVx1_ASAP7_75t_L g145 ( .A(n_73), .Y(n_145) );
INVx1_ASAP7_75t_L g161 ( .A(n_73), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_74), .B(n_137), .Y(n_180) );
AND2x2_ASAP7_75t_L g229 ( .A(n_76), .B(n_131), .Y(n_229) );
INVx1_ASAP7_75t_L g209 ( .A(n_77), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_78), .A2(n_147), .B(n_226), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_79), .A2(n_147), .B(n_171), .C(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_80), .A2(n_85), .B1(n_137), .B2(n_508), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_81), .B(n_508), .Y(n_557) );
INVx1_ASAP7_75t_L g118 ( .A(n_83), .Y(n_118) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_84), .B(n_131), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_86), .A2(n_147), .B1(n_175), .B2(n_176), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_87), .B(n_214), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_88), .B(n_214), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_89), .A2(n_510), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g237 ( .A(n_91), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_92), .B(n_217), .Y(n_555) );
AND2x2_ASAP7_75t_L g181 ( .A(n_93), .B(n_131), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_94), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_95), .A2(n_265), .B(n_266), .C(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_96), .B(n_508), .Y(n_531) );
INVxp67_ASAP7_75t_L g583 ( .A(n_97), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_98), .B(n_217), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_99), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_SL g106 ( .A(n_100), .Y(n_106) );
BUFx2_ASAP7_75t_L g790 ( .A(n_100), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_101), .B(n_157), .Y(n_238) );
AO21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_786), .B(n_803), .Y(n_103) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_107), .C(n_778), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVxp33_ASAP7_75t_SL g781 ( .A(n_108), .Y(n_781) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_119), .B(n_495), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_112), .A2(n_120), .B1(n_499), .B2(n_780), .Y(n_779) );
CKINVDCx11_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
AND2x6_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OR2x6_ASAP7_75t_SL g497 ( .A(n_114), .B(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g785 ( .A(n_114), .B(n_115), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_114), .B(n_498), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_115), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_490), .Y(n_120) );
NOR4xp25_ASAP7_75t_L g121 ( .A(n_122), .B(n_369), .C(n_393), .D(n_459), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_122), .A2(n_393), .B1(n_493), .B2(n_819), .Y(n_494) );
INVx2_ASAP7_75t_L g799 ( .A(n_122), .Y(n_799) );
NAND3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_321), .C(n_355), .Y(n_122) );
NOR3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_280), .C(n_300), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_255), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_188), .B1(n_244), .B2(n_252), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_168), .Y(n_126) );
AND2x2_ASAP7_75t_L g419 ( .A(n_127), .B(n_349), .Y(n_419) );
INVx1_ASAP7_75t_L g426 ( .A(n_127), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_127), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_127), .B(n_289), .Y(n_478) );
OR2x2_ASAP7_75t_L g488 ( .A(n_127), .B(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_128), .B(n_246), .Y(n_309) );
AND2x4_ASAP7_75t_L g337 ( .A(n_128), .B(n_251), .Y(n_337) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g285 ( .A(n_129), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_129), .B(n_170), .Y(n_375) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_129), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_129), .B(n_262), .Y(n_412) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_135), .B(n_164), .Y(n_129) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_130), .A2(n_135), .B(n_164), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_130), .A2(n_131), .B1(n_264), .B2(n_269), .Y(n_263) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_132), .B(n_272), .Y(n_271) );
AOI21x1_ASAP7_75t_L g525 ( .A1(n_132), .A2(n_526), .B(n_532), .Y(n_525) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_134), .B(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g198 ( .A(n_134), .B(n_167), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_146), .Y(n_135) );
INVx1_ASAP7_75t_L g276 ( .A(n_137), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_137), .A2(n_147), .B1(n_577), .B2(n_579), .Y(n_576) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
OR2x6_ASAP7_75t_L g155 ( .A(n_139), .B(n_151), .Y(n_155) );
INVxp33_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g152 ( .A(n_140), .B(n_142), .Y(n_152) );
AND2x4_ASAP7_75t_L g217 ( .A(n_140), .B(n_160), .Y(n_217) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g196 ( .A(n_143), .Y(n_196) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g510 ( .A(n_144), .B(n_152), .Y(n_510) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
AND2x6_ASAP7_75t_L g214 ( .A(n_145), .B(n_158), .Y(n_214) );
INVxp67_ASAP7_75t_L g274 ( .A(n_147), .Y(n_274) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NOR2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_156), .C(n_162), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g184 ( .A1(n_155), .A2(n_162), .B(n_185), .C(n_186), .Y(n_184) );
INVx2_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_155), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g226 ( .A1(n_155), .A2(n_162), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_155), .A2(n_162), .B(n_237), .C(n_238), .Y(n_236) );
INVxp67_ASAP7_75t_L g265 ( .A(n_155), .Y(n_265) );
INVx1_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
AND2x4_ASAP7_75t_L g508 ( .A(n_157), .B(n_163), .Y(n_508) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_162), .A2(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_162), .B(n_198), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_162), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_162), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_162), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_162), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_162), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_162), .A2(n_564), .B(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_163), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_165), .Y(n_222) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_165), .A2(n_519), .B(n_523), .Y(n_518) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_168), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g483 ( .A(n_168), .B(n_320), .Y(n_483) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_L g473 ( .A(n_169), .B(n_412), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
INVx2_ASAP7_75t_L g251 ( .A(n_170), .Y(n_251) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_181), .Y(n_170) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_171), .A2(n_173), .B(n_181), .Y(n_279) );
AOI21x1_ASAP7_75t_L g536 ( .A1(n_171), .A2(n_537), .B(n_540), .Y(n_536) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_172), .A2(n_183), .B(n_187), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_172), .A2(n_507), .B(n_509), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_174), .B(n_180), .Y(n_173) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
INVx2_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_182), .Y(n_286) );
INVx1_ASAP7_75t_L g299 ( .A(n_182), .Y(n_299) );
INVxp67_ASAP7_75t_L g318 ( .A(n_182), .Y(n_318) );
AND2x4_ASAP7_75t_L g349 ( .A(n_182), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_230), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_219), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g391 ( .A(n_191), .B(n_378), .Y(n_391) );
AND2x2_ASAP7_75t_L g415 ( .A(n_191), .B(n_231), .Y(n_415) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_204), .Y(n_191) );
INVx2_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
INVx1_ASAP7_75t_L g315 ( .A(n_192), .Y(n_315) );
AND2x4_ASAP7_75t_L g324 ( .A(n_192), .B(n_242), .Y(n_324) );
AND2x2_ASAP7_75t_L g380 ( .A(n_192), .B(n_232), .Y(n_380) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_199), .Y(n_192) );
NOR3xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .C(n_197), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_198), .A2(n_235), .B(n_239), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_198), .A2(n_545), .B(n_546), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_198), .B(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_198), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_198), .B(n_583), .Y(n_582) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_198), .B(n_210), .C(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
AND2x2_ASAP7_75t_L g254 ( .A(n_204), .B(n_221), .Y(n_254) );
INVx2_ASAP7_75t_L g293 ( .A(n_204), .Y(n_293) );
NOR2x1_ASAP7_75t_SL g306 ( .A(n_204), .B(n_232), .Y(n_306) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_211), .B(n_218), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_210), .B(n_267), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B1(n_215), .B2(n_216), .Y(n_211) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g408 ( .A(n_219), .Y(n_408) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g331 ( .A(n_220), .Y(n_331) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_221), .Y(n_289) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_221), .Y(n_305) );
AND2x2_ASAP7_75t_L g313 ( .A(n_221), .B(n_242), .Y(n_313) );
INVx1_ASAP7_75t_L g353 ( .A(n_221), .Y(n_353) );
INVx1_ASAP7_75t_L g378 ( .A(n_221), .Y(n_378) );
OR2x2_ASAP7_75t_L g439 ( .A(n_221), .B(n_232), .Y(n_439) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_221) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_222), .A2(n_552), .B(n_558), .Y(n_551) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_222), .A2(n_561), .B(n_567), .Y(n_560) );
AO21x2_ASAP7_75t_L g605 ( .A1(n_222), .A2(n_561), .B(n_567), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
OA211x2_ASAP7_75t_L g460 ( .A1(n_230), .A2(n_461), .B(n_463), .C(n_470), .Y(n_460) );
OR2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_240), .Y(n_230) );
AND2x2_ASAP7_75t_L g381 ( .A(n_231), .B(n_254), .Y(n_381) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_231), .B(n_241), .Y(n_399) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx4_ASAP7_75t_L g253 ( .A(n_232), .Y(n_253) );
INVx2_ASAP7_75t_L g295 ( .A(n_232), .Y(n_295) );
AND2x4_ASAP7_75t_L g358 ( .A(n_232), .B(n_315), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_232), .B(n_354), .Y(n_409) );
AND2x2_ASAP7_75t_L g452 ( .A(n_232), .B(n_293), .Y(n_452) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_241), .B(n_353), .Y(n_446) );
AND2x2_ASAP7_75t_L g466 ( .A(n_241), .B(n_289), .Y(n_466) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g354 ( .A(n_242), .Y(n_354) );
INVx1_ASAP7_75t_L g328 ( .A(n_243), .Y(n_328) );
NOR2xp67_ASAP7_75t_SL g244 ( .A(n_245), .B(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g422 ( .A(n_245), .Y(n_422) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_245), .B(n_423), .Y(n_469) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g442 ( .A(n_247), .B(n_284), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_248), .A2(n_431), .B(n_434), .C(n_443), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_248), .A2(n_468), .B(n_475), .C(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g359 ( .A(n_249), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g278 ( .A(n_250), .Y(n_278) );
NOR2x1_ASAP7_75t_L g298 ( .A(n_250), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g334 ( .A(n_250), .B(n_284), .Y(n_334) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_250), .B(n_284), .Y(n_444) );
AND2x2_ASAP7_75t_L g317 ( .A(n_251), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g368 ( .A(n_251), .Y(n_368) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x4_ASAP7_75t_SL g257 ( .A(n_253), .B(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g314 ( .A(n_253), .B(n_315), .Y(n_314) );
NOR2x1_ASAP7_75t_L g343 ( .A(n_253), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g362 ( .A(n_253), .B(n_363), .Y(n_362) );
NOR2xp67_ASAP7_75t_SL g445 ( .A(n_253), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_254), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_SL g485 ( .A(n_254), .B(n_327), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
INVx2_ASAP7_75t_SL g453 ( .A(n_259), .Y(n_453) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_277), .Y(n_259) );
INVx3_ASAP7_75t_L g376 ( .A(n_260), .Y(n_376) );
AND2x2_ASAP7_75t_L g397 ( .A(n_260), .B(n_388), .Y(n_397) );
AND2x2_ASAP7_75t_L g455 ( .A(n_260), .B(n_337), .Y(n_455) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g284 ( .A(n_262), .Y(n_284) );
INVx1_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
INVx1_ASAP7_75t_L g340 ( .A(n_262), .Y(n_340) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B1(n_275), .B2(n_276), .Y(n_270) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g423 ( .A(n_277), .Y(n_423) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g283 ( .A(n_279), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g350 ( .A(n_279), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_287), .B1(n_290), .B2(n_296), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g357 ( .A(n_288), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g377 ( .A(n_292), .B(n_378), .Y(n_377) );
NOR2x1_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g385 ( .A(n_293), .Y(n_385) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g433 ( .A(n_295), .B(n_324), .Y(n_433) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_297), .A2(n_391), .B(n_392), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B(n_310), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_330), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_307), .A2(n_414), .B1(n_416), .B2(n_418), .Y(n_413) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_316), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_SL g363 ( .A(n_313), .Y(n_363) );
AND2x2_ASAP7_75t_L g392 ( .A(n_314), .B(n_330), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_314), .B(n_352), .Y(n_424) );
AND2x2_ASAP7_75t_L g428 ( .A(n_314), .B(n_385), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_316), .A2(n_373), .B(n_377), .Y(n_372) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x2_ASAP7_75t_L g333 ( .A(n_317), .B(n_334), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_317), .B(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g402 ( .A(n_320), .Y(n_402) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_345), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_332), .B1(n_335), .B2(n_341), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx4_ASAP7_75t_L g344 ( .A(n_324), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_324), .B(n_330), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_324), .B(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_327), .A2(n_351), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g450 ( .A(n_327), .B(n_352), .Y(n_450) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g432 ( .A(n_329), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g468 ( .A(n_330), .B(n_452), .Y(n_468) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g348 ( .A(n_334), .B(n_349), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_334), .B(n_368), .Y(n_367) );
OAI22xp5_ASAP7_75t_SL g345 ( .A1(n_335), .A2(n_346), .B1(n_347), .B2(n_351), .Y(n_345) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g462 ( .A(n_339), .B(n_349), .Y(n_462) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g360 ( .A(n_340), .Y(n_360) );
AND2x2_ASAP7_75t_L g386 ( .A(n_340), .B(n_349), .Y(n_386) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_342), .B(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_343), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g437 ( .A(n_344), .Y(n_437) );
INVx1_ASAP7_75t_L g449 ( .A(n_346), .Y(n_449) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_348), .A2(n_392), .B1(n_471), .B2(n_472), .Y(n_470) );
AND2x2_ASAP7_75t_L g387 ( .A(n_349), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g458 ( .A(n_349), .B(n_411), .Y(n_458) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI211xp5_ASAP7_75t_SL g361 ( .A1(n_352), .A2(n_362), .B(n_364), .C(n_365), .Y(n_361) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_352), .B(n_358), .Y(n_471) );
AND2x4_ASAP7_75t_SL g352 ( .A(n_353), .B(n_354), .Y(n_352) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_353), .Y(n_405) );
O2A1O1Ixp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B(n_359), .C(n_361), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_356), .A2(n_384), .B1(n_386), .B2(n_387), .Y(n_383) );
INVx2_ASAP7_75t_L g364 ( .A(n_358), .Y(n_364) );
AND2x2_ASAP7_75t_L g384 ( .A(n_358), .B(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_358), .Y(n_451) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g492 ( .A(n_370), .Y(n_492) );
NAND4xp75_ASAP7_75t_L g796 ( .A(n_370), .B(n_797), .C(n_798), .D(n_799), .Y(n_796) );
NOR2x1_ASAP7_75t_SL g370 ( .A(n_371), .B(n_382), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_379), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_373), .A2(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
INVx1_ASAP7_75t_L g479 ( .A(n_376), .Y(n_479) );
AND2x2_ASAP7_75t_L g417 ( .A(n_380), .B(n_405), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_381), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_383), .B(n_390), .Y(n_382) );
AND2x2_ASAP7_75t_L g484 ( .A(n_386), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g797 ( .A(n_393), .Y(n_797) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_429), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_413), .C(n_420), .Y(n_394) );
OAI222xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B1(n_400), .B2(n_404), .C1(n_406), .C2(n_410), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .B1(n_425), .B2(n_427), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR2xp67_ASAP7_75t_SL g429 ( .A(n_430), .B(n_447), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_437), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g489 ( .A(n_442), .Y(n_489) );
NAND2xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_453), .B1(n_454), .B2(n_456), .C(n_457), .Y(n_447) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .C(n_451), .D(n_452), .Y(n_448) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_459), .A2(n_492), .B(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g798 ( .A(n_459), .Y(n_798) );
NAND4xp75_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .C(n_480), .D(n_486), .Y(n_459) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_464), .B(n_469), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_484), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .Y(n_490) );
NAND2x1_ASAP7_75t_SL g495 ( .A(n_496), .B(n_499), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_496), .Y(n_780) );
CKINVDCx11_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_670), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_598), .C(n_648), .Y(n_501) );
OAI211xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_533), .B(n_568), .C(n_587), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
AND2x2_ASAP7_75t_L g597 ( .A(n_504), .B(n_516), .Y(n_597) );
INVx1_ASAP7_75t_L g728 ( .A(n_504), .Y(n_728) );
NOR2x1p5_ASAP7_75t_L g760 ( .A(n_504), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g573 ( .A(n_505), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g619 ( .A(n_505), .Y(n_619) );
OR2x2_ASAP7_75t_L g623 ( .A(n_505), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_505), .B(n_518), .Y(n_635) );
OR2x2_ASAP7_75t_L g657 ( .A(n_505), .B(n_518), .Y(n_657) );
AND2x4_ASAP7_75t_L g663 ( .A(n_505), .B(n_627), .Y(n_663) );
OR2x2_ASAP7_75t_L g680 ( .A(n_505), .B(n_575), .Y(n_680) );
INVx1_ASAP7_75t_L g715 ( .A(n_505), .Y(n_715) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_505), .Y(n_737) );
OR2x2_ASAP7_75t_L g751 ( .A(n_505), .B(n_684), .Y(n_751) );
AND2x4_ASAP7_75t_SL g755 ( .A(n_505), .B(n_575), .Y(n_755) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g707 ( .A(n_516), .B(n_663), .Y(n_707) );
AND2x2_ASAP7_75t_L g754 ( .A(n_516), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g572 ( .A(n_518), .Y(n_572) );
AND2x2_ASAP7_75t_L g617 ( .A(n_518), .B(n_524), .Y(n_617) );
INVx2_ASAP7_75t_L g624 ( .A(n_518), .Y(n_624) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_518), .Y(n_745) );
BUFx3_ASAP7_75t_L g761 ( .A(n_518), .Y(n_761) );
INVx2_ASAP7_75t_L g586 ( .A(n_524), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_524), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g684 ( .A(n_524), .B(n_624), .Y(n_684) );
INVx1_ASAP7_75t_L g702 ( .A(n_524), .Y(n_702) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_524), .Y(n_718) );
INVx1_ASAP7_75t_L g740 ( .A(n_524), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_524), .B(n_619), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_524), .B(n_575), .Y(n_777) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_541), .Y(n_534) );
AND2x4_ASAP7_75t_L g591 ( .A(n_535), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_535), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g642 ( .A(n_535), .B(n_550), .Y(n_642) );
AND2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_551), .Y(n_652) );
OR2x2_ASAP7_75t_L g732 ( .A(n_535), .B(n_647), .Y(n_732) );
OAI322xp33_ASAP7_75t_L g762 ( .A1(n_535), .A2(n_675), .A3(n_714), .B1(n_747), .B2(n_763), .C1(n_764), .C2(n_765), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_535), .B(n_745), .Y(n_763) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g596 ( .A(n_536), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_541), .A2(n_709), .B1(n_713), .B2(n_716), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g768 ( .A1(n_541), .A2(n_769), .B(n_770), .C(n_773), .Y(n_768) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_542), .B(n_550), .Y(n_541) );
AND2x4_ASAP7_75t_L g590 ( .A(n_542), .B(n_560), .Y(n_590) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_542), .Y(n_594) );
INVx5_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
INVx2_ASAP7_75t_L g615 ( .A(n_542), .Y(n_615) );
AND2x2_ASAP7_75t_L g638 ( .A(n_542), .B(n_551), .Y(n_638) );
AND2x2_ASAP7_75t_L g667 ( .A(n_542), .B(n_559), .Y(n_667) );
OR2x2_ASAP7_75t_L g676 ( .A(n_542), .B(n_596), .Y(n_676) );
OR2x2_ASAP7_75t_L g691 ( .A(n_542), .B(n_605), .Y(n_691) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_550), .B(n_569), .Y(n_568) );
INVx3_ASAP7_75t_SL g675 ( .A(n_550), .Y(n_675) );
AND2x2_ASAP7_75t_L g698 ( .A(n_550), .B(n_606), .Y(n_698) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_559), .Y(n_550) );
INVx2_ASAP7_75t_L g592 ( .A(n_551), .Y(n_592) );
AND2x2_ASAP7_75t_L g595 ( .A(n_551), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g609 ( .A(n_551), .B(n_560), .Y(n_609) );
INVx1_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_551), .B(n_560), .Y(n_647) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_551), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_551), .B(n_606), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_560), .Y(n_628) );
AND2x2_ASAP7_75t_L g712 ( .A(n_560), .B(n_596), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_570), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x6_ASAP7_75t_SL g776 ( .A(n_571), .B(n_777), .Y(n_776) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_572), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_572), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g724 ( .A(n_572), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_573), .A2(n_633), .B1(n_636), .B2(n_643), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_574), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g668 ( .A(n_574), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_574), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_574), .B(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_586), .Y(n_574) );
AND2x2_ASAP7_75t_L g618 ( .A(n_575), .B(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g627 ( .A(n_575), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_575), .A2(n_634), .B1(n_686), .B2(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g693 ( .A(n_575), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_575), .B(n_687), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_575), .B(n_617), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_575), .B(n_624), .Y(n_766) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_581), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_593), .B(n_597), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
NAND4xp25_ASAP7_75t_SL g636 ( .A(n_589), .B(n_637), .C(n_639), .D(n_641), .Y(n_636) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_590), .B(n_697), .Y(n_726) );
AND2x2_ASAP7_75t_L g753 ( .A(n_590), .B(n_591), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_590), .B(n_613), .Y(n_764) );
INVx1_ASAP7_75t_L g629 ( .A(n_591), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_591), .A2(n_654), .B1(n_665), .B2(n_668), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_591), .B(n_604), .C(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_591), .B(n_606), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_591), .B(n_614), .Y(n_757) );
AND2x2_ASAP7_75t_L g689 ( .A(n_592), .B(n_596), .Y(n_689) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_592), .Y(n_750) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g645 ( .A(n_594), .Y(n_645) );
INVx1_ASAP7_75t_L g735 ( .A(n_595), .Y(n_735) );
AND2x2_ASAP7_75t_L g742 ( .A(n_595), .B(n_606), .Y(n_742) );
BUFx2_ASAP7_75t_L g697 ( .A(n_596), .Y(n_697) );
NAND3xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_620), .C(n_632), .Y(n_598) );
OAI31xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_607), .A3(n_610), .B(n_616), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_600), .A2(n_654), .B1(n_658), .B2(n_659), .Y(n_653) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OR2x2_ASAP7_75t_L g639 ( .A(n_602), .B(n_640), .Y(n_639) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_602), .B(n_666), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_603), .A2(n_705), .B(n_735), .C(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_604), .B(n_750), .Y(n_749) );
AND2x4_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_605), .B(n_613), .Y(n_640) );
AND2x2_ASAP7_75t_L g658 ( .A(n_605), .B(n_638), .Y(n_658) );
AND2x2_ASAP7_75t_L g775 ( .A(n_608), .B(n_697), .Y(n_775) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g631 ( .A(n_609), .B(n_615), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g706 ( .A(n_614), .B(n_689), .Y(n_706) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_615), .B(n_689), .Y(n_695) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx2_ASAP7_75t_L g687 ( .A(n_617), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_618), .B(n_718), .Y(n_717) );
AOI32xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_628), .A3(n_629), .B1(n_630), .B2(n_820), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_621), .A2(n_706), .B1(n_742), .B2(n_743), .C(n_746), .Y(n_741) );
AND2x4_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_624), .Y(n_669) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g634 ( .A(n_626), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g739 ( .A(n_627), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_628), .B(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_630), .A2(n_673), .B1(n_677), .B2(n_681), .C(n_685), .Y(n_672) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g648 ( .A1(n_635), .A2(n_649), .B(n_653), .C(n_664), .Y(n_648) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI322xp33_ASAP7_75t_L g746 ( .A1(n_641), .A2(n_651), .A3(n_700), .B1(n_747), .B2(n_748), .C1(n_749), .C2(n_751), .Y(n_746) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI21xp33_ASAP7_75t_L g773 ( .A1(n_644), .A2(n_774), .B(n_776), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g730 ( .A1(n_650), .A2(n_731), .B(n_733), .C(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g772 ( .A(n_657), .B(n_738), .Y(n_772) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_663), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g747 ( .A(n_663), .Y(n_747) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI31xp33_ASAP7_75t_L g703 ( .A1(n_667), .A2(n_704), .A3(n_706), .B(n_707), .Y(n_703) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_729), .Y(n_670) );
NAND5xp2_ASAP7_75t_L g671 ( .A(n_672), .B(n_692), .C(n_703), .D(n_708), .E(n_719), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g770 ( .A1(n_675), .A2(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g743 ( .A(n_679), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_696), .C(n_699), .Y(n_692) );
INVxp33_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OR2x2_ASAP7_75t_L g721 ( .A(n_697), .B(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_700), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g771 ( .A(n_712), .Y(n_771) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_725), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI21xp33_ASAP7_75t_L g725 ( .A1(n_721), .A2(n_726), .B(n_727), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_730), .B(n_741), .C(n_752), .D(n_768), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_739), .B(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g769 ( .A(n_751), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_756), .B2(n_758), .C(n_762), .Y(n_752) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_781), .B(n_782), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
BUFx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI21xp5_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_791), .B(n_801), .Y(n_786) );
BUFx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2x1_ASAP7_75t_R g801 ( .A(n_790), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g800 ( .A(n_793), .Y(n_800) );
XNOR2x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
BUFx3_ASAP7_75t_L g807 ( .A(n_802), .Y(n_807) );
BUFx2_ASAP7_75t_L g812 ( .A(n_802), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_SL g817 ( .A(n_810), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
endmodule