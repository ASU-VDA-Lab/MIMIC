module real_aes_6938_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_1), .A2(n_146), .B(n_158), .C(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g265 ( .A(n_2), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_3), .A2(n_173), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_4), .B(n_169), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g172 ( .A1(n_5), .A2(n_173), .B(n_174), .Y(n_172) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_7), .A2(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_8), .B(n_44), .Y(n_117) );
INVx1_ASAP7_75t_L g473 ( .A(n_9), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_10), .B(n_179), .Y(n_461) );
INVx1_ASAP7_75t_L g181 ( .A(n_11), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_12), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g143 ( .A(n_13), .Y(n_143) );
INVx1_ASAP7_75t_L g247 ( .A(n_14), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_16), .A2(n_182), .B(n_248), .C(n_482), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_17), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_17), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_18), .B(n_169), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_19), .B(n_192), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_20), .B(n_173), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_21), .B(n_515), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_22), .A2(n_149), .B(n_233), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_23), .B(n_169), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_24), .B(n_179), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_25), .A2(n_245), .B(n_246), .C(n_248), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_26), .B(n_179), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_27), .Y(n_532) );
INVx1_ASAP7_75t_L g522 ( .A(n_28), .Y(n_522) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_29), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_30), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_31), .B(n_179), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g104 ( .A1(n_32), .A2(n_105), .B1(n_735), .B2(n_741), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_33), .A2(n_67), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_33), .Y(n_731) );
INVx1_ASAP7_75t_L g511 ( .A(n_34), .Y(n_511) );
INVx1_ASAP7_75t_L g157 ( .A(n_35), .Y(n_157) );
AOI222xp33_ASAP7_75t_SL g118 ( .A1(n_36), .A2(n_119), .B1(n_120), .B2(n_129), .C1(n_715), .C2(n_718), .Y(n_118) );
INVx2_ASAP7_75t_L g151 ( .A(n_37), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_38), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_39), .A2(n_183), .B(n_233), .C(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g512 ( .A(n_40), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_41), .A2(n_146), .B(n_158), .C(n_203), .Y(n_202) );
CKINVDCx14_ASAP7_75t_R g498 ( .A(n_42), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_43), .A2(n_158), .B(n_521), .C(n_525), .Y(n_520) );
INVx1_ASAP7_75t_L g155 ( .A(n_45), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_46), .A2(n_178), .B(n_208), .C(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_47), .B(n_179), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_48), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_49), .Y(n_508) );
INVx1_ASAP7_75t_L g488 ( .A(n_50), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_51), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_52), .B(n_173), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_53), .A2(n_149), .B1(n_152), .B2(n_158), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_54), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_55), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_56), .A2(n_178), .B(n_180), .C(n_183), .Y(n_177) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_57), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_58), .Y(n_222) );
INVx1_ASAP7_75t_L g175 ( .A(n_59), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_60), .A2(n_728), .B1(n_729), .B2(n_732), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_60), .Y(n_732) );
INVx1_ASAP7_75t_L g147 ( .A(n_61), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_62), .A2(n_78), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_62), .Y(n_127) );
INVx1_ASAP7_75t_L g142 ( .A(n_63), .Y(n_142) );
INVx1_ASAP7_75t_SL g501 ( .A(n_64), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_65), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_66), .B(n_169), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_67), .Y(n_730) );
INVx1_ASAP7_75t_L g535 ( .A(n_68), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_SL g191 ( .A1(n_69), .A2(n_183), .B(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_70), .Y(n_194) );
INVx1_ASAP7_75t_L g739 ( .A(n_71), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_72), .A2(n_173), .B(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_73), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_74), .Y(n_166) );
OAI22xp33_ASAP7_75t_SL g724 ( .A1(n_74), .A2(n_166), .B1(n_725), .B2(n_726), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_75), .A2(n_173), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g215 ( .A(n_76), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_77), .A2(n_241), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_78), .Y(n_126) );
INVx1_ASAP7_75t_L g480 ( .A(n_79), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_80), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_81), .A2(n_146), .B(n_158), .C(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_82), .A2(n_173), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g483 ( .A(n_83), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_84), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
INVx1_ASAP7_75t_L g459 ( .A(n_86), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_87), .B(n_192), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_88), .A2(n_146), .B(n_158), .C(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g113 ( .A(n_89), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g446 ( .A(n_89), .Y(n_446) );
OR2x2_ASAP7_75t_L g714 ( .A(n_89), .B(n_115), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_90), .A2(n_158), .B(n_534), .C(n_537), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_91), .B(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_92), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_93), .A2(n_146), .B(n_158), .C(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_94), .Y(n_237) );
INVx1_ASAP7_75t_L g190 ( .A(n_95), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_96), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_97), .B(n_205), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_98), .B(n_171), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_99), .B(n_171), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_100), .A2(n_173), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g491 ( .A(n_101), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_102), .B(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_103), .A2(n_121), .B1(n_122), .B2(n_128), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_103), .Y(n_128) );
AOI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_118), .B1(n_722), .B2(n_723), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g722 ( .A(n_108), .Y(n_722) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_110), .A2(n_724), .B(n_733), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g734 ( .A(n_113), .Y(n_734) );
INVx1_ASAP7_75t_SL g740 ( .A(n_113), .Y(n_740) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_114), .B(n_446), .Y(n_717) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g445 ( .A(n_115), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_443), .B1(n_447), .B2(n_714), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_131), .A2(n_443), .B1(n_719), .B2(n_720), .Y(n_718) );
AND3x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_368), .C(n_417), .Y(n_131) );
NOR3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_275), .C(n_313), .Y(n_132) );
OAI222xp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_196), .B1(n_250), .B2(n_256), .C1(n_270), .C2(n_273), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_167), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_135), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_135), .B(n_318), .Y(n_409) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g286 ( .A(n_136), .B(n_187), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_136), .B(n_168), .Y(n_294) );
AND2x2_ASAP7_75t_L g329 ( .A(n_136), .B(n_306), .Y(n_329) );
OR2x2_ASAP7_75t_L g353 ( .A(n_136), .B(n_168), .Y(n_353) );
OR2x2_ASAP7_75t_L g361 ( .A(n_136), .B(n_260), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_136), .B(n_187), .Y(n_364) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g258 ( .A(n_137), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_137), .B(n_187), .Y(n_272) );
AND2x2_ASAP7_75t_L g322 ( .A(n_137), .B(n_260), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_137), .B(n_168), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_137), .B(n_421), .Y(n_442) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_165), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_138), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_138), .A2(n_261), .B(n_268), .Y(n_260) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_140), .B(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B1(n_161), .B2(n_162), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_145), .A2(n_175), .B(n_176), .C(n_177), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_145), .A2(n_176), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_145), .A2(n_176), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g469 ( .A1(n_145), .A2(n_176), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_145), .A2(n_176), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g487 ( .A1(n_145), .A2(n_176), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_145), .A2(n_176), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_145), .A2(n_176), .B(n_508), .C(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g537 ( .A(n_145), .Y(n_537) );
INVx4_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_146), .B(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g173 ( .A(n_146), .B(n_163), .Y(n_173) );
BUFx3_ASAP7_75t_L g525 ( .A(n_146), .Y(n_525) );
INVx2_ASAP7_75t_L g267 ( .A(n_149), .Y(n_267) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx1_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g152 ( .A1(n_153), .A2(n_155), .B1(n_156), .B2(n_157), .Y(n_152) );
INVx2_ASAP7_75t_L g156 ( .A(n_153), .Y(n_156) );
INVx4_ASAP7_75t_L g245 ( .A(n_153), .Y(n_245) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
AND2x2_ASAP7_75t_L g163 ( .A(n_154), .B(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx3_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx2_ASAP7_75t_L g460 ( .A(n_156), .Y(n_460) );
INVx5_ASAP7_75t_L g176 ( .A(n_158), .Y(n_176) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
BUFx3_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_162), .A2(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_162), .A2(n_262), .B(n_263), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_162), .A2(n_456), .B(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_162), .A2(n_186), .B(n_519), .C(n_520), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_162), .A2(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g513 ( .A(n_164), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_167), .A2(n_361), .B(n_362), .C(n_365), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_167), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_167), .B(n_305), .Y(n_427) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_187), .Y(n_167) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_168), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g285 ( .A(n_168), .Y(n_285) );
AND2x2_ASAP7_75t_L g312 ( .A(n_168), .B(n_306), .Y(n_312) );
INVx1_ASAP7_75t_SL g320 ( .A(n_168), .Y(n_320) );
AND2x2_ASAP7_75t_L g343 ( .A(n_168), .B(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g421 ( .A(n_168), .Y(n_421) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_185), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_170), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_170), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_170), .B(n_527), .Y(n_526) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_170), .A2(n_531), .B(n_538), .Y(n_530) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_171), .A2(n_188), .B(n_195), .Y(n_187) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_171), .Y(n_477) );
BUFx2_ASAP7_75t_L g241 ( .A(n_173), .Y(n_241) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_182), .B(n_194), .Y(n_193) );
INVx5_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_182), .B(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
INVx1_ASAP7_75t_L g223 ( .A(n_186), .Y(n_223) );
INVx2_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_186), .A2(n_240), .B(n_249), .Y(n_239) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_186), .A2(n_468), .B(n_474), .Y(n_467) );
BUFx2_ASAP7_75t_L g257 ( .A(n_187), .Y(n_257) );
INVx1_ASAP7_75t_L g319 ( .A(n_187), .Y(n_319) );
INVx3_ASAP7_75t_L g344 ( .A(n_187), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_196), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_224), .Y(n_196) );
INVx1_ASAP7_75t_L g340 ( .A(n_197), .Y(n_340) );
OAI32xp33_ASAP7_75t_L g346 ( .A1(n_197), .A2(n_285), .A3(n_347), .B1(n_348), .B2(n_349), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_197), .A2(n_351), .B1(n_354), .B2(n_359), .Y(n_350) );
INVx4_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g288 ( .A(n_198), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g366 ( .A(n_198), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g436 ( .A(n_198), .B(n_382), .Y(n_436) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
AND2x2_ASAP7_75t_L g251 ( .A(n_199), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g281 ( .A(n_199), .Y(n_281) );
INVx1_ASAP7_75t_L g300 ( .A(n_199), .Y(n_300) );
OR2x2_ASAP7_75t_L g308 ( .A(n_199), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_199), .B(n_289), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_199), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g336 ( .A(n_199), .B(n_254), .Y(n_336) );
INVx3_ASAP7_75t_L g358 ( .A(n_199), .Y(n_358) );
AND2x2_ASAP7_75t_L g383 ( .A(n_199), .B(n_255), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_199), .B(n_348), .Y(n_431) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_211), .Y(n_199) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_202), .B(n_210), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B(n_207), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_205), .A2(n_265), .B(n_266), .C(n_267), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_205), .A2(n_245), .B1(n_511), .B2(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_205), .A2(n_522), .B(n_523), .C(n_524), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_207), .A2(n_218), .B(n_219), .Y(n_217) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_207), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_207), .A2(n_460), .B(n_535), .C(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
INVx1_ASAP7_75t_L g220 ( .A(n_210), .Y(n_220) );
INVx2_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
AND2x2_ASAP7_75t_L g387 ( .A(n_213), .B(n_225), .Y(n_387) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_213) );
INVx1_ASAP7_75t_L g505 ( .A(n_220), .Y(n_505) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_220), .A2(n_558), .B(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_223), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_223), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_223), .A2(n_455), .B(n_462), .Y(n_454) );
INVx2_ASAP7_75t_L g429 ( .A(n_224), .Y(n_429) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_238), .Y(n_224) );
INVx1_ASAP7_75t_L g274 ( .A(n_225), .Y(n_274) );
AND2x2_ASAP7_75t_L g301 ( .A(n_225), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_225), .B(n_255), .Y(n_309) );
AND2x2_ASAP7_75t_L g367 ( .A(n_225), .B(n_290), .Y(n_367) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g253 ( .A(n_226), .Y(n_253) );
AND2x2_ASAP7_75t_L g280 ( .A(n_226), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g289 ( .A(n_226), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_226), .B(n_255), .Y(n_355) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_236), .Y(n_226) );
INVx1_ASAP7_75t_L g515 ( .A(n_227), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_227), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_234), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_233), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_238), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_238), .B(n_255), .Y(n_348) );
AND2x2_ASAP7_75t_L g357 ( .A(n_238), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g382 ( .A(n_238), .Y(n_382) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g254 ( .A(n_239), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g290 ( .A(n_239), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_245), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_245), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_245), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_250), .A2(n_260), .B1(n_419), .B2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_252), .A2(n_363), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_253), .B(n_358), .Y(n_375) );
INVx1_ASAP7_75t_L g400 ( .A(n_253), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_254), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g327 ( .A(n_254), .B(n_280), .Y(n_327) );
INVx2_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
INVx1_ASAP7_75t_L g333 ( .A(n_255), .Y(n_333) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_256), .A2(n_408), .B1(n_425), .B2(n_428), .C(n_430), .Y(n_424) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_257), .B(n_306), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_258), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g349 ( .A(n_258), .B(n_295), .Y(n_349) );
INVx3_ASAP7_75t_SL g390 ( .A(n_258), .Y(n_390) );
AND2x2_ASAP7_75t_L g334 ( .A(n_259), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g363 ( .A(n_259), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_259), .B(n_272), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_259), .B(n_318), .Y(n_404) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g306 ( .A(n_260), .Y(n_306) );
OAI322xp33_ASAP7_75t_L g401 ( .A1(n_260), .A2(n_332), .A3(n_354), .B1(n_402), .B2(n_404), .C1(n_405), .C2(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_271), .A2(n_274), .B(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_272), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g373 ( .A(n_272), .B(n_285), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_272), .B(n_312), .Y(n_388) );
INVxp67_ASAP7_75t_L g339 ( .A(n_274), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_274), .A2(n_346), .B(n_350), .C(n_360), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g275 ( .A1(n_276), .A2(n_284), .B1(n_287), .B2(n_291), .C(n_296), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g299 ( .A(n_283), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g416 ( .A(n_283), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_284), .A2(n_433), .B1(n_438), .B2(n_439), .C(n_441), .Y(n_432) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g332 ( .A(n_285), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_285), .B(n_363), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_285), .B(n_390), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_286), .B(n_311), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_286), .A2(n_298), .B1(n_408), .B2(n_409), .Y(n_407) );
OR2x2_ASAP7_75t_L g438 ( .A(n_286), .B(n_306), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g415 ( .A(n_289), .Y(n_415) );
AND2x2_ASAP7_75t_L g440 ( .A(n_289), .B(n_383), .Y(n_440) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g304 ( .A(n_294), .B(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_303), .B1(n_307), .B2(n_310), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g371 ( .A(n_299), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_299), .B(n_339), .Y(n_406) );
AOI322xp5_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_331), .A3(n_333), .B1(n_334), .B2(n_336), .C1(n_337), .C2(n_341), .Y(n_330) );
INVxp67_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_304), .A2(n_309), .B1(n_326), .B2(n_328), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_305), .B(n_318), .Y(n_405) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_306), .B(n_344), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_306), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g402 ( .A(n_308), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NAND3xp33_ASAP7_75t_SL g313 ( .A(n_314), .B(n_330), .C(n_345), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_321), .B2(n_323), .C(n_325), .Y(n_314) );
AND2x2_ASAP7_75t_L g321 ( .A(n_317), .B(n_322), .Y(n_321) );
INVx3_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_324), .Y(n_403) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_329), .B(n_343), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_332), .B(n_390), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_333), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g408 ( .A(n_336), .Y(n_408) );
AND2x2_ASAP7_75t_L g423 ( .A(n_336), .B(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_347), .A2(n_418), .B(n_424), .C(n_432), .Y(n_417) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g386 ( .A(n_357), .B(n_387), .Y(n_386) );
NAND2x1_ASAP7_75t_SL g428 ( .A(n_358), .B(n_429), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g393 ( .A(n_367), .Y(n_393) );
AND2x2_ASAP7_75t_L g397 ( .A(n_367), .B(n_383), .Y(n_397) );
NOR5xp2_ASAP7_75t_L g368 ( .A(n_369), .B(n_384), .C(n_401), .D(n_407), .E(n_410), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_372), .B2(n_374), .C(n_376), .Y(n_369) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_373), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g399 ( .A(n_383), .B(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_388), .B1(n_389), .B2(n_391), .C(n_394), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
AOI211xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_413), .B(n_415), .C(n_416), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
CKINVDCx14_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g719 ( .A(n_447), .Y(n_719) );
XNOR2xp5_ASAP7_75t_L g726 ( .A(n_447), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_669), .Y(n_447) );
NAND5xp2_ASAP7_75t_L g448 ( .A(n_449), .B(n_581), .C(n_619), .D(n_640), .E(n_657), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_553), .C(n_574), .Y(n_449) );
OAI221xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_493), .B1(n_516), .B2(n_540), .C(n_544), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_464), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_453), .B(n_542), .Y(n_561) );
OR2x2_ASAP7_75t_L g588 ( .A(n_453), .B(n_476), .Y(n_588) );
AND2x2_ASAP7_75t_L g602 ( .A(n_453), .B(n_476), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_453), .B(n_467), .Y(n_616) );
AND2x2_ASAP7_75t_L g654 ( .A(n_453), .B(n_618), .Y(n_654) );
AND2x2_ASAP7_75t_L g683 ( .A(n_453), .B(n_593), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_453), .B(n_565), .Y(n_700) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g580 ( .A(n_454), .B(n_475), .Y(n_580) );
BUFx3_ASAP7_75t_L g605 ( .A(n_454), .Y(n_605) );
AND2x2_ASAP7_75t_L g634 ( .A(n_454), .B(n_476), .Y(n_634) );
AND3x2_ASAP7_75t_L g647 ( .A(n_454), .B(n_648), .C(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g570 ( .A(n_464), .Y(n_570) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AOI32xp33_ASAP7_75t_L g625 ( .A1(n_465), .A2(n_577), .A3(n_626), .B1(n_629), .B2(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g552 ( .A(n_466), .B(n_475), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_466), .B(n_580), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_466), .B(n_602), .Y(n_630) );
OR2x2_ASAP7_75t_L g636 ( .A(n_466), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_466), .B(n_591), .Y(n_661) );
OR2x2_ASAP7_75t_L g679 ( .A(n_466), .B(n_504), .Y(n_679) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g543 ( .A(n_467), .B(n_485), .Y(n_543) );
INVx2_ASAP7_75t_L g565 ( .A(n_467), .Y(n_565) );
OR2x2_ASAP7_75t_L g587 ( .A(n_467), .B(n_485), .Y(n_587) );
AND2x2_ASAP7_75t_L g592 ( .A(n_467), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_467), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_467), .B(n_542), .Y(n_648) );
INVx1_ASAP7_75t_SL g699 ( .A(n_475), .Y(n_699) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
INVx1_ASAP7_75t_SL g542 ( .A(n_476), .Y(n_542) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_476), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_476), .B(n_628), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_476), .B(n_565), .C(n_683), .Y(n_694) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_477), .A2(n_486), .B(n_492), .Y(n_485) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_477), .A2(n_496), .B(n_502), .Y(n_495) );
INVx2_ASAP7_75t_L g593 ( .A(n_485), .Y(n_593) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_485), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
INVx1_ASAP7_75t_L g629 ( .A(n_494), .Y(n_629) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g547 ( .A(n_495), .B(n_529), .Y(n_547) );
INVx2_ASAP7_75t_L g564 ( .A(n_495), .Y(n_564) );
AND2x2_ASAP7_75t_L g569 ( .A(n_495), .B(n_530), .Y(n_569) );
AND2x2_ASAP7_75t_L g584 ( .A(n_495), .B(n_517), .Y(n_584) );
AND2x2_ASAP7_75t_L g596 ( .A(n_495), .B(n_568), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_503), .B(n_612), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_503), .B(n_569), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_503), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_503), .B(n_563), .Y(n_691) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g528 ( .A(n_504), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_504), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g573 ( .A(n_504), .B(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g599 ( .A(n_504), .B(n_529), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_504), .B(n_639), .Y(n_638) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_514), .Y(n_504) );
INVx1_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_510), .B(n_513), .Y(n_509) );
INVx2_ASAP7_75t_L g524 ( .A(n_513), .Y(n_524) );
INVx1_ASAP7_75t_L g559 ( .A(n_514), .Y(n_559) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_517), .B(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g563 ( .A(n_517), .B(n_564), .Y(n_563) );
INVx3_ASAP7_75t_SL g568 ( .A(n_517), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_517), .B(n_555), .Y(n_621) );
OR2x2_ASAP7_75t_L g631 ( .A(n_517), .B(n_557), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_517), .B(n_599), .Y(n_659) );
OR2x2_ASAP7_75t_L g689 ( .A(n_517), .B(n_529), .Y(n_689) );
AND2x2_ASAP7_75t_L g693 ( .A(n_517), .B(n_530), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_517), .B(n_569), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_517), .B(n_595), .Y(n_713) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_526), .Y(n_517) );
INVx1_ASAP7_75t_SL g656 ( .A(n_528), .Y(n_656) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_557), .Y(n_595) );
AND2x2_ASAP7_75t_L g609 ( .A(n_529), .B(n_564), .Y(n_609) );
AND2x2_ASAP7_75t_L g612 ( .A(n_529), .B(n_568), .Y(n_612) );
INVx1_ASAP7_75t_L g639 ( .A(n_529), .Y(n_639) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g551 ( .A(n_530), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_541), .A2(n_587), .B(n_711), .C(n_712), .Y(n_710) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_543), .B(n_560), .Y(n_575) );
AND2x2_ASAP7_75t_L g601 ( .A(n_543), .B(n_602), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_545), .A2(n_548), .B(n_552), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_546), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g572 ( .A(n_547), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_547), .B(n_568), .Y(n_613) );
AND2x2_ASAP7_75t_L g704 ( .A(n_547), .B(n_555), .Y(n_704) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g577 ( .A(n_551), .B(n_564), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_551), .B(n_562), .Y(n_578) );
OAI322xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_561), .A3(n_562), .B1(n_565), .B2(n_566), .C1(n_570), .C2(n_571), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
AND2x2_ASAP7_75t_L g665 ( .A(n_555), .B(n_577), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_555), .B(n_629), .Y(n_711) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g608 ( .A(n_557), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g674 ( .A(n_561), .B(n_587), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_562), .B(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_563), .B(n_595), .Y(n_652) );
AND2x2_ASAP7_75t_L g598 ( .A(n_564), .B(n_568), .Y(n_598) );
AND2x2_ASAP7_75t_L g606 ( .A(n_565), .B(n_607), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_565), .A2(n_644), .B(n_704), .C(n_705), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_566), .A2(n_579), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_568), .B(n_595), .Y(n_635) );
AND2x2_ASAP7_75t_L g641 ( .A(n_568), .B(n_609), .Y(n_641) );
AND2x2_ASAP7_75t_L g675 ( .A(n_568), .B(n_577), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_569), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_SL g685 ( .A(n_569), .Y(n_685) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_573), .A2(n_601), .B1(n_603), .B2(n_608), .Y(n_600) );
OAI22xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_576), .B1(n_578), .B2(n_579), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_575), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_610) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_580), .A2(n_682), .B1(n_684), .B2(n_686), .C(n_690), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_589), .C(n_610), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g651 ( .A(n_587), .B(n_604), .Y(n_651) );
INVx1_ASAP7_75t_L g702 ( .A(n_587), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_588), .A2(n_590), .B1(n_594), .B2(n_597), .C(n_600), .Y(n_589) );
INVx2_ASAP7_75t_SL g644 ( .A(n_588), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
AND2x2_ASAP7_75t_L g633 ( .A(n_592), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g618 ( .A(n_593), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g680 ( .A(n_596), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_604), .B(n_706), .Y(n_705) );
CKINVDCx16_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g649 ( .A(n_607), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_608), .A2(n_620), .B(n_622), .C(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g697 ( .A(n_611), .Y(n_697) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_615), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g628 ( .A(n_618), .Y(n_628) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI222xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_631), .B1(n_632), .B2(n_635), .C1(n_636), .C2(n_638), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g664 ( .A(n_628), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_631), .B(n_685), .Y(n_684) );
NAND2xp33_ASAP7_75t_SL g662 ( .A(n_632), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g637 ( .A(n_634), .Y(n_637) );
AND2x2_ASAP7_75t_L g701 ( .A(n_634), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g667 ( .A(n_637), .B(n_664), .Y(n_667) );
INVx1_ASAP7_75t_L g696 ( .A(n_638), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_645), .C(n_650), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_644), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_647), .A2(n_675), .A3(n_680), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_701), .Y(n_695) );
AND2x2_ASAP7_75t_L g682 ( .A(n_648), .B(n_683), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_655), .Y(n_650) );
INVxp33_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_662), .B2(n_665), .C(n_666), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND5xp2_ASAP7_75t_L g669 ( .A(n_670), .B(n_681), .C(n_695), .D(n_703), .E(n_707), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B(n_676), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVxp33_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_683), .A2(n_708), .B(n_709), .C(n_710), .Y(n_707) );
AOI31xp33_ASAP7_75t_L g690 ( .A1(n_685), .A2(n_691), .A3(n_692), .B(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g708 ( .A(n_706), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g721 ( .A(n_714), .Y(n_721) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_736), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
endmodule