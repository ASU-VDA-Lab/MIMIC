module fake_jpeg_27920_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_31),
.B1(n_33),
.B2(n_32),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_31),
.B1(n_20),
.B2(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_48),
.B1(n_56),
.B2(n_58),
.Y(n_83)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_33),
.B1(n_32),
.B2(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_67),
.Y(n_68)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_33),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_29),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_29),
.B1(n_30),
.B2(n_19),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_41),
.B1(n_42),
.B2(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_84),
.B1(n_56),
.B2(n_60),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_42),
.B1(n_35),
.B2(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_64),
.B1(n_58),
.B2(n_45),
.Y(n_95)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_17),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_29),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_87),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_38),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_102),
.B1(n_111),
.B2(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_98),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_103),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_66),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_114),
.C(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_113),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_67),
.B(n_50),
.C(n_47),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_51),
.B(n_47),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_65),
.B1(n_53),
.B2(n_19),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_66),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_65),
.B1(n_53),
.B2(n_50),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_92),
.Y(n_125)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_83),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_91),
.B1(n_83),
.B2(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_126),
.B1(n_137),
.B2(n_109),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_30),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_80),
.B1(n_81),
.B2(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_135),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_81),
.B1(n_74),
.B2(n_76),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_74),
.B1(n_73),
.B2(n_51),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_52),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_140),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_52),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_86),
.B(n_106),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_52),
.C(n_89),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_110),
.C(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_116),
.B(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_151),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_158),
.B1(n_133),
.B2(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_124),
.B1(n_121),
.B2(n_137),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_129),
.B1(n_138),
.B2(n_143),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_156),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_165),
.C(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_97),
.B1(n_116),
.B2(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_167),
.B1(n_168),
.B2(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_163),
.B(n_164),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_112),
.B(n_98),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_138),
.C(n_141),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_106),
.C(n_117),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_94),
.B1(n_106),
.B2(n_30),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_192),
.B1(n_167),
.B2(n_168),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_150),
.B1(n_152),
.B2(n_156),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_174),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_173),
.B(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_135),
.C(n_125),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_183),
.C(n_186),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_160),
.B(n_155),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_128),
.C(n_123),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_123),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_38),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_144),
.C(n_130),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_144),
.B(n_130),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_163),
.B(n_159),
.Y(n_207)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_21),
.A3(n_23),
.B1(n_8),
.B2(n_15),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_148),
.A2(n_21),
.B1(n_38),
.B2(n_23),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_205),
.B1(n_209),
.B2(n_192),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_176),
.B(n_154),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_206),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_150),
.B1(n_153),
.B2(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_23),
.B(n_2),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_181),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_154),
.C(n_146),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_215),
.C(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_145),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_200),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_21),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_187),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_170),
.B1(n_190),
.B2(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_215),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_185),
.C(n_191),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_212),
.C(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_0),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_202),
.B(n_196),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_1),
.B(n_2),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_239),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

OAI322xp33_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_207),
.A3(n_210),
.B1(n_9),
.B2(n_10),
.C1(n_5),
.C2(n_6),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_244),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_210),
.A3(n_21),
.B1(n_8),
.B2(n_10),
.C1(n_5),
.C2(n_6),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_7),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_227),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_225),
.C(n_221),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_220),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_216),
.C(n_232),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_216),
.C(n_235),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_224),
.B(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_217),
.C(n_231),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_237),
.B1(n_243),
.B2(n_251),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_264),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_226),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_237),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_267),
.C(n_252),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_228),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_233),
.B(n_250),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_242),
.B1(n_220),
.B2(n_222),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_270),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_275),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_274),
.B(n_276),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_265),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_238),
.C(n_9),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_5),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_261),
.B(n_9),
.Y(n_284)
);

NOR2x1_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_266),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_285),
.B(n_12),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_284),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_11),
.B(n_12),
.C(n_15),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_11),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.C(n_285),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_282),
.C(n_2),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_15),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_291),
.B1(n_286),
.B2(n_3),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_4),
.B(n_1),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_1),
.Y(n_295)
);


endmodule