module fake_jpeg_15625_n_365 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_365);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_365;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_45),
.B(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_61),
.Y(n_103)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_59),
.Y(n_95)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_75),
.B(n_77),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_26),
.B1(n_37),
.B2(n_36),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_79),
.A2(n_98),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_42),
.B(n_20),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_90),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_24),
.B1(n_28),
.B2(n_20),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_33),
.B1(n_23),
.B2(n_34),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_41),
.A2(n_35),
.B1(n_32),
.B2(n_28),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_35),
.B1(n_24),
.B2(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_105),
.Y(n_149)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_49),
.A2(n_23),
.B(n_22),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_48),
.B(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_17),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_119),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_117),
.A2(n_144),
.B1(n_158),
.B2(n_138),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_30),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_30),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_123),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_12),
.B1(n_11),
.B2(n_23),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_132),
.B1(n_92),
.B2(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_30),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_12),
.B(n_25),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_R g170 ( 
.A(n_124),
.B(n_134),
.Y(n_170)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_34),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_142),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_25),
.B1(n_34),
.B2(n_2),
.Y(n_132)
);

OR2x2_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_25),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_70),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_83),
.B(n_0),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_145),
.Y(n_176)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_1),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_5),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_146),
.B(n_150),
.Y(n_192)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_4),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_82),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_72),
.B(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_154),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_85),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_79),
.B(n_10),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_5),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_146),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_102),
.B1(n_99),
.B2(n_72),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_167),
.A2(n_145),
.B1(n_139),
.B2(n_135),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_114),
.B(n_69),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_139),
.C(n_117),
.Y(n_207)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_178),
.A2(n_186),
.B(n_193),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_118),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_112),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_201),
.Y(n_216)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_65),
.B(n_71),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_127),
.A2(n_86),
.B1(n_78),
.B2(n_109),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_188),
.A2(n_198),
.B1(n_128),
.B2(n_129),
.Y(n_230)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_190),
.Y(n_226)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_5),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_199),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_202),
.B1(n_149),
.B2(n_137),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_123),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_148),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_131),
.B(n_143),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_142),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_220),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_181),
.B(n_168),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_235),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_231),
.B1(n_180),
.B2(n_187),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_147),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_210),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_147),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_214),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_143),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_219),
.B1(n_230),
.B2(n_235),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_136),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_145),
.B1(n_120),
.B2(n_118),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_130),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_229),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_140),
.C(n_116),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_165),
.C(n_187),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_227),
.B(n_233),
.Y(n_266)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

AO21x2_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_128),
.B(n_141),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_232),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_164),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_156),
.B1(n_7),
.B2(n_10),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_179),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_176),
.A2(n_10),
.B1(n_178),
.B2(n_186),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_166),
.A2(n_172),
.B1(n_170),
.B2(n_202),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_170),
.A2(n_198),
.B1(n_176),
.B2(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_163),
.B(n_175),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_249),
.C(n_251),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_161),
.B1(n_194),
.B2(n_189),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_244),
.A2(n_261),
.B(n_263),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_246),
.B(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_247),
.A2(n_248),
.B1(n_264),
.B2(n_269),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_195),
.B1(n_185),
.B2(n_168),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_220),
.C(n_238),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_191),
.C(n_169),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_169),
.C(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_236),
.C(n_219),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_215),
.B(n_234),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_SL g262 ( 
.A(n_231),
.B(n_216),
.C(n_237),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_250),
.B(n_246),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_206),
.A2(n_231),
.B(n_230),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_206),
.B1(n_229),
.B2(n_205),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_203),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_213),
.C(n_221),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_223),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_284),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_247),
.B1(n_264),
.B2(n_244),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_277),
.A2(n_279),
.B1(n_287),
.B2(n_289),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_260),
.B1(n_257),
.B2(n_262),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_223),
.B(n_228),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_203),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_268),
.B(n_248),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_294),
.B1(n_281),
.B2(n_277),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_245),
.A2(n_249),
.B1(n_265),
.B2(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_297),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_241),
.A2(n_259),
.B1(n_270),
.B2(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_264),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_204),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_258),
.B(n_255),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_300),
.A2(n_307),
.B1(n_306),
.B2(n_312),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_293),
.C(n_275),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_315),
.C(n_287),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_295),
.B1(n_278),
.B2(n_273),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_304),
.B1(n_300),
.B2(n_315),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_316),
.Y(n_324)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_286),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_285),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_292),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_278),
.C(n_289),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_280),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_327),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_311),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_320),
.B(n_322),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_325),
.C(n_332),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_328),
.Y(n_343)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_326),
.A2(n_331),
.B(n_335),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_284),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_291),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_274),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_312),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_306),
.B(n_274),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_330),
.B(n_334),
.Y(n_339)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_297),
.C(n_281),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_298),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_304),
.A2(n_280),
.B(n_283),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_333),
.B(n_308),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_341),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_301),
.B(n_305),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_345),
.C(n_339),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_317),
.C(n_305),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_324),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_347),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_318),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_340),
.C(n_337),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_339),
.A2(n_328),
.B(n_322),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_338),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_350),
.B(n_340),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_354),
.Y(n_356)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_353),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_356),
.A2(n_354),
.B(n_345),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_358),
.B(n_355),
.C(n_332),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_360),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_361),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_359),
.B(n_355),
.C(n_347),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_363),
.A2(n_331),
.B1(n_318),
.B2(n_326),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_342),
.Y(n_365)
);


endmodule