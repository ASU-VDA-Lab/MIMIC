module fake_jpeg_16431_n_355 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_355);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_37),
.B1(n_31),
.B2(n_26),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_69),
.B1(n_82),
.B2(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_20),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_37),
.B1(n_26),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_37),
.B1(n_26),
.B2(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_77),
.B1(n_23),
.B2(n_38),
.Y(n_101)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_21),
.B1(n_30),
.B2(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_40),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_33),
.Y(n_85)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_90),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_93),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_79),
.Y(n_93)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_108),
.B1(n_21),
.B2(n_70),
.Y(n_140)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_107),
.B1(n_112),
.B2(n_64),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_40),
.B1(n_35),
.B2(n_39),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_64),
.B1(n_77),
.B2(n_55),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_39),
.B1(n_29),
.B2(n_76),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_126),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_77),
.B(n_69),
.C(n_60),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_118),
.A2(n_127),
.B(n_36),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_131),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_146),
.B1(n_102),
.B2(n_97),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_42),
.C(n_46),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_111),
.C(n_94),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_94),
.C(n_53),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_68),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_68),
.B1(n_101),
.B2(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_144),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_82),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_62),
.C(n_66),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_29),
.B(n_77),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_110),
.B(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_21),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_141),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_140),
.A2(n_148),
.B1(n_116),
.B2(n_96),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_27),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_61),
.B1(n_30),
.B2(n_36),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_57),
.B1(n_61),
.B2(n_30),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_173),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_93),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_158),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_160),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_127),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_165),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_136),
.B1(n_142),
.B2(n_141),
.Y(n_176)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_145),
.B(n_131),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_27),
.B(n_1),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_176),
.A2(n_178),
.B1(n_186),
.B2(n_192),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_197),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_124),
.B1(n_118),
.B2(n_125),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_117),
.B1(n_130),
.B2(n_126),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_135),
.CI(n_121),
.CON(n_185),
.SN(n_185)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_189),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_161),
.B1(n_169),
.B2(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_136),
.B(n_123),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_133),
.B(n_144),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_165),
.B1(n_164),
.B2(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_172),
.B1(n_151),
.B2(n_150),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_159),
.B1(n_154),
.B2(n_152),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_148),
.Y(n_192)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_145),
.A3(n_147),
.B1(n_115),
.B2(n_134),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_168),
.Y(n_213)
);

AND2x4_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_147),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_170),
.C(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_203),
.C(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_202),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_166),
.C(n_155),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_158),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_206),
.A2(n_213),
.B(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_208),
.B(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_163),
.Y(n_211)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_188),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_168),
.Y(n_216)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_219),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_63),
.C(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_182),
.B(n_27),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_182),
.B(n_27),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_100),
.C(n_103),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_223),
.C(n_224),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_147),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_100),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_210),
.B1(n_178),
.B2(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_227),
.A2(n_244),
.B1(n_0),
.B2(n_1),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_174),
.B1(n_197),
.B2(n_190),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_234),
.B1(n_198),
.B2(n_214),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_231),
.B(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_197),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_176),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_241),
.A2(n_242),
.B1(n_215),
.B2(n_217),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_174),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_174),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_192),
.C(n_194),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_27),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_184),
.B(n_134),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_220),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_0),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_251),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_262),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_198),
.B1(n_218),
.B2(n_222),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_260),
.B1(n_269),
.B2(n_237),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_209),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_103),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_230),
.A2(n_36),
.B1(n_30),
.B2(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_228),
.C(n_246),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_284),
.C(n_288),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_228),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_235),
.C(n_243),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_286),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_225),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_289),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_245),
.C(n_248),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_252),
.B1(n_271),
.B2(n_241),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_303),
.B1(n_305),
.B2(n_242),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_300),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_253),
.B(n_255),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_297),
.A2(n_299),
.B(n_242),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_234),
.B(n_252),
.C(n_231),
.D(n_264),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_298),
.A2(n_301),
.B1(n_247),
.B2(n_276),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_233),
.B(n_268),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_272),
.A2(n_281),
.B1(n_273),
.B2(n_236),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_277),
.B(n_238),
.CI(n_230),
.CON(n_302),
.SN(n_302)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_232),
.B(n_247),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_254),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_313),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_267),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_315),
.C(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_284),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_285),
.C(n_274),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_320),
.C(n_319),
.Y(n_331)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_275),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_299),
.B(n_291),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_275),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_265),
.C(n_3),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_330),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_324),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_300),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_325),
.A2(n_11),
.B(n_16),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_305),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_297),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_318),
.B(n_295),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_302),
.C(n_3),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_333),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_303),
.B1(n_302),
.B2(n_5),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_340),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_12),
.B1(n_17),
.B2(n_6),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_337),
.Y(n_341)
);

AOI31xp67_ASAP7_75t_L g338 ( 
.A1(n_325),
.A2(n_11),
.A3(n_16),
.B(n_6),
.Y(n_338)
);

AOI21x1_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_10),
.B(n_15),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_12),
.C(n_16),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_326),
.B1(n_12),
.B2(n_6),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_343),
.C(n_13),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_10),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_344),
.A2(n_7),
.B(n_10),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_L g347 ( 
.A1(n_345),
.A2(n_337),
.B(n_334),
.C(n_7),
.D(n_9),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_348),
.A3(n_349),
.B1(n_346),
.B2(n_345),
.C1(n_341),
.C2(n_14),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_18),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_353),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_355)
);


endmodule