module fake_jpeg_1717_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_0),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_21),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_6),
.Y(n_22)
);

CKINVDCx12_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_8),
.C(n_11),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_18),
.B(n_10),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_27),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_20),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_29),
.C(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_37),
.CI(n_14),
.CON(n_39),
.SN(n_39)
);

AO22x1_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_33),
.B1(n_19),
.B2(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_19),
.C(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_16),
.B1(n_14),
.B2(n_1),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_40),
.B(n_39),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_41),
.C(n_39),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_38),
.B(n_6),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_38),
.Y(n_46)
);


endmodule