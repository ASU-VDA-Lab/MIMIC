module fake_jpeg_24794_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_17),
.Y(n_22)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_16),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_10),
.C(n_12),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_27),
.C(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_26),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_9),
.B(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_15),
.B1(n_19),
.B2(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_32),
.B1(n_0),
.B2(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_22),
.A2(n_15),
.B1(n_20),
.B2(n_18),
.Y(n_32)
);

XNOR2x1_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_36),
.C(n_35),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_29),
.B1(n_2),
.B2(n_1),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_11),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.C(n_29),
.Y(n_39)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_33),
.B(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AOI221xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_2),
.B1(n_4),
.B2(n_41),
.C(n_43),
.Y(n_45)
);


endmodule