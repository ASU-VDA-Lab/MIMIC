module fake_jpeg_3233_n_225 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_225);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_52),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_92),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_65),
.B(n_72),
.C(n_74),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_66),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_84),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_53),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_115),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_82),
.B1(n_78),
.B2(n_63),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_112),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_63),
.B1(n_55),
.B2(n_73),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_76),
.B1(n_59),
.B2(n_71),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_79),
.B1(n_59),
.B2(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_129),
.B1(n_132),
.B2(n_110),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_110),
.Y(n_144)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_130),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_76),
.B(n_60),
.C(n_67),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_102),
.B(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_69),
.B1(n_60),
.B2(n_67),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_33),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_23),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_155),
.B1(n_134),
.B2(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_149),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.C(n_153),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_60),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_1),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_1),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_64),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_2),
.Y(n_154)
);

NOR4xp25_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_54),
.B1(n_64),
.B2(n_4),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_64),
.B(n_54),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_40),
.B(n_39),
.C(n_38),
.D(n_37),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_126),
.B1(n_124),
.B2(n_121),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_162),
.B(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_49),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_179),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_48),
.B1(n_47),
.B2(n_44),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_175),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_140),
.B1(n_36),
.B2(n_35),
.C(n_34),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_8),
.B(n_9),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_183),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_30),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_187),
.Y(n_200)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_171),
.B1(n_160),
.B2(n_175),
.C(n_165),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_26),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_25),
.C(n_15),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_18),
.Y(n_203)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

AO221x1_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_178),
.B1(n_163),
.B2(n_168),
.C(n_17),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_198),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_14),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_203),
.C(n_193),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_191),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_190),
.B1(n_182),
.B2(n_187),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_16),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_205),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_18),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_212),
.C(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_190),
.B(n_186),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_19),
.B(n_20),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_186),
.C(n_183),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_216),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_204),
.C(n_203),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_208),
.C(n_20),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_21),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_208),
.C(n_218),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_21),
.Y(n_225)
);


endmodule