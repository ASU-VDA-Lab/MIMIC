module real_aes_9057_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_1), .A2(n_142), .B(n_146), .C(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g195 ( .A(n_2), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_3), .A2(n_137), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_4), .B(n_159), .Y(n_476) );
AOI21xp33_ASAP7_75t_L g163 ( .A1(n_5), .A2(n_137), .B(n_164), .Y(n_163) );
AND2x6_ASAP7_75t_L g142 ( .A(n_6), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_7), .A2(n_245), .B(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_40), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_8), .B(n_40), .Y(n_734) );
INVx1_ASAP7_75t_L g532 ( .A(n_9), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_10), .B(n_168), .Y(n_511) );
INVx1_ASAP7_75t_L g170 ( .A(n_11), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_12), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
INVx1_ASAP7_75t_L g251 ( .A(n_14), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_15), .A2(n_154), .B(n_252), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_16), .B(n_159), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_17), .B(n_151), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_18), .B(n_137), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_19), .B(n_560), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_20), .A2(n_178), .B(n_237), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_21), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_22), .B(n_168), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_23), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_24), .B(n_168), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_25), .Y(n_456) );
INVx1_ASAP7_75t_L g482 ( .A(n_26), .Y(n_482) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_27), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_28), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_29), .B(n_168), .Y(n_197) );
INVx1_ASAP7_75t_L g557 ( .A(n_30), .Y(n_557) );
INVx1_ASAP7_75t_L g184 ( .A(n_31), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_32), .A2(n_92), .B1(n_751), .B2(n_752), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_32), .Y(n_752) );
INVx2_ASAP7_75t_L g140 ( .A(n_33), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_34), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_35), .A2(n_155), .B(n_237), .C(n_474), .Y(n_473) );
INVxp67_ASAP7_75t_L g558 ( .A(n_36), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_37), .A2(n_142), .B(n_146), .C(n_209), .Y(n_208) );
CKINVDCx14_ASAP7_75t_R g472 ( .A(n_38), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_39), .A2(n_146), .B(n_481), .C(n_486), .Y(n_480) );
INVx1_ASAP7_75t_L g182 ( .A(n_41), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_42), .A2(n_49), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_42), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_43), .A2(n_63), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_43), .Y(n_730) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_44), .A2(n_727), .B1(n_728), .B2(n_731), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_44), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_45), .A2(n_167), .B(n_213), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_46), .B(n_168), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_47), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_48), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_49), .Y(n_747) );
INVx1_ASAP7_75t_L g497 ( .A(n_50), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_51), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_52), .B(n_137), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_53), .A2(n_146), .B1(n_178), .B2(n_180), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_54), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_55), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_56), .A2(n_155), .B(n_167), .C(n_169), .Y(n_166) );
CKINVDCx14_ASAP7_75t_R g529 ( .A(n_57), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_58), .Y(n_227) );
INVx1_ASAP7_75t_L g165 ( .A(n_59), .Y(n_165) );
INVx1_ASAP7_75t_L g143 ( .A(n_60), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_61), .Y(n_738) );
INVx1_ASAP7_75t_L g134 ( .A(n_62), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_63), .Y(n_729) );
INVx1_ASAP7_75t_SL g475 ( .A(n_64), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_65), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_66), .B(n_159), .Y(n_501) );
INVx1_ASAP7_75t_L g459 ( .A(n_67), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_68), .A2(n_105), .B1(n_113), .B2(n_763), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_69), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_SL g150 ( .A1(n_70), .A2(n_151), .B(n_152), .C(n_155), .Y(n_150) );
INVxp67_ASAP7_75t_L g153 ( .A(n_71), .Y(n_153) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_73), .A2(n_137), .B(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_74), .A2(n_725), .B1(n_726), .B2(n_732), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_74), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_75), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_76), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_77), .A2(n_137), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g220 ( .A(n_78), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_79), .A2(n_245), .B(n_553), .Y(n_552) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_80), .Y(n_479) );
INVx1_ASAP7_75t_L g517 ( .A(n_81), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_82), .A2(n_142), .B(n_146), .C(n_222), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_83), .A2(n_137), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g520 ( .A(n_84), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_85), .B(n_196), .Y(n_210) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g510 ( .A(n_87), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_88), .B(n_151), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_89), .A2(n_142), .B(n_146), .C(n_194), .Y(n_193) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_90), .B(n_109), .C(n_110), .Y(n_108) );
INVx2_ASAP7_75t_L g119 ( .A(n_90), .Y(n_119) );
OR2x2_ASAP7_75t_L g758 ( .A(n_90), .B(n_737), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_91), .A2(n_146), .B(n_458), .C(n_462), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_92), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_92), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_93), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_94), .A2(n_142), .B(n_146), .C(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_95), .Y(n_241) );
INVx1_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_97), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_98), .B(n_196), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_99), .B(n_130), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_100), .B(n_130), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_101), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_102), .A2(n_137), .B(n_144), .Y(n_136) );
INVx2_ASAP7_75t_L g500 ( .A(n_103), .Y(n_500) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g764 ( .A(n_106), .Y(n_764) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g733 ( .A(n_109), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO221x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_739), .B1(n_744), .B2(n_754), .C(n_759), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_733), .B1(n_735), .B2(n_738), .Y(n_114) );
XOR2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_724), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B1(n_446), .B2(n_447), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g446 ( .A(n_119), .Y(n_446) );
NOR2x2_ASAP7_75t_L g736 ( .A(n_119), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND4x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_364), .C(n_411), .D(n_431), .Y(n_122) );
NOR3xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_294), .C(n_319), .Y(n_123) );
OAI211xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_202), .B(n_254), .C(n_284), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_173), .Y(n_126) );
INVx3_ASAP7_75t_SL g336 ( .A(n_127), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_127), .B(n_267), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_127), .B(n_189), .Y(n_417) );
AND2x2_ASAP7_75t_L g440 ( .A(n_127), .B(n_306), .Y(n_440) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_161), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g258 ( .A(n_129), .B(n_162), .Y(n_258) );
INVx3_ASAP7_75t_L g271 ( .A(n_129), .Y(n_271) );
AND2x2_ASAP7_75t_L g276 ( .A(n_129), .B(n_161), .Y(n_276) );
OR2x2_ASAP7_75t_L g327 ( .A(n_129), .B(n_268), .Y(n_327) );
BUFx2_ASAP7_75t_L g347 ( .A(n_129), .Y(n_347) );
AND2x2_ASAP7_75t_L g357 ( .A(n_129), .B(n_268), .Y(n_357) );
AND2x2_ASAP7_75t_L g363 ( .A(n_129), .B(n_174), .Y(n_363) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_136), .B(n_158), .Y(n_129) );
INVx4_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_130), .Y(n_469) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_132), .B(n_133), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx2_ASAP7_75t_L g245 ( .A(n_137), .Y(n_245) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_138), .B(n_142), .Y(n_186) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g485 ( .A(n_139), .Y(n_485) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g179 ( .A(n_140), .Y(n_179) );
INVx1_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
INVx1_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
INVx3_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_141), .Y(n_181) );
INVx4_ASAP7_75t_SL g157 ( .A(n_142), .Y(n_157) );
BUFx3_ASAP7_75t_L g486 ( .A(n_142), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B(n_150), .C(n_157), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_145), .A2(n_157), .B(n_165), .C(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_145), .A2(n_157), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_145), .A2(n_157), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_145), .A2(n_157), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_145), .A2(n_157), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_145), .A2(n_157), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_145), .A2(n_157), .B(n_554), .C(n_555), .Y(n_553) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
BUFx3_ASAP7_75t_L g214 ( .A(n_147), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_154), .B(n_170), .Y(n_169) );
INVx5_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_154), .B(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_156), .Y(n_238) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_157), .A2(n_177), .B1(n_185), .B2(n_186), .Y(n_176) );
INVx1_ASAP7_75t_L g462 ( .A(n_157), .Y(n_462) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_159), .A2(n_163), .B(n_171), .Y(n_162) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_160), .B(n_217), .Y(n_216) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_160), .A2(n_455), .B(n_463), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_160), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_160), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_162), .B(n_268), .Y(n_282) );
INVx2_ASAP7_75t_L g292 ( .A(n_162), .Y(n_292) );
AND2x2_ASAP7_75t_L g305 ( .A(n_162), .B(n_271), .Y(n_305) );
OR2x2_ASAP7_75t_L g316 ( .A(n_162), .B(n_268), .Y(n_316) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_162), .B(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g374 ( .A(n_162), .Y(n_374) );
AND2x2_ASAP7_75t_L g420 ( .A(n_162), .B(n_174), .Y(n_420) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
INVx1_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
INVx2_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_172), .A2(n_244), .B(n_253), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_172), .A2(n_186), .B(n_479), .C(n_480), .Y(n_478) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_172), .A2(n_527), .B(n_533), .Y(n_526) );
INVx3_ASAP7_75t_SL g293 ( .A(n_173), .Y(n_293) );
OR2x2_ASAP7_75t_L g346 ( .A(n_173), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_189), .Y(n_173) );
INVx3_ASAP7_75t_L g268 ( .A(n_174), .Y(n_268) );
AND2x2_ASAP7_75t_L g335 ( .A(n_174), .B(n_190), .Y(n_335) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_174), .Y(n_403) );
AOI33xp33_ASAP7_75t_L g407 ( .A1(n_174), .A2(n_336), .A3(n_343), .B1(n_352), .B2(n_408), .B3(n_409), .Y(n_407) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_187), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_175), .B(n_188), .Y(n_187) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_175), .A2(n_191), .B(n_199), .Y(n_190) );
INVx2_ASAP7_75t_L g215 ( .A(n_175), .Y(n_215) );
INVx2_ASAP7_75t_L g198 ( .A(n_178), .Y(n_198) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_180) );
INVx2_ASAP7_75t_L g183 ( .A(n_181), .Y(n_183) );
INVx4_ASAP7_75t_L g249 ( .A(n_181), .Y(n_249) );
INVx2_ASAP7_75t_L g460 ( .A(n_183), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_220), .B(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_186), .A2(n_456), .B(n_457), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_186), .A2(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g256 ( .A(n_189), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_189), .B(n_271), .Y(n_270) );
NOR3xp33_ASAP7_75t_L g330 ( .A(n_189), .B(n_331), .C(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g356 ( .A(n_189), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_189), .B(n_363), .Y(n_366) );
AND2x2_ASAP7_75t_L g419 ( .A(n_189), .B(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g275 ( .A(n_190), .Y(n_275) );
OR2x2_ASAP7_75t_L g369 ( .A(n_190), .B(n_268), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .C(n_198), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_196), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_196), .A2(n_249), .B1(n_557), .B2(n_558), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_201), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_201), .B(n_241), .Y(n_240) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_201), .A2(n_506), .B(n_512), .Y(n_505) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_228), .Y(n_202) );
AOI32xp33_ASAP7_75t_L g320 ( .A1(n_203), .A2(n_321), .A3(n_323), .B1(n_325), .B2(n_328), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_203), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g423 ( .A(n_203), .Y(n_423) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g355 ( .A(n_204), .B(n_339), .Y(n_355) );
AND2x2_ASAP7_75t_L g375 ( .A(n_204), .B(n_301), .Y(n_375) );
AND2x2_ASAP7_75t_L g443 ( .A(n_204), .B(n_361), .Y(n_443) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_218), .Y(n_204) );
INVx3_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
AND2x2_ASAP7_75t_L g278 ( .A(n_205), .B(n_262), .Y(n_278) );
OR2x2_ASAP7_75t_L g283 ( .A(n_205), .B(n_261), .Y(n_283) );
INVx1_ASAP7_75t_L g290 ( .A(n_205), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_205), .B(n_272), .Y(n_298) );
AND2x2_ASAP7_75t_L g300 ( .A(n_205), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_205), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g353 ( .A(n_205), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_205), .B(n_438), .Y(n_437) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
AOI21xp5_ASAP7_75t_SL g206 ( .A1(n_207), .A2(n_208), .B(n_215), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_212), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_212), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
O2A1O1Ixp5_ASAP7_75t_L g509 ( .A1(n_212), .A2(n_460), .B(n_510), .C(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
INVx1_ASAP7_75t_L g225 ( .A(n_215), .Y(n_225) );
INVx2_ASAP7_75t_L g262 ( .A(n_218), .Y(n_262) );
AND2x2_ASAP7_75t_L g308 ( .A(n_218), .B(n_229), .Y(n_308) );
AND2x2_ASAP7_75t_L g318 ( .A(n_218), .B(n_243), .Y(n_318) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_225), .B(n_226), .Y(n_218) );
INVx1_ASAP7_75t_L g551 ( .A(n_225), .Y(n_551) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_225), .A2(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g438 ( .A(n_228), .Y(n_438) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_242), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_229), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
AND2x2_ASAP7_75t_L g323 ( .A(n_229), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g339 ( .A(n_229), .B(n_302), .Y(n_339) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g287 ( .A(n_230), .Y(n_287) );
AND2x2_ASAP7_75t_L g301 ( .A(n_230), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g352 ( .A(n_230), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_230), .B(n_262), .Y(n_384) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_240), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_231), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g560 ( .A(n_231), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_238), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_237), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g263 ( .A(n_242), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g324 ( .A(n_242), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_242), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g361 ( .A(n_242), .Y(n_361) );
INVx1_ASAP7_75t_L g394 ( .A(n_242), .Y(n_394) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g272 ( .A(n_243), .B(n_262), .Y(n_272) );
INVx1_ASAP7_75t_L g302 ( .A(n_243), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_249), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_249), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_249), .B(n_520), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B1(n_265), .B2(n_272), .C(n_273), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_256), .B(n_276), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_256), .B(n_339), .Y(n_416) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_258), .B(n_306), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_258), .B(n_267), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_258), .B(n_281), .Y(n_410) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g332 ( .A(n_262), .Y(n_332) );
AND2x2_ASAP7_75t_L g307 ( .A(n_263), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
AND2x2_ASAP7_75t_L g317 ( .A(n_264), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_264), .B(n_287), .Y(n_333) );
AND2x2_ASAP7_75t_L g397 ( .A(n_264), .B(n_323), .Y(n_397) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g306 ( .A(n_268), .B(n_275), .Y(n_306) );
AND2x2_ASAP7_75t_L g402 ( .A(n_269), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_271), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_272), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_272), .B(n_279), .Y(n_367) );
AND2x2_ASAP7_75t_L g387 ( .A(n_272), .B(n_287), .Y(n_387) );
AND2x2_ASAP7_75t_L g408 ( .A(n_272), .B(n_352), .Y(n_408) );
OAI32xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .A3(n_279), .B1(n_280), .B2(n_283), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_SL g281 ( .A(n_275), .Y(n_281) );
NAND2x1_ASAP7_75t_L g322 ( .A(n_275), .B(n_305), .Y(n_322) );
OR2x2_ASAP7_75t_L g326 ( .A(n_275), .B(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_275), .B(n_374), .Y(n_427) );
INVx1_ASAP7_75t_L g295 ( .A(n_276), .Y(n_295) );
OAI221xp5_ASAP7_75t_SL g413 ( .A1(n_277), .A2(n_368), .B1(n_414), .B2(n_417), .C(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g285 ( .A(n_278), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g328 ( .A(n_278), .B(n_301), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_278), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g406 ( .A(n_278), .B(n_339), .Y(n_406) );
INVxp67_ASAP7_75t_L g342 ( .A(n_279), .Y(n_342) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g412 ( .A(n_281), .B(n_399), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_281), .B(n_362), .Y(n_435) );
INVx1_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_283), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g428 ( .A(n_283), .B(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B(n_291), .Y(n_284) );
AND2x2_ASAP7_75t_L g297 ( .A(n_286), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g381 ( .A(n_290), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g399 ( .A(n_292), .B(n_357), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_292), .B(n_356), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_293), .B(n_305), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_299), .C(n_309), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_295), .A2(n_330), .B1(n_334), .B2(n_337), .C(n_340), .Y(n_329) );
AOI31xp33_ASAP7_75t_L g424 ( .A1(n_295), .A2(n_425), .A3(n_426), .B(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B1(n_305), .B2(n_307), .Y(n_299) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g425 ( .A(n_305), .Y(n_425) );
INVx1_ASAP7_75t_L g388 ( .A(n_306), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_308), .A2(n_432), .B(n_434), .C(n_436), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_313), .B2(n_317), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_314), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_316), .A2(n_350), .B1(n_369), .B2(n_405), .C(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g400 ( .A(n_317), .Y(n_400) );
INVx1_ASAP7_75t_L g354 ( .A(n_318), .Y(n_354) );
NAND3xp33_ASAP7_75t_SL g319 ( .A(n_320), .B(n_329), .C(n_344), .Y(n_319) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_321), .A2(n_371), .B(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_323), .B(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g430 ( .A(n_324), .Y(n_430) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g368 ( .A(n_331), .B(n_351), .Y(n_368) );
INVx1_ASAP7_75t_L g343 ( .A(n_332), .Y(n_343) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g341 ( .A(n_335), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_335), .B(n_373), .Y(n_372) );
NOR4xp25_ASAP7_75t_L g340 ( .A(n_336), .B(n_341), .C(n_342), .D(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B1(n_355), .B2(n_356), .C1(n_358), .C2(n_362), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g442 ( .A(n_346), .Y(n_442) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_358), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g418 ( .A1(n_363), .A2(n_419), .B(n_421), .Y(n_418) );
NOR4xp25_ASAP7_75t_L g364 ( .A(n_365), .B(n_376), .C(n_389), .D(n_404), .Y(n_364) );
OAI221xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B1(n_368), .B2(n_369), .C(n_370), .Y(n_365) );
INVx1_ASAP7_75t_L g445 ( .A(n_366), .Y(n_445) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_373), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
OAI222xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B1(n_382), .B2(n_383), .C1(n_386), .C2(n_388), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_412), .B(n_413), .C(n_424), .Y(n_411) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .B1(n_396), .B2(n_398), .C1(n_400), .C2(n_401), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_406), .A2(n_409), .B1(n_442), .B2(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_439), .B(n_441), .C(n_444), .Y(n_436) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_447), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_679), .Y(n_447) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_616), .C(n_650), .D(n_666), .Y(n_448) );
NAND4xp25_ASAP7_75t_SL g449 ( .A(n_450), .B(n_546), .C(n_580), .D(n_596), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_489), .B1(n_522), .B2(n_534), .C1(n_539), .C2(n_545), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI31xp33_ASAP7_75t_L g712 ( .A1(n_452), .A2(n_713), .A3(n_714), .B(n_716), .Y(n_712) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_465), .Y(n_452) );
AND2x2_ASAP7_75t_L g687 ( .A(n_453), .B(n_467), .Y(n_687) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_SL g538 ( .A(n_454), .Y(n_538) );
AND2x2_ASAP7_75t_L g545 ( .A(n_454), .B(n_477), .Y(n_545) );
AND2x2_ASAP7_75t_L g601 ( .A(n_454), .B(n_468), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_465), .B(n_631), .Y(n_630) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_466), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_466), .B(n_549), .Y(n_591) );
AND2x2_ASAP7_75t_L g684 ( .A(n_466), .B(n_624), .Y(n_684) );
OAI321xp33_ASAP7_75t_L g718 ( .A1(n_466), .A2(n_538), .A3(n_691), .B1(n_719), .B2(n_721), .C(n_722), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_466), .B(n_525), .C(n_631), .D(n_723), .Y(n_722) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
AND2x2_ASAP7_75t_L g586 ( .A(n_467), .B(n_536), .Y(n_586) );
AND2x2_ASAP7_75t_L g605 ( .A(n_467), .B(n_538), .Y(n_605) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g537 ( .A(n_468), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g561 ( .A(n_468), .B(n_477), .Y(n_561) );
AND2x2_ASAP7_75t_L g647 ( .A(n_468), .B(n_536), .Y(n_647) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_476), .Y(n_468) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_469), .A2(n_495), .B(n_501), .Y(n_494) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_469), .A2(n_515), .B(n_521), .Y(n_514) );
INVx3_ASAP7_75t_SL g536 ( .A(n_477), .Y(n_536) );
AND2x2_ASAP7_75t_L g579 ( .A(n_477), .B(n_566), .Y(n_579) );
OR2x2_ASAP7_75t_L g612 ( .A(n_477), .B(n_538), .Y(n_612) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_477), .Y(n_619) );
AND2x2_ASAP7_75t_L g648 ( .A(n_477), .B(n_537), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_477), .B(n_621), .Y(n_663) );
AND2x2_ASAP7_75t_L g695 ( .A(n_477), .B(n_687), .Y(n_695) );
AND2x2_ASAP7_75t_L g704 ( .A(n_477), .B(n_550), .Y(n_704) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_485), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .Y(n_490) );
INVx1_ASAP7_75t_SL g672 ( .A(n_491), .Y(n_672) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g541 ( .A(n_492), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g524 ( .A(n_493), .B(n_504), .Y(n_524) );
AND2x2_ASAP7_75t_L g608 ( .A(n_493), .B(n_526), .Y(n_608) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g578 ( .A(n_494), .B(n_514), .Y(n_578) );
OR2x2_ASAP7_75t_L g589 ( .A(n_494), .B(n_526), .Y(n_589) );
AND2x2_ASAP7_75t_L g615 ( .A(n_494), .B(n_526), .Y(n_615) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_494), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_502), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_502), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g588 ( .A(n_503), .B(n_589), .Y(n_588) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_503), .A2(n_578), .A3(n_584), .B1(n_615), .B2(n_665), .C1(n_675), .C2(n_677), .Y(n_674) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_504), .B(n_525), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_504), .B(n_526), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_504), .B(n_542), .Y(n_595) );
AND2x2_ASAP7_75t_L g649 ( .A(n_504), .B(n_615), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_504), .Y(n_653) );
AND2x2_ASAP7_75t_L g665 ( .A(n_504), .B(n_514), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_504), .B(n_541), .Y(n_697) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_514), .Y(n_562) );
BUFx3_ASAP7_75t_L g576 ( .A(n_505), .Y(n_576) );
AND3x2_ASAP7_75t_L g658 ( .A(n_505), .B(n_638), .C(n_659), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_514), .B(n_524), .C(n_525), .Y(n_523) );
INVx1_ASAP7_75t_SL g542 ( .A(n_514), .Y(n_542) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_514), .Y(n_643) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g637 ( .A(n_524), .B(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g644 ( .A(n_524), .Y(n_644) );
AND2x2_ASAP7_75t_L g682 ( .A(n_525), .B(n_660), .Y(n_682) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
AND2x2_ASAP7_75t_L g638 ( .A(n_526), .B(n_542), .Y(n_638) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OR2x2_ASAP7_75t_L g582 ( .A(n_536), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g701 ( .A(n_536), .B(n_601), .Y(n_701) );
AND2x2_ASAP7_75t_L g715 ( .A(n_536), .B(n_538), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_537), .B(n_550), .Y(n_656) );
AND2x2_ASAP7_75t_L g703 ( .A(n_537), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g566 ( .A(n_538), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g583 ( .A(n_538), .B(n_550), .Y(n_583) );
INVx1_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
AND2x2_ASAP7_75t_L g624 ( .A(n_538), .B(n_550), .Y(n_624) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_540), .A2(n_667), .B1(n_671), .B2(n_673), .C(n_674), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x2_ASAP7_75t_L g570 ( .A(n_541), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_544), .B(n_577), .Y(n_720) );
AOI322xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_562), .A3(n_563), .B1(n_564), .B2(n_570), .C1(n_572), .C2(n_579), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_561), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_549), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_549), .B(n_611), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_549), .A2(n_561), .B(n_635), .C(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_549), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_549), .B(n_605), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_549), .B(n_687), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_549), .B(n_715), .Y(n_714) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_550), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_550), .B(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g676 ( .A(n_550), .B(n_563), .Y(n_676) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B(n_559), .Y(n_550) );
INVx1_ASAP7_75t_L g568 ( .A(n_552), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_559), .Y(n_569) );
INVx1_ASAP7_75t_L g651 ( .A(n_561), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g661 ( .A1(n_561), .A2(n_586), .A3(n_662), .B(n_664), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_561), .B(n_567), .Y(n_713) );
INVx1_ASAP7_75t_SL g574 ( .A(n_562), .Y(n_574) );
AND2x2_ASAP7_75t_L g607 ( .A(n_562), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g688 ( .A(n_562), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g573 ( .A(n_563), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g598 ( .A(n_563), .Y(n_598) );
AND2x2_ASAP7_75t_L g625 ( .A(n_563), .B(n_578), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_563), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g717 ( .A(n_563), .B(n_665), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_565), .B(n_635), .Y(n_708) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g604 ( .A(n_567), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g622 ( .A(n_567), .Y(n_622) );
NAND2xp33_ASAP7_75t_SL g572 ( .A(n_573), .B(n_575), .Y(n_572) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_574), .A2(n_617), .B(n_623), .C(n_639), .Y(n_616) );
OR2x2_ASAP7_75t_L g691 ( .A(n_574), .B(n_672), .Y(n_691) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
CKINVDCx16_ASAP7_75t_R g628 ( .A(n_576), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_576), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g597 ( .A(n_578), .B(n_598), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B(n_587), .C(n_590), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g631 ( .A(n_583), .Y(n_631) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_586), .B(n_624), .Y(n_629) );
INVx1_ASAP7_75t_L g635 ( .A(n_586), .Y(n_635) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g594 ( .A(n_589), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g627 ( .A(n_589), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g689 ( .A(n_589), .Y(n_689) );
AOI21xp33_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_592), .B(n_594), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_592), .A2(n_603), .B(n_606), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .B(n_602), .C(n_609), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_597), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_600), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g613 ( .A(n_601), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_603), .A2(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_608), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g633 ( .A(n_608), .Y(n_633) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_613), .B(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g664 ( .A(n_615), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_621), .B(n_647), .Y(n_673) );
AND2x2_ASAP7_75t_L g686 ( .A(n_621), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g700 ( .A(n_621), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g710 ( .A(n_621), .B(n_648), .Y(n_710) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_626), .C(n_634), .Y(n_623) );
INVx1_ASAP7_75t_L g670 ( .A(n_624), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_630), .B2(n_632), .Y(n_626) );
OR2x2_ASAP7_75t_L g632 ( .A(n_628), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_628), .B(n_689), .Y(n_711) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g705 ( .A(n_638), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_645), .B1(n_648), .B2(n_649), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g723 ( .A(n_643), .Y(n_723) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g669 ( .A(n_647), .Y(n_669) );
OAI211xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_654), .C(n_661), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_669), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR5xp2_ASAP7_75t_L g679 ( .A(n_680), .B(n_698), .C(n_706), .D(n_712), .E(n_718), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_683), .B(n_685), .C(n_692), .Y(n_680) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_690), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_695), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .B(n_705), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g721 ( .A(n_701), .Y(n_721) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_711), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g737 ( .A(n_733), .Y(n_737) );
INVx3_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g755 ( .A(n_743), .Y(n_755) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_749), .B1(n_750), .B2(n_753), .Y(n_744) );
INVx1_ASAP7_75t_L g753 ( .A(n_745), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g762 ( .A(n_758), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
endmodule