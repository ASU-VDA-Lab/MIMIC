module fake_jpeg_4984_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_16),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_46),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_21),
.B1(n_19),
.B2(n_36),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_67),
.B1(n_20),
.B2(n_26),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_32),
.B(n_21),
.C(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_37),
.B1(n_26),
.B2(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_19),
.B1(n_36),
.B2(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_69),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_73),
.B(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_28),
.B(n_35),
.C(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_54),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_46),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_33),
.Y(n_110)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_37),
.B1(n_19),
.B2(n_61),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_99),
.B1(n_56),
.B2(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_62),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_25),
.B(n_54),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_80),
.CI(n_72),
.CON(n_134),
.SN(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_62),
.B1(n_60),
.B2(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_115),
.B1(n_116),
.B2(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_110),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_58),
.B1(n_42),
.B2(n_60),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_72),
.B1(n_76),
.B2(n_93),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_82),
.B1(n_78),
.B2(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_25),
.B1(n_20),
.B2(n_34),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_33),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_97),
.B(n_76),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_35),
.B1(n_23),
.B2(n_27),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_35),
.B1(n_23),
.B2(n_27),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_92),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_35),
.B1(n_23),
.B2(n_27),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_81),
.B1(n_71),
.B2(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_132),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_113),
.B1(n_122),
.B2(n_111),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_72),
.C(n_80),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_39),
.C(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_136),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_79),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_141),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_138),
.A2(n_17),
.B1(n_28),
.B2(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_108),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_154),
.B1(n_157),
.B2(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_146),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_90),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_152),
.B1(n_106),
.B2(n_105),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_49),
.B1(n_98),
.B2(n_91),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_98),
.B1(n_49),
.B2(n_83),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_96),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_117),
.B(n_126),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_159),
.A2(n_164),
.B(n_186),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_117),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_176),
.C(n_180),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_189),
.B(n_192),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_126),
.B(n_104),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_104),
.A3(n_115),
.B1(n_127),
.B2(n_124),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_169),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_168),
.B1(n_175),
.B2(n_178),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_40),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_138),
.B1(n_153),
.B2(n_148),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_114),
.B1(n_118),
.B2(n_90),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_42),
.B1(n_17),
.B2(n_28),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_12),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_28),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_150),
.B1(n_143),
.B2(n_139),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_17),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_187),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_0),
.C(n_1),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_146),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_14),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_188),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_0),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_153),
.A2(n_11),
.B1(n_12),
.B2(n_4),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_138),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_197),
.B1(n_210),
.B2(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_201),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_144),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_202),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_134),
.B1(n_151),
.B2(n_140),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_215),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_213),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_135),
.B1(n_134),
.B2(n_151),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_168),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_135),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_162),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_214),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_164),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_180),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_2),
.B(n_3),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_186),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_160),
.B(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_185),
.Y(n_226)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_220),
.A2(n_181),
.B1(n_191),
.B2(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_229),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_176),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_198),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_227),
.C(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_207),
.B(n_159),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_220),
.A2(n_191),
.B1(n_204),
.B2(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_165),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_234),
.B(n_5),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

AOI22x1_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_177),
.B1(n_189),
.B2(n_192),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_239),
.B(n_224),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_204),
.A2(n_173),
.B1(n_161),
.B2(n_4),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_7),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_173),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_244),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_5),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_221),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_198),
.C(n_193),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_230),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_222),
.C(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_253),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_222),
.C(n_208),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_203),
.B1(n_201),
.B2(n_208),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_231),
.B1(n_233),
.B2(n_235),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_269),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_205),
.C(n_196),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_264),
.C(n_248),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_196),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_214),
.B1(n_6),
.B2(n_7),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_223),
.B1(n_229),
.B2(n_228),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_6),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_241),
.B(n_245),
.C(n_9),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_6),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_224),
.B(n_245),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_281),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_264),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_231),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_258),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_286),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_226),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_236),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_236),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_267),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_279),
.A2(n_268),
.B1(n_261),
.B2(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_292),
.B1(n_299),
.B2(n_272),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_255),
.B1(n_259),
.B2(n_257),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_251),
.C(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.C(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_252),
.C(n_238),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_300),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_10),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_277),
.B(n_10),
.CI(n_281),
.CON(n_302),
.SN(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_276),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_310),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_274),
.C(n_284),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_277),
.B(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_313),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_271),
.B(n_280),
.C(n_274),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_315),
.B1(n_295),
.B2(n_296),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_10),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_297),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_312),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_324),
.B1(n_304),
.B2(n_312),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_290),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_305),
.B(n_293),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_311),
.Y(n_325)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_329),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_303),
.B1(n_308),
.B2(n_307),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_314),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_327),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_330),
.B(n_331),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_319),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_333),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_334),
.B(n_317),
.Y(n_340)
);


endmodule