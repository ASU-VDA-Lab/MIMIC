module fake_jpeg_6555_n_166 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_3),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_26),
.Y(n_55)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_40),
.Y(n_45)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_2),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_24),
.B(n_22),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_20),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_29),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_76)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_32),
.A2(n_15),
.B1(n_17),
.B2(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_15),
.B1(n_25),
.B2(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_25),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_3),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_79),
.B1(n_88),
.B2(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_60),
.B1(n_55),
.B2(n_45),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_57),
.B(n_70),
.C(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_89),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_10),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_92),
.B(n_78),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_11),
.B1(n_53),
.B2(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_98),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AO22x2_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_52),
.B1(n_59),
.B2(n_48),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_52),
.C(n_69),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_103),
.C(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_71),
.C(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_71),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_114),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_121),
.C(n_123),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_92),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_76),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_87),
.C(n_73),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_105),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_99),
.C(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_108),
.C(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_133),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_99),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_132),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_120),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_135),
.B(n_138),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_89),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_111),
.C(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_138),
.A2(n_117),
.B1(n_125),
.B2(n_118),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_146),
.Y(n_150)
);

AOI21x1_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_125),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_141),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_130),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_121),
.C(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_144),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_135),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_128),
.C(n_116),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_142),
.B(n_143),
.C(n_148),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_156),
.B(n_78),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_158),
.B(n_109),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_160),
.B(n_161),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_157),
.B(n_84),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_84),
.C(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_164),
.Y(n_166)
);


endmodule