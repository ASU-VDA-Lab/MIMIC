module real_jpeg_24885_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_21),
.B1(n_25),
.B2(n_34),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_21),
.B1(n_25),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_52),
.B1(n_80),
.B2(n_81),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_25),
.B(n_43),
.C(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_24),
.B(n_79),
.C(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_37),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_33),
.C(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_4),
.B(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_11),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_4),
.B(n_65),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_21),
.B1(n_25),
.B2(n_37),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_116),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_115),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_73),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_73),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_53),
.C(n_60),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_17),
.B(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_39),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_26),
.C(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_20),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_21),
.A2(n_25),
.B1(n_43),
.B2(n_46),
.Y(n_49)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_23),
.A2(n_25),
.B(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_23),
.A2(n_24),
.B1(n_99),
.B2(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_35),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_27),
.B(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_33),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_32),
.A2(n_33),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_33),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_35),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_38),
.B(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_36),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_44),
.B(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_38),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_41),
.B(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_45),
.B1(n_66),
.B2(n_67),
.Y(n_72)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_45),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_48),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_53),
.B(n_60),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_54),
.A2(n_56),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_54),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_56),
.Y(n_176)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_59),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_62),
.A2(n_64),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_63),
.B(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_65),
.B(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_69),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_71),
.B(n_133),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_90),
.B2(n_91),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_89),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_103),
.B1(n_104),
.B2(n_114),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_109),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_179),
.B(n_183),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_165),
.B(n_178),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_145),
.B(n_164),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_136),
.B2(n_144),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_135),
.C(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_153),
.B(n_163),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_159),
.B(n_162),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_173),
.C(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);


endmodule