module real_jpeg_17122_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_295;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_7),
.B1(n_19),
.B2(n_21),
.Y(n_18)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_1),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_1),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_1),
.B(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_2),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_3),
.Y(n_262)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_4),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_5),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_5),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_9),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_10),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_11),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_39),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_12),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_12),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_12),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_12),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_12),
.B(n_255),
.Y(n_254)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_15),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_16),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_16),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_16),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_16),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_16),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_16),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_177),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_176),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_148),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_24),
.B(n_148),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_104),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_67),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_48),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_47),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_35),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_35),
.B(n_118),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_35),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.C(n_56),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_82),
.C(n_93),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_68),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_77),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

MAJx3_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_74),
.C(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_81),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_85),
.Y(n_238)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_85),
.Y(n_253)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_91),
.Y(n_276)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_94),
.A2(n_100),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_95),
.B(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_99),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_101),
.Y(n_270)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_135),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_123),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_110),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_116),
.B(n_122),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_130),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_125),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_126),
.B(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_127),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_156),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_149),
.A2(n_150),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_152),
.A2(n_153),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.C(n_163),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_157),
.B(n_161),
.C(n_163),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_163),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.C(n_174),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_164),
.A2(n_165),
.B1(n_174),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_168),
.B(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21x1_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_287),
.B(n_295),
.Y(n_178)
);

AOI21x1_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_231),
.B(n_286),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_207),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_181),
.B(n_207),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_205),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_183),
.B(n_187),
.C(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.C(n_198),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_205),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_228),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_220),
.C(n_224),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_247),
.B(n_285),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_245),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_233),
.B(n_245),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.C(n_243),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_243),
.B1(n_244),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_239),
.Y(n_257)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_279),
.B(n_284),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_267),
.B(n_278),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_250),
.B(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_272),
.B(n_277),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_271),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_293),
.Y(n_295)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);


endmodule