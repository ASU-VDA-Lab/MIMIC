module fake_jpeg_21923_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_240;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_41),
.Y(n_57)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AND2x4_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_1),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_50),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_19),
.B1(n_30),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_36),
.B1(n_30),
.B2(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_62),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_65),
.B1(n_42),
.B2(n_35),
.Y(n_72)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_75),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_53),
.B(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_33),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_76),
.B1(n_20),
.B2(n_27),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_36),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_57),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_111),
.B(n_90),
.C(n_102),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_49),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_99),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_57),
.B1(n_36),
.B2(n_55),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_38),
.B1(n_40),
.B2(n_47),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_36),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_84),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_66),
.B1(n_47),
.B2(n_56),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_83),
.B1(n_89),
.B2(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_122),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_126),
.B1(n_130),
.B2(n_136),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_20),
.B(n_17),
.Y(n_157)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_120),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_88),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_44),
.B(n_30),
.C(n_35),
.D(n_48),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_58),
.C(n_41),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_44),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_129),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_96),
.B1(n_90),
.B2(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

AO21x2_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_86),
.B(n_69),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_106),
.B1(n_77),
.B2(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_77),
.B1(n_69),
.B2(n_35),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_78),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_78),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_142),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_82),
.B(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_147),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_52),
.B1(n_58),
.B2(n_77),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_130),
.B1(n_118),
.B2(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_131),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_150),
.B1(n_156),
.B2(n_162),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_132),
.B1(n_123),
.B2(n_116),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_35),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_130),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_38),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_105),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_40),
.B1(n_100),
.B2(n_82),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_126),
.C(n_117),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_175),
.C(n_150),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_178),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_130),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_130),
.B(n_86),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_185),
.B1(n_149),
.B2(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_120),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_164),
.B(n_24),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_3),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_201),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_194),
.B1(n_208),
.B2(n_171),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_151),
.C(n_140),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_157),
.B1(n_153),
.B2(n_143),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_153),
.C(n_43),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_43),
.C(n_68),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_209),
.C(n_22),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_68),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_24),
.B1(n_20),
.B2(n_31),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_185),
.B1(n_177),
.B2(n_21),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_94),
.B1(n_31),
.B2(n_28),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_94),
.Y(n_209)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_172),
.B1(n_173),
.B2(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_218),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_171),
.B1(n_28),
.B2(n_23),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_189),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_23),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_14),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_223),
.C(n_195),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_22),
.C(n_21),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_224),
.B(n_200),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_204),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_225),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_4),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_191),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.C(n_222),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_201),
.C(n_15),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_7),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_4),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_223),
.C(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_219),
.C(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_218),
.C(n_217),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_217),
.C(n_225),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_233),
.B1(n_228),
.B2(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_255),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_239),
.B(n_229),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_256),
.B(n_8),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_7),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_7),
.B(n_8),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_8),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_9),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_260),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_263),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_10),
.C(n_11),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_10),
.B(n_11),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_255),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_253),
.B(n_11),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_264),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_266),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_270),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_268),
.B(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_10),
.C(n_12),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_273),
.A2(n_12),
.B(n_13),
.Y(n_274)
);


endmodule