module fake_jpeg_32058_n_532 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_532);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_17),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_22),
.A2(n_8),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_58),
.B(n_9),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_18),
.B(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_7),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_7),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_80),
.Y(n_134)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_7),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_21),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_101),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_25),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_39),
.B(n_29),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_107),
.A2(n_154),
.B1(n_160),
.B2(n_165),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_59),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_130),
.B(n_140),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_80),
.A2(n_47),
.B1(n_37),
.B2(n_44),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_153),
.B1(n_97),
.B2(n_102),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_28),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_24),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_49),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_146),
.B(n_149),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_28),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_54),
.A2(n_37),
.B1(n_44),
.B2(n_36),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_56),
.A2(n_52),
.B1(n_21),
.B2(n_50),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_52),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_57),
.A2(n_49),
.B1(n_45),
.B2(n_31),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_75),
.A2(n_51),
.B1(n_37),
.B2(n_38),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_167),
.A2(n_176),
.B1(n_197),
.B2(n_217),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_169),
.B(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_183),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_109),
.A2(n_67),
.B1(n_100),
.B2(n_89),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_181),
.B(n_190),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_117),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_182),
.B(n_187),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_134),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_87),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_24),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_196),
.B(n_200),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_125),
.A2(n_74),
.B1(n_88),
.B2(n_84),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_198),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_134),
.B(n_29),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_143),
.A2(n_73),
.A3(n_33),
.B1(n_22),
.B2(n_27),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_178),
.Y(n_222)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_208),
.B(n_215),
.Y(n_249)
);

BUFx4f_ASAP7_75t_SL g209 ( 
.A(n_142),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_133),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_219),
.B1(n_220),
.B2(n_145),
.Y(n_224)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

BUFx4f_ASAP7_75t_SL g214 ( 
.A(n_113),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_144),
.A2(n_83),
.B1(n_79),
.B2(n_78),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_222),
.B(n_121),
.Y(n_273)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_167),
.B1(n_197),
.B2(n_163),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_229),
.A2(n_231),
.B1(n_251),
.B2(n_179),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_153),
.B1(n_135),
.B2(n_132),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_129),
.B(n_113),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_253),
.B(n_209),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_135),
.B1(n_151),
.B2(n_163),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_258),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_151),
.B1(n_145),
.B2(n_161),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_244),
.A2(n_198),
.B1(n_164),
.B2(n_194),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_180),
.A2(n_133),
.B1(n_156),
.B2(n_147),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_177),
.A2(n_129),
.B(n_101),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_33),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_26),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_147),
.B1(n_156),
.B2(n_161),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_264),
.A2(n_271),
.B1(n_276),
.B2(n_277),
.Y(n_312)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_207),
.C(n_27),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_266),
.B(n_288),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_231),
.A2(n_207),
.B1(n_199),
.B2(n_174),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_168),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_278),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_272),
.B1(n_298),
.B2(n_262),
.Y(n_303)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_273),
.B(n_279),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_188),
.C(n_220),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_281),
.C(n_257),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_209),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_296),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_222),
.A2(n_72),
.B1(n_165),
.B2(n_211),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_246),
.A2(n_206),
.B1(n_152),
.B2(n_213),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_38),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_280),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_234),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_226),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_283),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_240),
.B1(n_256),
.B2(n_242),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_235),
.A2(n_195),
.B1(n_173),
.B2(n_189),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_293),
.B1(n_242),
.B2(n_257),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_214),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_286),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_214),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_241),
.A2(n_26),
.A3(n_40),
.B1(n_30),
.B2(n_66),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_248),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_40),
.B(n_30),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_292),
.B(n_262),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_40),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_300),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_251),
.A2(n_30),
.B1(n_51),
.B2(n_48),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_235),
.A2(n_262),
.B1(n_228),
.B2(n_254),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_221),
.B(n_9),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_5),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_48),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_221),
.B(n_9),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_297),
.B(n_0),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_48),
.B1(n_10),
.B2(n_2),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_243),
.B(n_256),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_303),
.A2(n_299),
.B1(n_271),
.B2(n_264),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_305),
.B(n_322),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_296),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_227),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_324),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_321),
.B1(n_283),
.B2(n_259),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_240),
.B(n_252),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_313),
.A2(n_292),
.B(n_282),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_315),
.A2(n_267),
.B1(n_278),
.B2(n_279),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_272),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_252),
.C(n_232),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_296),
.C(n_271),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_228),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_319),
.B(n_259),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_284),
.A2(n_260),
.B1(n_227),
.B2(n_232),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_291),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_330),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_236),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_268),
.B(n_236),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_328),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_260),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_334),
.A2(n_299),
.B1(n_276),
.B2(n_270),
.Y(n_346)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_337),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_343),
.B1(n_334),
.B2(n_321),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_347),
.C(n_354),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_340),
.A2(n_360),
.B(n_309),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_328),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_344),
.B(n_351),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_346),
.A2(n_350),
.B1(n_331),
.B2(n_333),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_297),
.Y(n_349)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_280),
.C(n_225),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_289),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_310),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_326),
.Y(n_371)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_294),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_364),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_287),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_365),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_263),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_318),
.C(n_306),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_263),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_312),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_287),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_316),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_371),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_377),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_306),
.C(n_313),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_376),
.B(n_378),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_352),
.B(n_320),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_330),
.C(n_302),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_302),
.C(n_312),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_379),
.B(n_382),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_395),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_332),
.C(n_309),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_304),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_400),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_387),
.A2(n_389),
.B1(n_350),
.B2(n_346),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_343),
.A2(n_309),
.B1(n_316),
.B2(n_329),
.Y(n_389)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_393),
.A2(n_399),
.B(n_340),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_323),
.Y(n_394)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_305),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_397),
.A2(n_336),
.B1(n_356),
.B2(n_355),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_348),
.B(n_329),
.Y(n_398)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_398),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_360),
.A2(n_230),
.B(n_223),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_368),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_339),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_410),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_340),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_404),
.Y(n_441)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_407),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_409),
.A2(n_372),
.B1(n_387),
.B2(n_369),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_358),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_411),
.A2(n_414),
.B1(n_416),
.B2(n_418),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_336),
.B1(n_358),
.B2(n_359),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_381),
.A2(n_364),
.B(n_342),
.Y(n_415)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_384),
.A2(n_365),
.B1(n_362),
.B2(n_345),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_357),
.B1(n_345),
.B2(n_342),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_382),
.A2(n_363),
.B(n_337),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_SL g429 ( 
.A1(n_419),
.A2(n_425),
.B(n_399),
.C(n_389),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_390),
.Y(n_422)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_223),
.Y(n_423)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

AOI22x1_ASAP7_75t_SL g425 ( 
.A1(n_393),
.A2(n_223),
.B1(n_238),
.B2(n_230),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_378),
.A2(n_261),
.B(n_225),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_426),
.B(n_427),
.Y(n_431)
);

NOR3xp33_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_223),
.C(n_238),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_428),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_429),
.B(n_432),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_376),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_434),
.A2(n_449),
.B1(n_411),
.B2(n_418),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_420),
.B(n_377),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_437),
.B(n_445),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_401),
.B(n_379),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_419),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_375),
.C(n_395),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_443),
.C(n_446),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_372),
.C(n_388),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_423),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_410),
.C(n_402),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_369),
.C(n_385),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_416),
.C(n_422),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_413),
.Y(n_448)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_448),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_409),
.A2(n_370),
.B1(n_385),
.B2(n_396),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_449),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_435),
.A2(n_405),
.B(n_425),
.Y(n_454)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_456),
.B(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_450),
.Y(n_457)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_442),
.A2(n_406),
.B1(n_421),
.B2(n_404),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_461),
.B1(n_467),
.B2(n_434),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_404),
.B1(n_407),
.B2(n_414),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_462),
.B(n_463),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_448),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_447),
.B(n_370),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_465),
.Y(n_482)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_415),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_438),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_441),
.B1(n_435),
.B2(n_430),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_431),
.A2(n_374),
.B(n_261),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_469),
.A2(n_374),
.B(n_433),
.Y(n_473)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_473),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_472),
.A2(n_478),
.B1(n_454),
.B2(n_459),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_436),
.C(n_432),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_484),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_477),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_440),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_429),
.B1(n_446),
.B2(n_238),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_468),
.Y(n_489)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_483),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_238),
.C(n_48),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_10),
.Y(n_486)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

INVx11_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_487),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_502),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_453),
.Y(n_490)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_490),
.B1(n_500),
.B2(n_488),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_458),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_499),
.Y(n_507)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_462),
.B(n_467),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_494),
.A2(n_3),
.B(n_5),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_457),
.Y(n_495)
);

OAI22x1_ASAP7_75t_L g508 ( 
.A1(n_495),
.A2(n_473),
.B1(n_487),
.B2(n_472),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_474),
.A2(n_461),
.B1(n_456),
.B2(n_2),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_480),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_48),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_504),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_475),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_509),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_508),
.A2(n_496),
.B1(n_3),
.B2(n_11),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_497),
.B(n_484),
.Y(n_509)
);

BUFx4f_ASAP7_75t_SL g510 ( 
.A(n_499),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_513),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_498),
.A2(n_477),
.B(n_476),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_512),
.B(n_498),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_514),
.A2(n_516),
.B(n_509),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_505),
.A2(n_507),
.B(n_506),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_502),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_515),
.C(n_517),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_520),
.A2(n_510),
.B1(n_518),
.B2(n_516),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_524),
.C(n_16),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_523),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_SL g524 ( 
.A1(n_519),
.A2(n_3),
.B(n_14),
.C(n_16),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_16),
.B(n_0),
.Y(n_527)
);

AOI21xp33_ASAP7_75t_SL g528 ( 
.A1(n_527),
.A2(n_525),
.B(n_16),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_0),
.C(n_1),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_0),
.B(n_1),
.Y(n_530)
);

NAND2x1_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_1),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_1),
.Y(n_532)
);


endmodule