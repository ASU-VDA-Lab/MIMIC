module fake_jpeg_8844_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx8_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_70),
.Y(n_75)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_0),
.Y(n_77)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_37),
.B1(n_61),
.B2(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_98),
.B1(n_99),
.B2(n_60),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_97),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_80),
.B(n_56),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_51),
.B1(n_62),
.B2(n_48),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_57),
.B1(n_58),
.B2(n_45),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_112),
.B1(n_119),
.B2(n_122),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_44),
.B(n_43),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_44),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_3),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_125)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_74),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_42),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_102),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_127),
.B(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_111),
.C(n_110),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_106),
.B(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_6),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_8),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_115),
.B(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_95),
.B1(n_114),
.B2(n_103),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_59),
.A3(n_40),
.B1(n_120),
.B2(n_47),
.C(n_17),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_107),
.B(n_104),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_10),
.B(n_12),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_13),
.B(n_16),
.Y(n_143)
);


endmodule