module fake_jpeg_22990_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_49),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_32),
.B1(n_23),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_67),
.B1(n_29),
.B2(n_19),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_32),
.B1(n_23),
.B2(n_19),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_73),
.B1(n_48),
.B2(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_35),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_25),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_32),
.B1(n_23),
.B2(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_23),
.B1(n_29),
.B2(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_82),
.Y(n_144)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_83),
.Y(n_139)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_85),
.A2(n_99),
.B1(n_100),
.B2(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_93),
.B1(n_34),
.B2(n_26),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_63),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

NAND2xp67_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_48),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_29),
.B1(n_20),
.B2(n_35),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_97),
.B1(n_109),
.B2(n_30),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_37),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_101),
.C(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_51),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_48),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_113),
.B(n_34),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_45),
.A3(n_35),
.B1(n_21),
.B2(n_28),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_30),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_40),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_57),
.A2(n_28),
.B1(n_21),
.B2(n_34),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_46),
.C(n_43),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_69),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_74),
.B(n_46),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_21),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_63),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_18),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_50),
.B1(n_43),
.B2(n_18),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_103),
.B1(n_99),
.B2(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_93),
.B1(n_97),
.B2(n_89),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_132),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_149),
.Y(n_168)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_76),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_85),
.B1(n_111),
.B2(n_102),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_78),
.B(n_31),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_81),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_79),
.A2(n_22),
.B(n_30),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_158),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_159),
.B1(n_164),
.B2(n_144),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_157),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_89),
.B1(n_118),
.B2(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_166),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_131),
.C(n_120),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_178),
.C(n_180),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_101),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_144),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_119),
.B1(n_127),
.B2(n_132),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_139),
.B1(n_133),
.B2(n_88),
.Y(n_208)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_169),
.B(n_172),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_89),
.B1(n_118),
.B2(n_110),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_126),
.B1(n_147),
.B2(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_114),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_75),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_173),
.B(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_112),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_122),
.A2(n_105),
.B(n_118),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_18),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_96),
.C(n_84),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_96),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_160),
.B(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_117),
.C(n_82),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_190),
.B1(n_198),
.B2(n_208),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_186),
.B(n_188),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_147),
.B(n_136),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_136),
.B(n_138),
.Y(n_188)
);

XOR2x2_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_134),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_123),
.B1(n_148),
.B2(n_142),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_148),
.C(n_101),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_18),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_162),
.C(n_172),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_150),
.C(n_161),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_195),
.A2(n_196),
.B(n_206),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_130),
.B(n_7),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_142),
.B1(n_94),
.B2(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_204),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

OAI22x1_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_94),
.B1(n_31),
.B2(n_24),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_213),
.B1(n_124),
.B2(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_124),
.B1(n_116),
.B2(n_22),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_179),
.B(n_180),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_218),
.B(n_222),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_168),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_164),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_228),
.C(n_242),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_179),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_153),
.B(n_151),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_239),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_227),
.A2(n_231),
.B1(n_237),
.B2(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_22),
.C(n_26),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_27),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_26),
.B(n_27),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_31),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_236),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_183),
.B(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_186),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_31),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_185),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_0),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_9),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_24),
.C(n_1),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_243),
.B(n_251),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_182),
.C(n_187),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.C(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_187),
.C(n_205),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_201),
.B1(n_208),
.B2(n_213),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_226),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_205),
.C(n_188),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_207),
.B1(n_200),
.B2(n_210),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_255),
.B1(n_266),
.B2(n_227),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_200),
.B1(n_212),
.B2(n_24),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_7),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_263),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_225),
.A2(n_0),
.B(n_1),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_10),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_221),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_222),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_278),
.Y(n_298)
);

XOR2x2_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_240),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_271),
.B(n_287),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_225),
.C(n_228),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_218),
.C(n_221),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_242),
.C(n_214),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_214),
.B1(n_224),
.B2(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_233),
.B1(n_234),
.B2(n_4),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_258),
.B1(n_257),
.B2(n_254),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_2),
.C(n_3),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_2),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_259),
.C(n_249),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_296),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_264),
.B(n_245),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_300),
.B(n_302),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_281),
.A2(n_245),
.B(n_4),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_12),
.B(n_15),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_274),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_287),
.B1(n_284),
.B2(n_272),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_306),
.B(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_269),
.C(n_270),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.C(n_316),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_317),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_271),
.B(n_268),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_277),
.B1(n_283),
.B2(n_276),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_269),
.B(n_285),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_279),
.CI(n_6),
.CON(n_314),
.SN(n_314)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_297),
.B1(n_303),
.B2(n_12),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_288),
.C(n_299),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_11),
.B(n_12),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_298),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_300),
.Y(n_319)
);

OAI22x1_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_321),
.B1(n_328),
.B2(n_307),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_296),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_327),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_304),
.B1(n_289),
.B2(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_302),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_315),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_316),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_319),
.B(n_308),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_324),
.C(n_323),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_314),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_13),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_11),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_337),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_323),
.B(n_321),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_340),
.B(n_329),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_338),
.B(n_336),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_342),
.B1(n_338),
.B2(n_14),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_344),
.Y(n_345)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_345),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_13),
.Y(n_347)
);


endmodule