module fake_netlist_1_1245_n_33 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_6), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_7), .B(n_9), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_5), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
OR2x2_ASAP7_75t_L g20 ( .A(n_12), .B(n_0), .Y(n_20) );
NAND3xp33_ASAP7_75t_SL g21 ( .A(n_14), .B(n_0), .C(n_1), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_13), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_13), .Y(n_23) );
OAI321xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_21), .A3(n_19), .B1(n_18), .B2(n_16), .C(n_17), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_26), .B(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_18), .Y(n_28) );
AND2x2_ASAP7_75t_SL g29 ( .A(n_28), .B(n_1), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_15), .B1(n_2), .B2(n_3), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
AOI22xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_7), .B1(n_30), .B2(n_11), .Y(n_33) );
endmodule