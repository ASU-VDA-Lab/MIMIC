module fake_jpeg_29732_n_356 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_17),
.Y(n_82)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_16),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_67),
.Y(n_75)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_40),
.B1(n_21),
.B2(n_2),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_61),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_62),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_13),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_25),
.A2(n_14),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_26),
.Y(n_83)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_42),
.B1(n_37),
.B2(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_74),
.A2(n_91),
.B1(n_96),
.B2(n_115),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_33),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_86),
.B(n_88),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_33),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_105),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_42),
.B1(n_31),
.B2(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_92),
.B(n_4),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_44),
.A2(n_42),
.B1(n_24),
.B2(n_18),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_44),
.A2(n_24),
.B1(n_18),
.B2(n_33),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_110),
.B1(n_73),
.B2(n_87),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_18),
.C(n_23),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_76),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_34),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_47),
.A2(n_30),
.B1(n_23),
.B2(n_39),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_27),
.B1(n_39),
.B2(n_22),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_0),
.B(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_39),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_40),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_47),
.A2(n_40),
.B1(n_21),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_116),
.A2(n_62),
.B1(n_60),
.B2(n_21),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_127),
.B1(n_136),
.B2(n_142),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_70),
.B1(n_54),
.B2(n_60),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_133),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_76),
.B(n_81),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_65),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_104),
.B1(n_102),
.B2(n_111),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_54),
.B1(n_70),
.B2(n_49),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_27),
.B1(n_21),
.B2(n_40),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_40),
.A3(n_21),
.B1(n_11),
.B2(n_10),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_143),
.A3(n_138),
.B1(n_131),
.B2(n_135),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_99),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_87),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_0),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_151),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_73),
.B1(n_114),
.B2(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_4),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_157),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_4),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_121),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_133),
.B(n_126),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_168),
.C(n_190),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_111),
.B(n_102),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_136),
.B1(n_135),
.B2(n_129),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_169),
.A2(n_195),
.B(n_6),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_171),
.B(n_181),
.C(n_160),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_180),
.B1(n_191),
.B2(n_193),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_186),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_119),
.A2(n_98),
.B1(n_118),
.B2(n_94),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_189),
.B1(n_139),
.B2(n_154),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_122),
.A2(n_84),
.B1(n_94),
.B2(n_104),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_181),
.B(n_137),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_124),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_84),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_131),
.B(n_95),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_95),
.B1(n_72),
.B2(n_106),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_103),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_130),
.A2(n_106),
.B1(n_117),
.B2(n_73),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_103),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_117),
.B(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_9),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_6),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_129),
.C(n_123),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_142),
.C(n_149),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_208),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_139),
.B1(n_140),
.B2(n_153),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_211),
.B1(n_224),
.B2(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_220),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_157),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_176),
.C(n_184),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_139),
.B1(n_150),
.B2(n_156),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_218),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_195),
.B(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_174),
.B(n_141),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_182),
.B(n_141),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_176),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_182),
.B(n_155),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_187),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_164),
.A2(n_158),
.B1(n_124),
.B2(n_9),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_169),
.A2(n_8),
.B1(n_9),
.B2(n_170),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_161),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_230),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.C(n_171),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_194),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_160),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_250),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_247),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_257),
.B(n_225),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_197),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_239),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_170),
.B1(n_177),
.B2(n_186),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_253),
.B1(n_240),
.B2(n_215),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_193),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_251),
.B(n_204),
.C(n_214),
.D(n_221),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_196),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_197),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_207),
.A2(n_191),
.B1(n_172),
.B2(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_200),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_183),
.B(n_184),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_241),
.B1(n_240),
.B2(n_239),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_247),
.B(n_249),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_204),
.Y(n_266)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_251),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_199),
.C(n_198),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_277),
.C(n_280),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_212),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_275),
.A2(n_244),
.B1(n_201),
.B2(n_205),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_242),
.B(n_245),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_278),
.B(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_210),
.C(n_223),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_224),
.CI(n_215),
.CON(n_278),
.SN(n_278)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_211),
.CI(n_213),
.CON(n_279),
.SN(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_208),
.C(n_222),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_277),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_283),
.A2(n_299),
.B1(n_266),
.B2(n_262),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_295),
.B(n_276),
.Y(n_300)
);

OAI322xp33_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_237),
.A3(n_252),
.B1(n_232),
.B2(n_233),
.C1(n_258),
.C2(n_238),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_288),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_250),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_253),
.B1(n_236),
.B2(n_238),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_296),
.B1(n_260),
.B2(n_278),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_257),
.B(n_255),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_292),
.B(n_298),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_244),
.B(n_229),
.C(n_218),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_250),
.C(n_231),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_297),
.C(n_261),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_231),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_255),
.B(n_237),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_234),
.B1(n_206),
.B2(n_217),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_300),
.A2(n_291),
.B(n_298),
.Y(n_322)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_305),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_274),
.B1(n_267),
.B2(n_271),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_307),
.B1(n_315),
.B2(n_290),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_263),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_306),
.A2(n_310),
.B1(n_312),
.B2(n_314),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_280),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_261),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_260),
.C(n_259),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_259),
.C(n_279),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_293),
.C(n_297),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_283),
.A2(n_278),
.B1(n_279),
.B2(n_275),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_281),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_319),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_321),
.C(n_324),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_289),
.B1(n_284),
.B2(n_294),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_304),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_286),
.C(n_294),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_300),
.B1(n_314),
.B2(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_284),
.B(n_299),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_326),
.A2(n_310),
.B(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_318),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_272),
.B1(n_312),
.B2(n_303),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_329),
.A2(n_331),
.B1(n_321),
.B2(n_326),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_295),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_268),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_324),
.A2(n_303),
.B(n_308),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_340),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_341),
.A2(n_342),
.B(n_344),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_332),
.A2(n_328),
.B(n_336),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_318),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_343),
.B(n_339),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_163),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_188),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_334),
.C(n_331),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_348),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_349),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_353),
.A2(n_342),
.B(n_350),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_352),
.C(n_351),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_348),
.Y(n_356)
);


endmodule