module fake_jpeg_27688_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_SL g59 ( 
.A(n_19),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_15),
.B1(n_40),
.B2(n_39),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_58),
.B1(n_61),
.B2(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_47),
.B1(n_46),
.B2(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_62),
.B1(n_60),
.B2(n_54),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_13),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_61),
.B1(n_50),
.B2(n_65),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_52),
.B1(n_51),
.B2(n_53),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_101),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_64),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_86),
.B1(n_1),
.B2(n_2),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_3),
.Y(n_115)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_99),
.B1(n_105),
.B2(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_115),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_98),
.B1(n_97),
.B2(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_122),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_103),
.C(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_121),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_116),
.B(n_92),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_126),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_128),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_4),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_138),
.B1(n_140),
.B2(n_7),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_18),
.B(n_31),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_24),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_139),
.CI(n_129),
.CON(n_145),
.SN(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_147),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_155),
.B1(n_151),
.B2(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_149),
.B1(n_134),
.B2(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_27),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_25),
.C(n_45),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_22),
.B(n_30),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_16),
.Y(n_165)
);


endmodule