module fake_ariane_2161_n_3113 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_844, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_371, n_845, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_255, n_560, n_450, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_849, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_3113);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_371;
input n_845;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_255;
input n_560;
input n_450;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_849;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_3113;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2702;
wire n_2461;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_3063;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_2867;
wire n_1917;
wire n_2769;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_2909;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_2791;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2683;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_2598;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3052;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_2853;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2774;
wire n_2707;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_3085;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_3024;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_1748;
wire n_873;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3097;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2785;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_2656;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_2723;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_1321;
wire n_3050;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_3107;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2605;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_1116;
wire n_3043;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_2647;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3101;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_3091;
wire n_1024;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_2967;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3111;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_2736;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_2917;
wire n_2544;
wire n_2085;
wire n_2432;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1821;
wire n_1168;
wire n_1310;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_1474;
wire n_937;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_64),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_574),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_667),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_707),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_426),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_671),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_5),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_100),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_130),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_169),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_736),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_735),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_478),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_306),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_782),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_249),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_809),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_773),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_799),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_747),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_316),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_43),
.Y(n_873)
);

INVxp67_ASAP7_75t_R g874 ( 
.A(n_524),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_30),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_192),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_387),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_711),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_336),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_2),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_443),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_389),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_713),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_439),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_726),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_757),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_737),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_47),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_777),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_835),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_719),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_810),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_310),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_686),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_69),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_776),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_119),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_823),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_650),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_291),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_610),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_816),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_341),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_795),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_718),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_813),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_701),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_693),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_753),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_842),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_326),
.Y(n_912)
);

CKINVDCx16_ASAP7_75t_R g913 ( 
.A(n_802),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_355),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_86),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_156),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_812),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_321),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_727),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_195),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_26),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_715),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_140),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_492),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_698),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_441),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_804),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_516),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_526),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_183),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_312),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_331),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_749),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_798),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_699),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_223),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_785),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_70),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_754),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_714),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_594),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_277),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_756),
.Y(n_943)
);

CKINVDCx16_ASAP7_75t_R g944 ( 
.A(n_599),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_771),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_267),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_708),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_55),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_648),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_37),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_225),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_763),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_22),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_349),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_338),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_268),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_515),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_838),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_796),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_636),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_386),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_811),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_712),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_69),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_299),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_740),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_748),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_725),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_298),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_846),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_147),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_284),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_808),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_696),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_697),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_257),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_836),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_797),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_768),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_817),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_761),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_723),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_592),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_502),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_281),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_654),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_681),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_709),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_196),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_783),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_625),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_751),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_722),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_170),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_744),
.Y(n_995)
);

CKINVDCx14_ASAP7_75t_R g996 ( 
.A(n_843),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_703),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_60),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_566),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_334),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_767),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_720),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_194),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_824),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_694),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_39),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_56),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_423),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_787),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_134),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_790),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_732),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_611),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_180),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_779),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_208),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_734),
.Y(n_1017)
);

INVxp33_ASAP7_75t_L g1018 ( 
.A(n_487),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_242),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_745),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_695),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_57),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_833),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_700),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_792),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_414),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_721),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_677),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_605),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_688),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_781),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_772),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_628),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_156),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_704),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_435),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_88),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_358),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_398),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_390),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_774),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_759),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_449),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_324),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_819),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_706),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_769),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_638),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_22),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_15),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_728),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_764),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_512),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_805),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_153),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_433),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_752),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_342),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_620),
.Y(n_1059)
);

BUFx10_ASAP7_75t_L g1060 ( 
.A(n_613),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_755),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_184),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_175),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_248),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_122),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_762),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_786),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_678),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_717),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_504),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_675),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_669),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_730),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_351),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_108),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_658),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_775),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_807),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_292),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_716),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_608),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_832),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_760),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_731),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_821),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_742),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_750),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_187),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_319),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_452),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_477),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_153),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_743),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_680),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_480),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_484),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_333),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_493),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_849),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_814),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_778),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_126),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_765),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_827),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_267),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_40),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_102),
.Y(n_1107)
);

BUFx10_ASAP7_75t_L g1108 ( 
.A(n_788),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_46),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_403),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_826),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_258),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_17),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_325),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_634),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_710),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_357),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_374),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_822),
.Y(n_1119)
);

CKINVDCx14_ASAP7_75t_R g1120 ( 
.A(n_82),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_582),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_766),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_118),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_215),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_724),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_845),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_375),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_583),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_471),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_313),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_784),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_95),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_828),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_365),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_586),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_396),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_152),
.Y(n_1137)
);

CKINVDCx14_ASAP7_75t_R g1138 ( 
.A(n_472),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_550),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_206),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_733),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_653),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_839),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_4),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_430),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_705),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_356),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_87),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_434),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_465),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_400),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_803),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_820),
.Y(n_1153)
);

CKINVDCx16_ASAP7_75t_R g1154 ( 
.A(n_121),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_245),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_746),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_674),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_380),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_758),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_770),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_626),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_266),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_234),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_318),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_825),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_247),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_154),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_800),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_806),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_789),
.Y(n_1170)
);

BUFx2_ASAP7_75t_SL g1171 ( 
.A(n_739),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_794),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_563),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_738),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_829),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_847),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_780),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_195),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_455),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_729),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_831),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_590),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_285),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_322),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_818),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_95),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_110),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_607),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_834),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_29),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_205),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_598),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_18),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_837),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_801),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_793),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_791),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_18),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_848),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_840),
.Y(n_1200)
);

CKINVDCx14_ASAP7_75t_R g1201 ( 
.A(n_297),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_830),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_702),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_97),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_741),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1154),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_921),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_858),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_859),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_861),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1061),
.B(n_0),
.Y(n_1211)
);

INVxp33_ASAP7_75t_L g1212 ( 
.A(n_951),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_875),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1080),
.Y(n_1214)
);

CKINVDCx16_ASAP7_75t_R g1215 ( 
.A(n_1120),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_888),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1201),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_916),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_856),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_892),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_893),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_942),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_976),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_994),
.Y(n_1224)
);

CKINVDCx14_ASAP7_75t_R g1225 ( 
.A(n_996),
.Y(n_1225)
);

INVxp33_ASAP7_75t_SL g1226 ( 
.A(n_860),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1003),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_921),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1010),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1019),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_L g1231 ( 
.A(n_1132),
.B(n_0),
.Y(n_1231)
);

INVxp33_ASAP7_75t_SL g1232 ( 
.A(n_873),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1037),
.B(n_1049),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1063),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1064),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1092),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1102),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1106),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1112),
.Y(n_1239)
);

INVxp33_ASAP7_75t_SL g1240 ( 
.A(n_876),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1144),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_921),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1162),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_909),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1183),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1187),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1204),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_920),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_929),
.Y(n_1249)
);

XOR2xp5_ASAP7_75t_L g1250 ( 
.A(n_852),
.B(n_1),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1124),
.Y(n_1251)
);

INVxp33_ASAP7_75t_L g1252 ( 
.A(n_953),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_964),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_985),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_865),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1050),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1099),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1018),
.Y(n_1258)
);

INVxp33_ASAP7_75t_SL g1259 ( 
.A(n_880),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_952),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1115),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_957),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1028),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_904),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_966),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1242),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1207),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1228),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1248),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1265),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1208),
.Y(n_1272)
);

CKINVDCx16_ASAP7_75t_R g1273 ( 
.A(n_1215),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1254),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1214),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1217),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1258),
.B(n_1138),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1233),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1251),
.Y(n_1279)
);

BUFx8_ASAP7_75t_L g1280 ( 
.A(n_1264),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1209),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1210),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1225),
.B(n_1255),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1213),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1257),
.B(n_913),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1211),
.A2(n_872),
.B(n_857),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1253),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1219),
.Y(n_1288)
);

AND2x6_ASAP7_75t_L g1289 ( 
.A(n_1262),
.B(n_1253),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1216),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1226),
.B(n_944),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1218),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1222),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1256),
.B(n_906),
.Y(n_1294)
);

BUFx8_ASAP7_75t_L g1295 ( 
.A(n_1223),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1206),
.A2(n_956),
.B1(n_867),
.B2(n_1148),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1224),
.Y(n_1297)
);

BUFx8_ASAP7_75t_SL g1298 ( 
.A(n_1249),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1261),
.B(n_927),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1227),
.Y(n_1300)
);

BUFx8_ASAP7_75t_L g1301 ( 
.A(n_1229),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1212),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1230),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1234),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1235),
.B(n_1133),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1232),
.A2(n_1178),
.B1(n_1062),
.B2(n_895),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1236),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1252),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1240),
.A2(n_1195),
.B1(n_1051),
.B2(n_1066),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1237),
.B(n_1028),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1238),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1271),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1277),
.B(n_1259),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1287),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1302),
.B(n_1220),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1275),
.B(n_1278),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1308),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1282),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1273),
.B(n_1221),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1297),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1293),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1270),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1300),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1274),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1269),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1303),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1310),
.B(n_1239),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1304),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1268),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1307),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1272),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1281),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1269),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1284),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1305),
.B(n_1267),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1292),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1279),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1290),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1311),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1289),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1286),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1276),
.B(n_1263),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1289),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1283),
.A2(n_884),
.B(n_881),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1299),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1285),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1294),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1291),
.B(n_1241),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1296),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1288),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1294),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1306),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1295),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1309),
.B(n_1243),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1298),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1301),
.B(n_1244),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1280),
.Y(n_1357)
);

NAND2xp33_ASAP7_75t_SL g1358 ( 
.A(n_1288),
.B(n_1041),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1270),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1271),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1271),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1271),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1271),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1270),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1287),
.B(n_1260),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1271),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1271),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1270),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1287),
.B(n_1266),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1271),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1302),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1286),
.A2(n_889),
.B(n_885),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1271),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1271),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1270),
.Y(n_1375)
);

BUFx8_ASAP7_75t_L g1376 ( 
.A(n_1278),
.Y(n_1376)
);

AND2x6_ASAP7_75t_L g1377 ( 
.A(n_1351),
.B(n_1347),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1322),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1371),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1313),
.B(n_1068),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1371),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1317),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1355),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1346),
.A2(n_1071),
.B1(n_1231),
.B2(n_1042),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1348),
.A2(n_1197),
.B1(n_924),
.B2(n_864),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1359),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1365),
.B(n_1245),
.Y(n_1387)
);

XNOR2xp5_ASAP7_75t_L g1388 ( 
.A(n_1350),
.B(n_1342),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1246),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1364),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1331),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1340),
.B(n_1190),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1343),
.B(n_1191),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1368),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1376),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1351),
.B(n_1193),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1355),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1332),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1334),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1316),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1315),
.Y(n_1401)
);

NOR2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1319),
.B(n_1357),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1369),
.Y(n_1403)
);

BUFx10_ASAP7_75t_L g1404 ( 
.A(n_1337),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1314),
.B(n_1198),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1337),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1375),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1358),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1349),
.B(n_1247),
.Y(n_1409)
);

INVx4_ASAP7_75t_SL g1410 ( 
.A(n_1329),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_SL g1411 ( 
.A(n_1327),
.B(n_897),
.Y(n_1411)
);

INVx4_ASAP7_75t_SL g1412 ( 
.A(n_1329),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1335),
.B(n_853),
.Y(n_1413)
);

BUFx10_ASAP7_75t_L g1414 ( 
.A(n_1352),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1345),
.B(n_900),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1338),
.A2(n_923),
.B1(n_930),
.B2(n_915),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1318),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1354),
.B(n_936),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1321),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1336),
.B(n_938),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1339),
.B(n_896),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1312),
.Y(n_1422)
);

INVxp33_ASAP7_75t_L g1423 ( 
.A(n_1356),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1360),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1324),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1320),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1323),
.B(n_948),
.C(n_946),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1325),
.Y(n_1428)
);

AND2x2_ASAP7_75t_SL g1429 ( 
.A(n_1333),
.B(n_1250),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1326),
.B(n_977),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1361),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1362),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1328),
.B(n_1186),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1330),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1341),
.A2(n_965),
.B1(n_969),
.B2(n_950),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1363),
.B(n_971),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1366),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1367),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1370),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1373),
.Y(n_1440)
);

INVxp67_ASAP7_75t_L g1441 ( 
.A(n_1374),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1344),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1372),
.B(n_1167),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1331),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1352),
.A2(n_1108),
.B1(n_1192),
.B2(n_1060),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1371),
.Y(n_1446)
);

AND2x6_ASAP7_75t_L g1447 ( 
.A(n_1351),
.B(n_890),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1322),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1346),
.B(n_1126),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1331),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1322),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1346),
.B(n_1128),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_L g1453 ( 
.A(n_1348),
.B(n_972),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1346),
.B(n_989),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1371),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1371),
.B(n_1171),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1346),
.B(n_998),
.Y(n_1457)
);

INVxp33_ASAP7_75t_L g1458 ( 
.A(n_1314),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1346),
.B(n_1006),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1371),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1371),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1314),
.B(n_1007),
.Y(n_1462)
);

INVx4_ASAP7_75t_L g1463 ( 
.A(n_1371),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1346),
.B(n_1014),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1348),
.B(n_1022),
.C(n_1016),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1322),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1346),
.B(n_1034),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1371),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1322),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1371),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1371),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1352),
.A2(n_1108),
.B1(n_1192),
.B2(n_1060),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1331),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1371),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1346),
.B(n_1055),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1371),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1331),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1371),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1371),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1346),
.B(n_1065),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1314),
.B(n_1075),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1346),
.B(n_1079),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1371),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1355),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1322),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1331),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1371),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1365),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1365),
.B(n_1088),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1343),
.B(n_967),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1391),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1413),
.B(n_1105),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1453),
.A2(n_874),
.B(n_862),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1387),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1378),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1454),
.A2(n_901),
.B(n_914),
.C(n_891),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1386),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1403),
.B(n_1107),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1409),
.B(n_1109),
.Y(n_1499)
);

AO22x2_ASAP7_75t_L g1500 ( 
.A1(n_1380),
.A2(n_918),
.B1(n_949),
.B2(n_939),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1398),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1488),
.B(n_1393),
.Y(n_1502)
);

NOR3xp33_ASAP7_75t_L g1503 ( 
.A(n_1405),
.B(n_1123),
.C(n_1113),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1397),
.B(n_1202),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1399),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1449),
.B(n_1137),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1418),
.B(n_1140),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1452),
.B(n_1489),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1444),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1471),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1457),
.B(n_1155),
.Y(n_1512)
);

BUFx4f_ASAP7_75t_L g1513 ( 
.A(n_1395),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1458),
.B(n_1163),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1464),
.B(n_1166),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1390),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1450),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1462),
.B(n_1),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1384),
.B(n_1414),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1481),
.B(n_2),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1467),
.B(n_1182),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1401),
.B(n_954),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1478),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1459),
.A2(n_955),
.B(n_961),
.C(n_960),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1477),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1478),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1394),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1482),
.B(n_1486),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1437),
.B(n_1194),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1388),
.B(n_3),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1400),
.B(n_1465),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1417),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1426),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1470),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1475),
.B(n_974),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_L g1537 ( 
.A(n_1411),
.B(n_993),
.C(n_975),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1480),
.B(n_995),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_L g1539 ( 
.A(n_1377),
.B(n_854),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1455),
.B(n_1474),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_SL g1541 ( 
.A(n_1383),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1392),
.B(n_863),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1404),
.B(n_866),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1385),
.A2(n_1000),
.B1(n_1008),
.B2(n_1002),
.C(n_1001),
.Y(n_1544)
);

OAI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1445),
.A2(n_1015),
.B1(n_1026),
.B2(n_1025),
.C(n_1017),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1434),
.B(n_1188),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1428),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1441),
.B(n_1036),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_SL g1549 ( 
.A(n_1383),
.B(n_882),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1440),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1406),
.B(n_868),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1421),
.B(n_1043),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1423),
.B(n_1044),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1422),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1435),
.B(n_1433),
.Y(n_1555)
);

BUFx5_ASAP7_75t_L g1556 ( 
.A(n_1377),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1484),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1436),
.B(n_869),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1377),
.B(n_1045),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1424),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1431),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1432),
.A2(n_1121),
.B1(n_1129),
.B2(n_1039),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1430),
.B(n_1180),
.Y(n_1563)
);

BUFx8_ASAP7_75t_L g1564 ( 
.A(n_1382),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1407),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1448),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1379),
.B(n_870),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1446),
.B(n_1057),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_L g1569 ( 
.A(n_1490),
.B(n_871),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1438),
.A2(n_1439),
.B1(n_1466),
.B2(n_1451),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1469),
.B(n_1059),
.Y(n_1571)
);

NOR3xp33_ASAP7_75t_L g1572 ( 
.A(n_1427),
.B(n_1073),
.C(n_1070),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1485),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1472),
.B(n_1074),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1476),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1460),
.B(n_877),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1483),
.B(n_1076),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1443),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1415),
.B(n_3),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1419),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1420),
.Y(n_1581)
);

AND2x6_ASAP7_75t_SL g1582 ( 
.A(n_1389),
.B(n_1082),
.Y(n_1582)
);

BUFx5_ASAP7_75t_L g1583 ( 
.A(n_1447),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1381),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1463),
.B(n_878),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1408),
.A2(n_1114),
.B1(n_1116),
.B2(n_1089),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1382),
.B(n_886),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1461),
.B(n_887),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1456),
.Y(n_1589)
);

O2A1O1Ixp5_ASAP7_75t_L g1590 ( 
.A1(n_1396),
.A2(n_1136),
.B(n_1139),
.C(n_1130),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1468),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1410),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1412),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1402),
.B(n_1141),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1447),
.B(n_1142),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1447),
.B(n_1150),
.Y(n_1596)
);

INVxp67_ASAP7_75t_SL g1597 ( 
.A(n_1479),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1425),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1487),
.B(n_894),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1416),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1442),
.B(n_1152),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1429),
.B(n_1157),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1403),
.B(n_898),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1403),
.B(n_899),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1378),
.Y(n_1605)
);

NOR2xp67_ASAP7_75t_L g1606 ( 
.A(n_1397),
.B(n_1176),
.Y(n_1606)
);

AND2x4_ASAP7_75t_SL g1607 ( 
.A(n_1397),
.B(n_1164),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1391),
.A2(n_1170),
.B1(n_1172),
.B2(n_1165),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1413),
.B(n_903),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1458),
.B(n_905),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1391),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1413),
.B(n_907),
.Y(n_1612)
);

NAND2x1_ASAP7_75t_L g1613 ( 
.A(n_1377),
.B(n_917),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1378),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1413),
.B(n_908),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1403),
.B(n_910),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1458),
.B(n_912),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1378),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1413),
.B(n_919),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1378),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1378),
.Y(n_1621)
);

AO22x1_ASAP7_75t_L g1622 ( 
.A1(n_1423),
.A2(n_879),
.B1(n_883),
.B2(n_855),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1391),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1413),
.B(n_922),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1391),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1378),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1401),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1391),
.A2(n_1185),
.B1(n_970),
.B2(n_902),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1403),
.B(n_925),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1378),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1403),
.B(n_926),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1378),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1391),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1413),
.B(n_931),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1413),
.B(n_932),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1484),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1413),
.B(n_933),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1413),
.B(n_934),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1471),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1418),
.A2(n_928),
.B(n_959),
.C(n_911),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1388),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1391),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1413),
.B(n_935),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_L g1644 ( 
.A(n_1488),
.B(n_1098),
.C(n_1027),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1413),
.B(n_937),
.Y(n_1645)
);

AND2x2_ASAP7_75t_SL g1646 ( 
.A(n_1397),
.B(n_1122),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1378),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1403),
.B(n_940),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1401),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1613),
.A2(n_1156),
.B(n_1153),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1491),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1529),
.B(n_941),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1547),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1500),
.A2(n_1160),
.B1(n_1012),
.B2(n_1021),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1494),
.B(n_4),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_5),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1540),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1646),
.A2(n_980),
.B1(n_990),
.B2(n_947),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1513),
.Y(n_1659)
);

AND2x6_ASAP7_75t_L g1660 ( 
.A(n_1578),
.B(n_917),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1509),
.B(n_1199),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1500),
.A2(n_1012),
.B1(n_1021),
.B2(n_917),
.Y(n_1662)
);

BUFx4f_ASAP7_75t_L g1663 ( 
.A(n_1557),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1512),
.B(n_6),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1509),
.B(n_1203),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1639),
.B(n_1205),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1515),
.B(n_6),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1501),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1598),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1505),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1554),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1560),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1510),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1555),
.A2(n_945),
.B1(n_958),
.B2(n_943),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1521),
.B(n_1507),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1636),
.B(n_963),
.C(n_962),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1508),
.B(n_1530),
.Y(n_1677)
);

CKINVDCx8_ASAP7_75t_R g1678 ( 
.A(n_1557),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1517),
.B(n_7),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_SL g1680 ( 
.A(n_1503),
.B(n_992),
.C(n_981),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1541),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1525),
.B(n_7),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1511),
.B(n_8),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1639),
.B(n_1177),
.Y(n_1684)
);

BUFx12f_ASAP7_75t_L g1685 ( 
.A(n_1564),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1561),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1627),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1649),
.B(n_8),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1602),
.A2(n_1021),
.B1(n_1029),
.B2(n_1012),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1607),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1495),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1526),
.B(n_9),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1641),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1611),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_R g1695 ( 
.A(n_1549),
.B(n_968),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1623),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1523),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1575),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1625),
.B(n_1633),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1642),
.B(n_9),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1497),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1533),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1499),
.B(n_10),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1544),
.A2(n_1011),
.B1(n_1032),
.B2(n_987),
.Y(n_1704)
);

NAND2x2_ASAP7_75t_L g1705 ( 
.A(n_1518),
.B(n_10),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1535),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1601),
.B(n_11),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_R g1708 ( 
.A(n_1583),
.B(n_1159),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1492),
.B(n_11),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1527),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1592),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1522),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1519),
.B(n_12),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1531),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1593),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1502),
.B(n_12),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1534),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1550),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1514),
.B(n_973),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1553),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1573),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1556),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1516),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1610),
.A2(n_979),
.B1(n_982),
.B2(n_978),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1577),
.Y(n_1725)
);

BUFx4_ASAP7_75t_SL g1726 ( 
.A(n_1582),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1584),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1617),
.A2(n_984),
.B1(n_986),
.B2(n_983),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1528),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1609),
.B(n_13),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1612),
.B(n_13),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1565),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1506),
.B(n_988),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1615),
.B(n_14),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1589),
.B(n_1029),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1532),
.A2(n_997),
.B1(n_999),
.B2(n_991),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1566),
.Y(n_1737)
);

BUFx4f_ASAP7_75t_L g1738 ( 
.A(n_1594),
.Y(n_1738)
);

NOR2x2_ASAP7_75t_L g1739 ( 
.A(n_1591),
.B(n_1580),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_R g1740 ( 
.A(n_1539),
.B(n_1004),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1579),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1605),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1619),
.B(n_14),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1537),
.B(n_1009),
.C(n_1005),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_L g1745 ( 
.A(n_1556),
.B(n_1013),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1520),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1597),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1624),
.B(n_1020),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1634),
.B(n_15),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1586),
.A2(n_1024),
.B1(n_1030),
.B2(n_1023),
.Y(n_1750)
);

NOR2x2_ASAP7_75t_L g1751 ( 
.A(n_1614),
.B(n_16),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1581),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1556),
.B(n_1184),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1635),
.B(n_16),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1618),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1583),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1620),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1498),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1637),
.B(n_17),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1556),
.B(n_1200),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1504),
.B(n_19),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1621),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1638),
.A2(n_1069),
.B1(n_1086),
.B2(n_1047),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1626),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1630),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1643),
.B(n_19),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1606),
.B(n_1151),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1653),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1671),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1710),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1672),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1720),
.B(n_1645),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1651),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1675),
.B(n_1583),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1659),
.Y(n_1775)
);

BUFx4f_ASAP7_75t_L g1776 ( 
.A(n_1685),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1686),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1687),
.B(n_1568),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1712),
.B(n_1574),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1678),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1747),
.B(n_1583),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1668),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1670),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1673),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1693),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1681),
.B(n_1632),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1663),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1695),
.B(n_1496),
.Y(n_1788)
);

A2O1A1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1719),
.A2(n_1524),
.B(n_1538),
.C(n_1536),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1652),
.B(n_1563),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1691),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1707),
.B(n_1558),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1677),
.B(n_1548),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1694),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1701),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1698),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1714),
.B(n_1552),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1738),
.B(n_1644),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1725),
.B(n_1647),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1715),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1726),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1706),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1715),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1748),
.B(n_1545),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1758),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1704),
.A2(n_1569),
.B1(n_1572),
.B2(n_1628),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1723),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1752),
.B(n_1559),
.Y(n_1808)
);

OR2x4_ASAP7_75t_L g1809 ( 
.A(n_1680),
.B(n_1595),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1711),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1690),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1696),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1764),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1702),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1657),
.B(n_1622),
.Y(n_1815)
);

NOR2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1713),
.B(n_1596),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1735),
.B(n_1543),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1697),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1729),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1746),
.B(n_1542),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1740),
.B(n_1546),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1765),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1699),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1717),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1739),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1658),
.A2(n_1608),
.B1(n_1551),
.B2(n_1604),
.Y(n_1826)
);

AND2x6_ASAP7_75t_SL g1827 ( 
.A(n_1683),
.B(n_1571),
.Y(n_1827)
);

OR2x6_ASAP7_75t_L g1828 ( 
.A(n_1735),
.B(n_1567),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1721),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1664),
.B(n_1493),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1741),
.A2(n_1616),
.B1(n_1629),
.B2(n_1603),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1718),
.B(n_1570),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1764),
.Y(n_1833)
);

AND3x1_ASAP7_75t_SL g1834 ( 
.A(n_1705),
.B(n_20),
.C(n_21),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1669),
.B(n_1587),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1732),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1727),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1716),
.B(n_1631),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1737),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1655),
.B(n_1703),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1688),
.Y(n_1841)
);

BUFx10_ASAP7_75t_L g1842 ( 
.A(n_1733),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1742),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1656),
.B(n_1648),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1755),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1757),
.B(n_1562),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1762),
.B(n_1640),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1679),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1661),
.B(n_1588),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1682),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1665),
.B(n_1576),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1666),
.B(n_1585),
.Y(n_1852)
);

INVxp67_ASAP7_75t_SL g1853 ( 
.A(n_1745),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1660),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1750),
.A2(n_1599),
.B1(n_1031),
.B2(n_1035),
.Y(n_1855)
);

AND2x6_ASAP7_75t_L g1856 ( 
.A(n_1761),
.B(n_1029),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1684),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1692),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1751),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1700),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1676),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1736),
.B(n_20),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1709),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1730),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1731),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1734),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1667),
.B(n_21),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1743),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1749),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1754),
.Y(n_1870)
);

INVxp67_ASAP7_75t_SL g1871 ( 
.A(n_1759),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1724),
.B(n_1033),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1766),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1662),
.B(n_1590),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1660),
.B(n_23),
.Y(n_1875)
);

AOI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1753),
.A2(n_1058),
.B(n_1040),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_SL g1877 ( 
.A(n_1728),
.B(n_1674),
.C(n_1654),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1660),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1708),
.Y(n_1879)
);

INVxp67_ASAP7_75t_L g1880 ( 
.A(n_1767),
.Y(n_1880)
);

AND2x6_ASAP7_75t_L g1881 ( 
.A(n_1722),
.B(n_1058),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1756),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1763),
.B(n_23),
.Y(n_1883)
);

BUFx4f_ASAP7_75t_SL g1884 ( 
.A(n_1760),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1744),
.A2(n_1046),
.B1(n_1048),
.B2(n_1038),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_L g1886 ( 
.A(n_1689),
.B(n_1052),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1650),
.Y(n_1887)
);

INVx5_ASAP7_75t_L g1888 ( 
.A(n_1685),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1671),
.Y(n_1889)
);

BUFx3_ASAP7_75t_L g1890 ( 
.A(n_1659),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1671),
.Y(n_1891)
);

OR2x6_ASAP7_75t_L g1892 ( 
.A(n_1685),
.B(n_1058),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1659),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1659),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1720),
.B(n_24),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1804),
.A2(n_1054),
.B(n_1053),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1823),
.B(n_24),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1895),
.B(n_25),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1789),
.A2(n_1830),
.B(n_1853),
.Y(n_1899)
);

O2A1O1Ixp5_ASAP7_75t_L g1900 ( 
.A1(n_1788),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1779),
.B(n_27),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1802),
.Y(n_1902)
);

INVx5_ASAP7_75t_L g1903 ( 
.A(n_1787),
.Y(n_1903)
);

OAI21x1_ASAP7_75t_L g1904 ( 
.A1(n_1887),
.A2(n_303),
.B(n_302),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1790),
.A2(n_1072),
.B(n_1056),
.Y(n_1905)
);

AO31x2_ASAP7_75t_L g1906 ( 
.A1(n_1878),
.A2(n_305),
.A3(n_307),
.B(n_304),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1768),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1774),
.A2(n_1077),
.B(n_1067),
.Y(n_1908)
);

AOI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1874),
.A2(n_1081),
.B(n_1078),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1769),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1792),
.A2(n_1084),
.B(n_1083),
.Y(n_1911)
);

OAI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1876),
.A2(n_1781),
.B(n_1847),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1773),
.A2(n_309),
.B(n_308),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1872),
.A2(n_1087),
.B(n_1085),
.Y(n_1914)
);

AND3x2_ASAP7_75t_L g1915 ( 
.A(n_1825),
.B(n_1091),
.C(n_1090),
.Y(n_1915)
);

AOI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1870),
.A2(n_1094),
.B(n_1093),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1772),
.B(n_28),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1890),
.B(n_1894),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1858),
.A2(n_1871),
.B(n_1806),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1793),
.B(n_28),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1771),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1797),
.B(n_1796),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1798),
.B(n_29),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1848),
.B(n_30),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1826),
.A2(n_1097),
.B1(n_1100),
.B2(n_1095),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1844),
.A2(n_1101),
.B(n_1096),
.Y(n_1926)
);

NOR2x1p5_ASAP7_75t_L g1927 ( 
.A(n_1780),
.B(n_1158),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1883),
.A2(n_1110),
.B(n_1103),
.Y(n_1928)
);

OAI21x1_ASAP7_75t_L g1929 ( 
.A1(n_1782),
.A2(n_314),
.B(n_311),
.Y(n_1929)
);

OAI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1783),
.A2(n_317),
.B(n_315),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1859),
.B(n_31),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1850),
.B(n_31),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1867),
.A2(n_1111),
.B1(n_1117),
.B2(n_1104),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1860),
.B(n_1118),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1863),
.A2(n_1125),
.B(n_1119),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1864),
.A2(n_1131),
.B(n_1127),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1784),
.A2(n_323),
.B(n_320),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1821),
.B(n_32),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1794),
.A2(n_328),
.B(n_327),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1882),
.B(n_1134),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1893),
.Y(n_1941)
);

AO22x2_ASAP7_75t_L g1942 ( 
.A1(n_1865),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_L g1943 ( 
.A1(n_1812),
.A2(n_330),
.B(n_329),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1814),
.A2(n_335),
.B(n_332),
.Y(n_1944)
);

AOI21x1_ASAP7_75t_SL g1945 ( 
.A1(n_1862),
.A2(n_33),
.B(n_34),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1877),
.A2(n_1145),
.B(n_1135),
.Y(n_1946)
);

AO21x1_ASAP7_75t_L g1947 ( 
.A1(n_1875),
.A2(n_35),
.B(n_36),
.Y(n_1947)
);

AOI21xp33_ASAP7_75t_L g1948 ( 
.A1(n_1838),
.A2(n_1146),
.B(n_1143),
.Y(n_1948)
);

AO31x2_ASAP7_75t_L g1949 ( 
.A1(n_1873),
.A2(n_339),
.A3(n_340),
.B(n_337),
.Y(n_1949)
);

AO21x2_ASAP7_75t_L g1950 ( 
.A1(n_1815),
.A2(n_1149),
.B(n_1147),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1866),
.A2(n_1168),
.B(n_1161),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1829),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1868),
.B(n_35),
.Y(n_1953)
);

NAND2x1_ASAP7_75t_L g1954 ( 
.A(n_1881),
.B(n_343),
.Y(n_1954)
);

AOI221x1_ASAP7_75t_L g1955 ( 
.A1(n_1869),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_1955)
);

OAI21x1_ASAP7_75t_L g1956 ( 
.A1(n_1824),
.A2(n_1832),
.B(n_1854),
.Y(n_1956)
);

AOI211x1_ASAP7_75t_L g1957 ( 
.A1(n_1820),
.A2(n_1840),
.B(n_1808),
.C(n_1834),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1785),
.B(n_38),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1810),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1831),
.A2(n_1173),
.B1(n_1175),
.B2(n_1169),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1836),
.Y(n_1961)
);

AOI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1839),
.A2(n_1179),
.B(n_1174),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1770),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1816),
.B(n_40),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1842),
.B(n_1778),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1818),
.B(n_41),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1805),
.B(n_1775),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1827),
.B(n_41),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1843),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1893),
.B(n_1861),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1800),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1845),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1884),
.B(n_42),
.Y(n_1973)
);

A2O1A1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1880),
.A2(n_1189),
.B(n_1196),
.C(n_1181),
.Y(n_1974)
);

OA21x2_ASAP7_75t_L g1975 ( 
.A1(n_1846),
.A2(n_42),
.B(n_43),
.Y(n_1975)
);

AO31x2_ASAP7_75t_L g1976 ( 
.A1(n_1791),
.A2(n_345),
.A3(n_346),
.B(n_344),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1941),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1961),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1952),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1902),
.B(n_1888),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1907),
.Y(n_1981)
);

OR2x6_ASAP7_75t_L g1982 ( 
.A(n_1965),
.B(n_1892),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1917),
.A2(n_1809),
.B1(n_1857),
.B2(n_1817),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1973),
.B(n_1801),
.Y(n_1984)
);

NOR2x1p5_ASAP7_75t_L g1985 ( 
.A(n_1968),
.B(n_1938),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1941),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1922),
.B(n_1777),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1918),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1959),
.Y(n_1989)
);

O2A1O1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1896),
.A2(n_1828),
.B(n_1817),
.C(n_1851),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1971),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1963),
.B(n_1889),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1925),
.A2(n_1828),
.B1(n_1852),
.B2(n_1849),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1897),
.B(n_1891),
.Y(n_1994)
);

A2O1A1Ixp33_ASAP7_75t_SL g1995 ( 
.A1(n_1967),
.A2(n_1879),
.B(n_1885),
.C(n_1855),
.Y(n_1995)
);

A2O1A1Ixp33_ASAP7_75t_L g1996 ( 
.A1(n_1919),
.A2(n_1835),
.B(n_1811),
.C(n_1886),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1972),
.B(n_1969),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1910),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1942),
.A2(n_1799),
.B1(n_1856),
.B2(n_1845),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1957),
.A2(n_1776),
.B1(n_1892),
.B2(n_1888),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1971),
.B(n_1803),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1903),
.Y(n_2002)
);

BUFx12f_ASAP7_75t_L g2003 ( 
.A(n_1927),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1903),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_SL g2005 ( 
.A(n_1970),
.B(n_1800),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1905),
.A2(n_1841),
.B1(n_1837),
.B2(n_1813),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1899),
.A2(n_1881),
.B(n_1807),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1966),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1923),
.B(n_1841),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1921),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1901),
.B(n_1833),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1946),
.A2(n_1881),
.B(n_1819),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1956),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1915),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1975),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1942),
.Y(n_2016)
);

OAI21x1_ASAP7_75t_L g2017 ( 
.A1(n_1912),
.A2(n_1822),
.B(n_1795),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1954),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1898),
.B(n_1833),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1920),
.A2(n_1786),
.B1(n_1856),
.B2(n_46),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1964),
.B(n_1856),
.Y(n_2021)
);

O2A1O1Ixp5_ASAP7_75t_SL g2022 ( 
.A1(n_1934),
.A2(n_47),
.B(n_44),
.C(n_45),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_1958),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1931),
.B(n_44),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1940),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1981),
.B(n_1989),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1986),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1979),
.Y(n_2028)
);

BUFx4_ASAP7_75t_SL g2029 ( 
.A(n_2023),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2019),
.B(n_1953),
.Y(n_2030)
);

A2O1A1Ixp33_ASAP7_75t_L g2031 ( 
.A1(n_2020),
.A2(n_1914),
.B(n_1928),
.C(n_1948),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1997),
.B(n_1924),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1978),
.B(n_1992),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1998),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1983),
.B(n_1947),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1980),
.B(n_1932),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_2003),
.Y(n_2037)
);

O2A1O1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_1995),
.A2(n_1960),
.B(n_1933),
.C(n_1951),
.Y(n_2038)
);

A2O1A1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1990),
.A2(n_1996),
.B(n_1985),
.C(n_1900),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1977),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1988),
.B(n_1906),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_2008),
.B(n_1916),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1994),
.B(n_1950),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_2007),
.A2(n_1955),
.B(n_1929),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2009),
.B(n_1913),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2010),
.Y(n_2046)
);

A2O1A1Ixp33_ASAP7_75t_L g2047 ( 
.A1(n_2024),
.A2(n_1936),
.B(n_1935),
.C(n_1926),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2011),
.B(n_1930),
.Y(n_2048)
);

A2O1A1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_2016),
.A2(n_1974),
.B(n_1911),
.C(n_1939),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1991),
.B(n_1937),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1977),
.B(n_1943),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1987),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2000),
.A2(n_1909),
.B1(n_1962),
.B2(n_1945),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2004),
.B(n_45),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1999),
.A2(n_1908),
.B1(n_1944),
.B2(n_1906),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2012),
.A2(n_1904),
.B(n_1949),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2005),
.B(n_1949),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2015),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2001),
.B(n_48),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_2002),
.B(n_1976),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_2013),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2017),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_2002),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_1982),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1982),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2025),
.B(n_48),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2021),
.B(n_49),
.Y(n_2067)
);

A2O1A1Ixp33_ASAP7_75t_L g2068 ( 
.A1(n_1993),
.A2(n_1976),
.B(n_51),
.C(n_49),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2006),
.B(n_50),
.Y(n_2069)
);

O2A1O1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1984),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_2070)
);

O2A1O1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_2018),
.A2(n_2022),
.B(n_54),
.C(n_52),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2014),
.A2(n_53),
.B(n_54),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2014),
.B(n_347),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1979),
.Y(n_2074)
);

A2O1A1Ixp33_ASAP7_75t_L g2075 ( 
.A1(n_2020),
.A2(n_56),
.B(n_53),
.C(n_55),
.Y(n_2075)
);

OAI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2020),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1981),
.B(n_58),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2028),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_2037),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2074),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2046),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2034),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_2026),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2058),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2061),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2033),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2052),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2043),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2026),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_2029),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2030),
.B(n_59),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2041),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2062),
.Y(n_2093)
);

INVx4_ASAP7_75t_L g2094 ( 
.A(n_2040),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2032),
.B(n_60),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_2045),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_2048),
.B(n_2065),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2077),
.B(n_61),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2050),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2057),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2064),
.Y(n_2101)
);

OR2x6_ASAP7_75t_L g2102 ( 
.A(n_2036),
.B(n_61),
.Y(n_2102)
);

INVx4_ASAP7_75t_SL g2103 ( 
.A(n_2073),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2063),
.B(n_62),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2060),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2051),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2035),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2067),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2054),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2066),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2069),
.Y(n_2111)
);

BUFx3_ASAP7_75t_L g2112 ( 
.A(n_2027),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2059),
.B(n_63),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2042),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2039),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2056),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2055),
.Y(n_2117)
);

INVx3_ASAP7_75t_L g2118 ( 
.A(n_2049),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_2068),
.B(n_2072),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_2044),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2053),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2075),
.B(n_65),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2076),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2070),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2047),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_2038),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_2031),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2071),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2028),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_2056),
.A2(n_65),
.B(n_66),
.Y(n_2130)
);

OAI221xp5_ASAP7_75t_L g2131 ( 
.A1(n_2039),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.C(n_70),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2035),
.A2(n_71),
.B1(n_67),
.B2(n_68),
.Y(n_2132)
);

OAI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_2039),
.A2(n_71),
.B(n_72),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_2061),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2028),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2028),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2028),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2028),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2028),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2028),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_2027),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_2026),
.Y(n_2142)
);

OR2x6_ASAP7_75t_L g2143 ( 
.A(n_2064),
.B(n_72),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2028),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_L g2145 ( 
.A1(n_2056),
.A2(n_73),
.B(n_74),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2033),
.B(n_73),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2028),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2028),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2028),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2028),
.Y(n_2150)
);

NOR2x1_ASAP7_75t_R g2151 ( 
.A(n_2037),
.B(n_74),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_2061),
.Y(n_2152)
);

OAI21x1_ASAP7_75t_L g2153 ( 
.A1(n_2056),
.A2(n_75),
.B(n_76),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2028),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_2097),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2083),
.B(n_75),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2085),
.B(n_76),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_2142),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2096),
.B(n_77),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2089),
.B(n_77),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2134),
.B(n_78),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_2079),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2152),
.B(n_2101),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2099),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2087),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2106),
.B(n_78),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2078),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2120),
.B(n_79),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_2127),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2126),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2084),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_2090),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2129),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2141),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_2114),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_2111),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2100),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2080),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2135),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2136),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2086),
.B(n_83),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2117),
.Y(n_2182)
);

AND2x4_ASAP7_75t_L g2183 ( 
.A(n_2092),
.B(n_2108),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2125),
.B(n_83),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_2112),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2138),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2126),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_2094),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2137),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_2109),
.Y(n_2190)
);

AOI22xp33_ASAP7_75t_L g2191 ( 
.A1(n_2118),
.A2(n_87),
.B1(n_84),
.B2(n_85),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2082),
.B(n_88),
.Y(n_2192)
);

INVx2_ASAP7_75t_SL g2193 ( 
.A(n_2091),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2148),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2154),
.Y(n_2195)
);

BUFx8_ASAP7_75t_SL g2196 ( 
.A(n_2143),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_2110),
.B(n_89),
.Y(n_2197)
);

BUFx2_ASAP7_75t_L g2198 ( 
.A(n_2121),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2088),
.B(n_2095),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_2104),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_2102),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2139),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2093),
.B(n_89),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2105),
.B(n_90),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2140),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2116),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2115),
.B(n_90),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2131),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_2102),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2144),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2113),
.B(n_91),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2147),
.Y(n_2212)
);

NAND3xp33_ASAP7_75t_L g2213 ( 
.A(n_2133),
.B(n_92),
.C(n_93),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_2143),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2146),
.B(n_94),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2149),
.B(n_94),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_2150),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2098),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2123),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2103),
.B(n_96),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2081),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2103),
.B(n_96),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2124),
.B(n_97),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2130),
.Y(n_2224)
);

OR2x2_ASAP7_75t_L g2225 ( 
.A(n_2128),
.B(n_2145),
.Y(n_2225)
);

OAI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_2107),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2153),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_2119),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2122),
.B(n_98),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2151),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2132),
.B(n_99),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2085),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2085),
.B(n_101),
.Y(n_2233)
);

INVx4_ASAP7_75t_L g2234 ( 
.A(n_2141),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2087),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2083),
.B(n_101),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2083),
.B(n_102),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_2085),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2085),
.B(n_103),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2083),
.B(n_103),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2085),
.B(n_104),
.Y(n_2241)
);

INVx2_ASAP7_75t_SL g2242 ( 
.A(n_2090),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2083),
.B(n_104),
.Y(n_2243)
);

AO31x2_ASAP7_75t_L g2244 ( 
.A1(n_2114),
.A2(n_107),
.A3(n_105),
.B(n_106),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2083),
.B(n_105),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2087),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_2126),
.B(n_106),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2083),
.B(n_107),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2099),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2083),
.B(n_108),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2083),
.B(n_109),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2087),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2083),
.B(n_109),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2225),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2167),
.Y(n_2255)
);

OAI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2228),
.A2(n_112),
.B1(n_113),
.B2(n_111),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2219),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2177),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_2238),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_2234),
.B(n_2184),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2198),
.B(n_2155),
.Y(n_2261)
);

INVx4_ASAP7_75t_L g2262 ( 
.A(n_2188),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_2182),
.B(n_2238),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2173),
.Y(n_2264)
);

BUFx3_ASAP7_75t_L g2265 ( 
.A(n_2196),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2224),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2190),
.B(n_110),
.Y(n_2267)
);

OAI222xp33_ASAP7_75t_L g2268 ( 
.A1(n_2224),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.C1(n_112),
.C2(n_114),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2171),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2178),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2206),
.B(n_111),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2180),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2168),
.B(n_114),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2179),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_2172),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2163),
.B(n_2193),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2186),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2232),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2194),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2195),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2165),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2158),
.B(n_115),
.Y(n_2282)
);

OR2x2_ASAP7_75t_L g2283 ( 
.A(n_2175),
.B(n_116),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2159),
.B(n_117),
.Y(n_2284)
);

AO21x2_ASAP7_75t_L g2285 ( 
.A1(n_2192),
.A2(n_117),
.B(n_118),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2189),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2235),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2246),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2205),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2199),
.B(n_119),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2162),
.B(n_120),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2200),
.B(n_120),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2201),
.B(n_121),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_L g2294 ( 
.A1(n_2213),
.A2(n_124),
.B1(n_126),
.B2(n_122),
.C1(n_123),
.C2(n_125),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2212),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2218),
.B(n_123),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2227),
.Y(n_2297)
);

INVx4_ASAP7_75t_L g2298 ( 
.A(n_2230),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2209),
.B(n_124),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2242),
.B(n_125),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2166),
.B(n_127),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2161),
.B(n_127),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2185),
.B(n_128),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2221),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2157),
.B(n_128),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2176),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2164),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2233),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2249),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2252),
.Y(n_2310)
);

AOI211xp5_ASAP7_75t_L g2311 ( 
.A1(n_2247),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2202),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2183),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2217),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2210),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2203),
.B(n_129),
.Y(n_2316)
);

AND2x4_ASAP7_75t_SL g2317 ( 
.A(n_2220),
.B(n_131),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_2222),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2181),
.B(n_132),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2216),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2239),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2197),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2241),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2160),
.B(n_132),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2207),
.B(n_2223),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2156),
.B(n_133),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2236),
.B(n_133),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2237),
.B(n_134),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2244),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2244),
.Y(n_2330)
);

AND2x4_ASAP7_75t_SL g2331 ( 
.A(n_2240),
.B(n_135),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2204),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2243),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2245),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2248),
.Y(n_2335)
);

HB1xp67_ASAP7_75t_L g2336 ( 
.A(n_2250),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2251),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2253),
.B(n_135),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2214),
.B(n_136),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2211),
.B(n_136),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2229),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_2215),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2208),
.B(n_137),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2231),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2174),
.Y(n_2345)
);

INVxp67_ASAP7_75t_SL g2346 ( 
.A(n_2169),
.Y(n_2346)
);

AND2x4_ASAP7_75t_SL g2347 ( 
.A(n_2170),
.B(n_137),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2226),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2191),
.B(n_138),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2187),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2167),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_2219),
.B(n_138),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2198),
.B(n_139),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_2196),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2182),
.B(n_139),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2182),
.B(n_140),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2182),
.B(n_141),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2167),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2182),
.B(n_141),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2167),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2172),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2198),
.B(n_142),
.Y(n_2362)
);

AOI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2213),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2238),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2198),
.B(n_143),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2198),
.B(n_144),
.Y(n_2366)
);

AO21x1_ASAP7_75t_L g2367 ( 
.A1(n_2168),
.A2(n_145),
.B(n_146),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2198),
.B(n_145),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2198),
.B(n_146),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2167),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2225),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2167),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2198),
.B(n_147),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2257),
.Y(n_2374)
);

OR2x2_ASAP7_75t_L g2375 ( 
.A(n_2263),
.B(n_148),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2361),
.B(n_148),
.Y(n_2376)
);

INVx1_ASAP7_75t_SL g2377 ( 
.A(n_2265),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2255),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2342),
.B(n_149),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2264),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2278),
.B(n_149),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2330),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2272),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2314),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2308),
.B(n_150),
.Y(n_2385)
);

NOR2xp67_ASAP7_75t_SL g2386 ( 
.A(n_2354),
.B(n_150),
.Y(n_2386)
);

BUFx2_ASAP7_75t_L g2387 ( 
.A(n_2275),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2277),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2313),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2279),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2261),
.B(n_151),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_2276),
.B(n_151),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_2298),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2334),
.B(n_152),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2321),
.B(n_154),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2280),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2259),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2341),
.B(n_155),
.Y(n_2398)
);

HB1xp67_ASAP7_75t_L g2399 ( 
.A(n_2364),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2351),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2271),
.B(n_155),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2297),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2358),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2355),
.B(n_157),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2323),
.B(n_157),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2360),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2306),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2370),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2372),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2356),
.B(n_158),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2329),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2270),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2336),
.B(n_158),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2359),
.B(n_2285),
.Y(n_2414)
);

AND2x4_ASAP7_75t_L g2415 ( 
.A(n_2352),
.B(n_159),
.Y(n_2415)
);

OR2x2_ASAP7_75t_L g2416 ( 
.A(n_2254),
.B(n_2371),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2281),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2353),
.B(n_159),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2290),
.B(n_160),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2362),
.B(n_160),
.Y(n_2420)
);

OR2x2_ASAP7_75t_L g2421 ( 
.A(n_2357),
.B(n_161),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2287),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2365),
.B(n_161),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2288),
.Y(n_2424)
);

BUFx2_ASAP7_75t_SL g2425 ( 
.A(n_2299),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2274),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_2266),
.Y(n_2427)
);

NAND2x1_ASAP7_75t_L g2428 ( 
.A(n_2373),
.B(n_162),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2286),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2289),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_2299),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2366),
.B(n_162),
.Y(n_2432)
);

NOR2x1_ASAP7_75t_SL g2433 ( 
.A(n_2283),
.B(n_163),
.Y(n_2433)
);

HB1xp67_ASAP7_75t_L g2434 ( 
.A(n_2348),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2291),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2368),
.B(n_163),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2310),
.B(n_164),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2312),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2315),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2258),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2369),
.B(n_164),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2282),
.B(n_165),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2345),
.Y(n_2443)
);

AND2x4_ASAP7_75t_L g2444 ( 
.A(n_2337),
.B(n_165),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2318),
.B(n_166),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2318),
.B(n_166),
.Y(n_2446)
);

BUFx2_ASAP7_75t_L g2447 ( 
.A(n_2262),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2267),
.B(n_167),
.Y(n_2448)
);

NAND2x1p5_ASAP7_75t_L g2449 ( 
.A(n_2292),
.B(n_167),
.Y(n_2449)
);

BUFx3_ASAP7_75t_L g2450 ( 
.A(n_2317),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2367),
.B(n_2296),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2260),
.B(n_168),
.Y(n_2452)
);

INVx3_ASAP7_75t_L g2453 ( 
.A(n_2331),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2344),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2332),
.B(n_168),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2295),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2333),
.B(n_2335),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2339),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2304),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2300),
.B(n_2293),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2269),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2320),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2325),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2303),
.B(n_169),
.Y(n_2464)
);

INVxp67_ASAP7_75t_SL g2465 ( 
.A(n_2346),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2301),
.B(n_170),
.Y(n_2466)
);

NOR2xp67_ASAP7_75t_L g2467 ( 
.A(n_2305),
.B(n_171),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2322),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2307),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2309),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2350),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2340),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2273),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2316),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2302),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2324),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2284),
.B(n_171),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2319),
.B(n_172),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2326),
.B(n_172),
.Y(n_2479)
);

NAND4xp25_ASAP7_75t_L g2480 ( 
.A(n_2294),
.B(n_175),
.C(n_173),
.D(n_174),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2327),
.Y(n_2481)
);

INVx2_ASAP7_75t_SL g2482 ( 
.A(n_2328),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2338),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2343),
.Y(n_2484)
);

INVxp67_ASAP7_75t_SL g2485 ( 
.A(n_2311),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2256),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2363),
.B(n_173),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2268),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2349),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2347),
.B(n_174),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2255),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2342),
.B(n_176),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2255),
.Y(n_2493)
);

OR2x2_ASAP7_75t_L g2494 ( 
.A(n_2263),
.B(n_176),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2257),
.Y(n_2495)
);

HB1xp67_ASAP7_75t_L g2496 ( 
.A(n_2278),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2342),
.B(n_177),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2278),
.Y(n_2498)
);

OR2x2_ASAP7_75t_L g2499 ( 
.A(n_2263),
.B(n_177),
.Y(n_2499)
);

NAND2x1p5_ASAP7_75t_L g2500 ( 
.A(n_2352),
.B(n_178),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2255),
.Y(n_2501)
);

NOR2xp67_ASAP7_75t_L g2502 ( 
.A(n_2263),
.B(n_178),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2342),
.B(n_179),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2342),
.B(n_179),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2257),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2255),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2261),
.B(n_180),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2261),
.B(n_181),
.Y(n_2508)
);

INVxp67_ASAP7_75t_SL g2509 ( 
.A(n_2367),
.Y(n_2509)
);

INVx3_ASAP7_75t_L g2510 ( 
.A(n_2265),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2263),
.B(n_181),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2257),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2257),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2261),
.B(n_182),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2265),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2257),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2261),
.B(n_182),
.Y(n_2517)
);

AND2x4_ASAP7_75t_SL g2518 ( 
.A(n_2361),
.B(n_183),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2261),
.B(n_184),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2361),
.B(n_185),
.Y(n_2520)
);

BUFx6f_ASAP7_75t_SL g2521 ( 
.A(n_2265),
.Y(n_2521)
);

INVxp67_ASAP7_75t_SL g2522 ( 
.A(n_2367),
.Y(n_2522)
);

AND2x4_ASAP7_75t_L g2523 ( 
.A(n_2361),
.B(n_185),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2342),
.B(n_186),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2342),
.B(n_186),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2261),
.B(n_187),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2342),
.B(n_188),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2255),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2255),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2261),
.B(n_188),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2255),
.Y(n_2531)
);

OR2x2_ASAP7_75t_L g2532 ( 
.A(n_2263),
.B(n_189),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2342),
.B(n_189),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2263),
.B(n_190),
.Y(n_2534)
);

INVxp67_ASAP7_75t_SL g2535 ( 
.A(n_2367),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2342),
.B(n_190),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2257),
.Y(n_2537)
);

AND3x1_ASAP7_75t_L g2538 ( 
.A(n_2361),
.B(n_191),
.C(n_192),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2255),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_2265),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_2265),
.Y(n_2541)
);

BUFx12f_ASAP7_75t_L g2542 ( 
.A(n_2299),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2257),
.Y(n_2543)
);

HB1xp67_ASAP7_75t_L g2544 ( 
.A(n_2443),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2393),
.B(n_191),
.Y(n_2545)
);

OA21x2_ASAP7_75t_L g2546 ( 
.A1(n_2465),
.A2(n_193),
.B(n_194),
.Y(n_2546)
);

OAI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2509),
.A2(n_203),
.B1(n_211),
.B2(n_193),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2496),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2541),
.Y(n_2549)
);

OAI211xp5_ASAP7_75t_L g2550 ( 
.A1(n_2522),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2535),
.B(n_197),
.Y(n_2551)
);

NAND4xp25_ASAP7_75t_L g2552 ( 
.A(n_2387),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2498),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2411),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2378),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2484),
.B(n_199),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2540),
.Y(n_2557)
);

AOI21x1_ASAP7_75t_L g2558 ( 
.A1(n_2451),
.A2(n_200),
.B(n_201),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2472),
.Y(n_2559)
);

AOI221xp5_ASAP7_75t_L g2560 ( 
.A1(n_2488),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_2560)
);

AOI31xp33_ASAP7_75t_L g2561 ( 
.A1(n_2485),
.A2(n_211),
.A3(n_219),
.B(n_202),
.Y(n_2561)
);

OA21x2_ASAP7_75t_L g2562 ( 
.A1(n_2414),
.A2(n_204),
.B(n_205),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2380),
.Y(n_2563)
);

BUFx2_ASAP7_75t_L g2564 ( 
.A(n_2510),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2457),
.B(n_206),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2458),
.Y(n_2566)
);

AOI221xp5_ASAP7_75t_L g2567 ( 
.A1(n_2480),
.A2(n_2538),
.B1(n_2487),
.B2(n_2486),
.C(n_2437),
.Y(n_2567)
);

BUFx2_ASAP7_75t_L g2568 ( 
.A(n_2542),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2431),
.B(n_207),
.Y(n_2569)
);

HB1xp67_ASAP7_75t_L g2570 ( 
.A(n_2397),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2476),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2383),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2388),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2460),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2515),
.B(n_207),
.Y(n_2575)
);

BUFx3_ASAP7_75t_L g2576 ( 
.A(n_2541),
.Y(n_2576)
);

INVx5_ASAP7_75t_L g2577 ( 
.A(n_2447),
.Y(n_2577)
);

OAI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2502),
.A2(n_208),
.B(n_209),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2390),
.Y(n_2579)
);

OAI31xp33_ASAP7_75t_L g2580 ( 
.A1(n_2489),
.A2(n_212),
.A3(n_209),
.B(n_210),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2471),
.A2(n_213),
.B1(n_210),
.B2(n_212),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2433),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2399),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2396),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2400),
.Y(n_2585)
);

AOI222xp33_ASAP7_75t_L g2586 ( 
.A1(n_2467),
.A2(n_237),
.B1(n_221),
.B2(n_245),
.C1(n_229),
.C2(n_213),
.Y(n_2586)
);

NOR3xp33_ASAP7_75t_SL g2587 ( 
.A(n_2445),
.B(n_214),
.C(n_215),
.Y(n_2587)
);

AO21x2_ASAP7_75t_L g2588 ( 
.A1(n_2381),
.A2(n_214),
.B(n_216),
.Y(n_2588)
);

INVx3_ASAP7_75t_L g2589 ( 
.A(n_2521),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2463),
.B(n_2434),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2473),
.B(n_216),
.Y(n_2591)
);

AO21x2_ASAP7_75t_L g2592 ( 
.A1(n_2385),
.A2(n_217),
.B(n_218),
.Y(n_2592)
);

AND2x4_ASAP7_75t_SL g2593 ( 
.A(n_2435),
.B(n_217),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2482),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2391),
.B(n_218),
.Y(n_2595)
);

OAI31xp33_ASAP7_75t_SL g2596 ( 
.A1(n_2446),
.A2(n_221),
.A3(n_219),
.B(n_220),
.Y(n_2596)
);

AO21x2_ASAP7_75t_L g2597 ( 
.A1(n_2379),
.A2(n_220),
.B(n_222),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2374),
.B(n_222),
.Y(n_2598)
);

AOI221xp5_ASAP7_75t_L g2599 ( 
.A1(n_2398),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.C(n_226),
.Y(n_2599)
);

AND2x2_ASAP7_75t_SL g2600 ( 
.A(n_2435),
.B(n_224),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2403),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2450),
.Y(n_2602)
);

AND2x4_ASAP7_75t_SL g2603 ( 
.A(n_2453),
.B(n_226),
.Y(n_2603)
);

INVx5_ASAP7_75t_L g2604 ( 
.A(n_2413),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2382),
.Y(n_2605)
);

AO21x2_ASAP7_75t_L g2606 ( 
.A1(n_2492),
.A2(n_227),
.B(n_228),
.Y(n_2606)
);

NAND3xp33_ASAP7_75t_L g2607 ( 
.A(n_2427),
.B(n_227),
.C(n_228),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2407),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2416),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2406),
.Y(n_2610)
);

OA21x2_ASAP7_75t_L g2611 ( 
.A1(n_2495),
.A2(n_229),
.B(n_230),
.Y(n_2611)
);

AO21x2_ASAP7_75t_L g2612 ( 
.A1(n_2497),
.A2(n_230),
.B(n_231),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2425),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2375),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2505),
.B(n_232),
.Y(n_2615)
);

OAI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2494),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2616)
);

NAND4xp25_ASAP7_75t_SL g2617 ( 
.A(n_2377),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2507),
.B(n_236),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2408),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2409),
.Y(n_2620)
);

OAI31xp33_ASAP7_75t_SL g2621 ( 
.A1(n_2418),
.A2(n_240),
.A3(n_238),
.B(n_239),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_2512),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2508),
.B(n_238),
.Y(n_2623)
);

AOI31xp33_ASAP7_75t_SL g2624 ( 
.A1(n_2513),
.A2(n_241),
.A3(n_239),
.B(n_240),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2491),
.Y(n_2625)
);

OAI211xp5_ASAP7_75t_L g2626 ( 
.A1(n_2428),
.A2(n_2499),
.B(n_2532),
.C(n_2511),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2516),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2493),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2501),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2389),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_SL g2631 ( 
.A1(n_2395),
.A2(n_246),
.B1(n_243),
.B2(n_244),
.Y(n_2631)
);

BUFx2_ASAP7_75t_L g2632 ( 
.A(n_2537),
.Y(n_2632)
);

AOI221xp5_ASAP7_75t_L g2633 ( 
.A1(n_2478),
.A2(n_247),
.B1(n_244),
.B2(n_246),
.C(n_248),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2506),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2528),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2529),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2543),
.B(n_249),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2534),
.Y(n_2638)
);

NAND3xp33_ASAP7_75t_L g2639 ( 
.A(n_2384),
.B(n_250),
.C(n_251),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2468),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2531),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2539),
.Y(n_2642)
);

AO21x2_ASAP7_75t_L g2643 ( 
.A1(n_2536),
.A2(n_250),
.B(n_251),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2417),
.Y(n_2644)
);

OR2x2_ASAP7_75t_L g2645 ( 
.A(n_2474),
.B(n_252),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2514),
.B(n_252),
.Y(n_2646)
);

AOI33xp33_ASAP7_75t_L g2647 ( 
.A1(n_2475),
.A2(n_2483),
.A3(n_2481),
.B1(n_2477),
.B2(n_2479),
.B3(n_2423),
.Y(n_2647)
);

AOI21x1_ASAP7_75t_L g2648 ( 
.A1(n_2517),
.A2(n_253),
.B(n_254),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2394),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2422),
.Y(n_2650)
);

NAND4xp25_ASAP7_75t_L g2651 ( 
.A(n_2519),
.B(n_255),
.C(n_253),
.D(n_254),
.Y(n_2651)
);

AO21x2_ASAP7_75t_L g2652 ( 
.A1(n_2533),
.A2(n_255),
.B(n_256),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2392),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2424),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2405),
.B(n_259),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2526),
.B(n_259),
.Y(n_2656)
);

BUFx6f_ASAP7_75t_L g2657 ( 
.A(n_2490),
.Y(n_2657)
);

INVx4_ASAP7_75t_L g2658 ( 
.A(n_2376),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2438),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2439),
.Y(n_2660)
);

INVx3_ASAP7_75t_L g2661 ( 
.A(n_2520),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2454),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2462),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2503),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2504),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2524),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2544),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2557),
.B(n_2530),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2546),
.A2(n_2455),
.B1(n_2444),
.B2(n_2440),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2638),
.B(n_2466),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2548),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2553),
.Y(n_2672)
);

INVxp67_ASAP7_75t_SL g2673 ( 
.A(n_2576),
.Y(n_2673)
);

AOI21xp33_ASAP7_75t_SL g2674 ( 
.A1(n_2561),
.A2(n_2500),
.B(n_2449),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2564),
.B(n_2452),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2570),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2657),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2568),
.B(n_2523),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2583),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2554),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2555),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2589),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2602),
.B(n_2420),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2647),
.B(n_2525),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2563),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2572),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2604),
.B(n_2415),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2657),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2573),
.Y(n_2689)
);

OR2x2_ASAP7_75t_L g2690 ( 
.A(n_2590),
.B(n_2527),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2614),
.B(n_2432),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2577),
.B(n_2436),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2579),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2584),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2585),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2601),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2577),
.B(n_2441),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2549),
.B(n_2518),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2562),
.B(n_2442),
.Y(n_2699)
);

OR2x6_ASAP7_75t_L g2700 ( 
.A(n_2551),
.B(n_2575),
.Y(n_2700)
);

OR2x2_ASAP7_75t_L g2701 ( 
.A(n_2664),
.B(n_2419),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2604),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2658),
.B(n_2464),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2611),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2610),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2665),
.B(n_2421),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2619),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2620),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2625),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2574),
.B(n_2386),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2666),
.B(n_2401),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2661),
.B(n_2448),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2649),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2628),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2582),
.B(n_2404),
.Y(n_2715)
);

OR2x2_ASAP7_75t_L g2716 ( 
.A(n_2571),
.B(n_2594),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2662),
.B(n_2410),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2603),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2629),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2566),
.B(n_2469),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2597),
.B(n_2412),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2634),
.Y(n_2722)
);

AND2x4_ASAP7_75t_L g2723 ( 
.A(n_2569),
.B(n_2426),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2635),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2636),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2565),
.B(n_2470),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2682),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2667),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2692),
.Y(n_2729)
);

OR2x2_ASAP7_75t_L g2730 ( 
.A(n_2670),
.B(n_2559),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2697),
.B(n_2545),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2726),
.B(n_2621),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2671),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2668),
.B(n_2606),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2683),
.B(n_2675),
.Y(n_2735)
);

OAI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2684),
.A2(n_2626),
.B1(n_2567),
.B2(n_2607),
.Y(n_2736)
);

OR2x6_ASAP7_75t_L g2737 ( 
.A(n_2702),
.B(n_2655),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2678),
.B(n_2641),
.Y(n_2738)
);

NAND2x1_ASAP7_75t_L g2739 ( 
.A(n_2703),
.B(n_2642),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2673),
.B(n_2644),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2699),
.B(n_2612),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2672),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2676),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2679),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2691),
.B(n_2643),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2700),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2700),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2701),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2718),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2698),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_SL g2751 ( 
.A(n_2712),
.B(n_2600),
.Y(n_2751)
);

INVxp67_ASAP7_75t_L g2752 ( 
.A(n_2687),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2710),
.B(n_2650),
.Y(n_2753)
);

NAND2x1p5_ASAP7_75t_L g2754 ( 
.A(n_2677),
.B(n_2595),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2706),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2717),
.B(n_2663),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2713),
.B(n_2654),
.Y(n_2757)
);

OR2x2_ASAP7_75t_L g2758 ( 
.A(n_2711),
.B(n_2659),
.Y(n_2758)
);

AND2x2_ASAP7_75t_SL g2759 ( 
.A(n_2731),
.B(n_2596),
.Y(n_2759)
);

AND2x4_ASAP7_75t_L g2760 ( 
.A(n_2727),
.B(n_2688),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2750),
.B(n_2674),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2754),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2735),
.B(n_2690),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2737),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2758),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2738),
.B(n_2715),
.Y(n_2766)
);

OAI21xp5_ASAP7_75t_SL g2767 ( 
.A1(n_2736),
.A2(n_2552),
.B(n_2550),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2740),
.B(n_2652),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2756),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2737),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2751),
.B(n_2732),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2752),
.B(n_2645),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2749),
.B(n_2720),
.Y(n_2773)
);

OR2x6_ASAP7_75t_L g2774 ( 
.A(n_2746),
.B(n_2716),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2748),
.Y(n_2775)
);

INVx4_ASAP7_75t_L g2776 ( 
.A(n_2729),
.Y(n_2776)
);

OR2x2_ASAP7_75t_L g2777 ( 
.A(n_2755),
.B(n_2734),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2728),
.Y(n_2778)
);

NAND2x1p5_ASAP7_75t_L g2779 ( 
.A(n_2760),
.B(n_2747),
.Y(n_2779)
);

NAND4xp25_ASAP7_75t_L g2780 ( 
.A(n_2761),
.B(n_2730),
.C(n_2742),
.D(n_2733),
.Y(n_2780)
);

AND4x1_ASAP7_75t_L g2781 ( 
.A(n_2771),
.B(n_2633),
.C(n_2587),
.D(n_2560),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2774),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2774),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2773),
.Y(n_2784)
);

INVx4_ASAP7_75t_L g2785 ( 
.A(n_2776),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2763),
.B(n_2753),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2759),
.B(n_2669),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2765),
.B(n_2743),
.Y(n_2788)
);

INVx1_ASAP7_75t_SL g2789 ( 
.A(n_2786),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2784),
.Y(n_2790)
);

OAI21xp33_ASAP7_75t_SL g2791 ( 
.A1(n_2780),
.A2(n_2766),
.B(n_2769),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2779),
.Y(n_2792)
);

OAI221xp5_ASAP7_75t_L g2793 ( 
.A1(n_2787),
.A2(n_2767),
.B1(n_2741),
.B2(n_2745),
.C(n_2768),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2782),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2783),
.Y(n_2795)
);

AOI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2785),
.A2(n_2739),
.B(n_2772),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2788),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2789),
.B(n_2764),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2797),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2792),
.B(n_2770),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2790),
.B(n_2781),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2794),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2796),
.B(n_2762),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2795),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2791),
.B(n_2757),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2793),
.B(n_2775),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2789),
.B(n_2777),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2789),
.B(n_2778),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2789),
.B(n_2744),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2789),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2789),
.B(n_2680),
.Y(n_2811)
);

OR2x2_ASAP7_75t_L g2812 ( 
.A(n_2789),
.B(n_2681),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2789),
.Y(n_2813)
);

INVxp67_ASAP7_75t_L g2814 ( 
.A(n_2792),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2789),
.B(n_2685),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2807),
.B(n_2686),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2805),
.B(n_2689),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2809),
.B(n_2815),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2810),
.B(n_2693),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2798),
.Y(n_2820)
);

XNOR2xp5_ASAP7_75t_L g2821 ( 
.A(n_2813),
.B(n_2651),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2812),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2808),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2802),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2803),
.Y(n_2825)
);

AOI32xp33_ASAP7_75t_L g2826 ( 
.A1(n_2806),
.A2(n_2547),
.A3(n_2613),
.B1(n_2725),
.B2(n_2724),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2804),
.B(n_2694),
.Y(n_2827)
);

CKINVDCx5p33_ASAP7_75t_R g2828 ( 
.A(n_2801),
.Y(n_2828)
);

OAI22xp33_ASAP7_75t_SL g2829 ( 
.A1(n_2800),
.A2(n_2721),
.B1(n_2704),
.B2(n_2695),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2799),
.B(n_2696),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2811),
.Y(n_2831)
);

INVxp67_ASAP7_75t_SL g2832 ( 
.A(n_2814),
.Y(n_2832)
);

INVx1_ASAP7_75t_SL g2833 ( 
.A(n_2807),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2807),
.B(n_2705),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2807),
.B(n_2707),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_L g2836 ( 
.A(n_2832),
.B(n_2558),
.C(n_2556),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2828),
.B(n_2709),
.C(n_2708),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2818),
.Y(n_2838)
);

NAND4xp25_ASAP7_75t_L g2839 ( 
.A(n_2833),
.B(n_2599),
.C(n_2719),
.D(n_2714),
.Y(n_2839)
);

AOI211xp5_ASAP7_75t_SL g2840 ( 
.A1(n_2822),
.A2(n_2722),
.B(n_2653),
.C(n_2616),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2816),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2820),
.A2(n_2588),
.B1(n_2592),
.B2(n_2618),
.Y(n_2842)
);

NOR3xp33_ASAP7_75t_L g2843 ( 
.A(n_2825),
.B(n_2639),
.C(n_2617),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2821),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2835),
.B(n_2823),
.Y(n_2845)
);

AOI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2829),
.A2(n_2646),
.B(n_2623),
.Y(n_2846)
);

AOI221xp5_ASAP7_75t_L g2847 ( 
.A1(n_2826),
.A2(n_2578),
.B1(n_2656),
.B2(n_2580),
.C(n_2591),
.Y(n_2847)
);

NOR3x1_ASAP7_75t_L g2848 ( 
.A(n_2817),
.B(n_2834),
.C(n_2819),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2831),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2824),
.B(n_2627),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2827),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_L g2852 ( 
.A(n_2830),
.B(n_2632),
.Y(n_2852)
);

NOR4xp25_ASAP7_75t_L g2853 ( 
.A(n_2833),
.B(n_2624),
.C(n_2660),
.D(n_2615),
.Y(n_2853)
);

INVxp67_ASAP7_75t_L g2854 ( 
.A(n_2818),
.Y(n_2854)
);

NAND4xp25_ASAP7_75t_L g2855 ( 
.A(n_2833),
.B(n_2631),
.C(n_2586),
.D(n_2581),
.Y(n_2855)
);

NOR2x1_ASAP7_75t_L g2856 ( 
.A(n_2818),
.B(n_2598),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2843),
.A2(n_2856),
.B1(n_2849),
.B2(n_2841),
.Y(n_2857)
);

AOI211x1_ASAP7_75t_L g2858 ( 
.A1(n_2846),
.A2(n_2648),
.B(n_2593),
.C(n_2622),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2853),
.B(n_2608),
.Y(n_2859)
);

NAND3xp33_ASAP7_75t_L g2860 ( 
.A(n_2854),
.B(n_2637),
.C(n_2723),
.Y(n_2860)
);

NOR3xp33_ASAP7_75t_SL g2861 ( 
.A(n_2845),
.B(n_260),
.C(n_261),
.Y(n_2861)
);

INVxp67_ASAP7_75t_SL g2862 ( 
.A(n_2848),
.Y(n_2862)
);

AOI211xp5_ASAP7_75t_SL g2863 ( 
.A1(n_2838),
.A2(n_2640),
.B(n_2609),
.C(n_2605),
.Y(n_2863)
);

NOR2x1_ASAP7_75t_L g2864 ( 
.A(n_2837),
.B(n_260),
.Y(n_2864)
);

NOR3xp33_ASAP7_75t_L g2865 ( 
.A(n_2844),
.B(n_2402),
.C(n_2429),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2850),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2840),
.B(n_2630),
.Y(n_2867)
);

NAND4xp25_ASAP7_75t_L g2868 ( 
.A(n_2852),
.B(n_263),
.C(n_261),
.D(n_262),
.Y(n_2868)
);

A2O1A1Ixp33_ASAP7_75t_SL g2869 ( 
.A1(n_2851),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_2869)
);

AOI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2839),
.A2(n_2456),
.B(n_2430),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2855),
.Y(n_2871)
);

NOR3xp33_ASAP7_75t_L g2872 ( 
.A(n_2836),
.B(n_2461),
.C(n_2459),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_SL g2873 ( 
.A(n_2847),
.B(n_264),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2842),
.B(n_265),
.Y(n_2874)
);

NAND4xp25_ASAP7_75t_L g2875 ( 
.A(n_2848),
.B(n_268),
.C(n_265),
.D(n_266),
.Y(n_2875)
);

AOI211xp5_ASAP7_75t_L g2876 ( 
.A1(n_2852),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2855),
.B(n_269),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2856),
.Y(n_2878)
);

NOR3xp33_ASAP7_75t_L g2879 ( 
.A(n_2854),
.B(n_270),
.C(n_271),
.Y(n_2879)
);

AOI311xp33_ASAP7_75t_L g2880 ( 
.A1(n_2838),
.A2(n_274),
.A3(n_272),
.B(n_273),
.C(n_275),
.Y(n_2880)
);

OAI211xp5_ASAP7_75t_L g2881 ( 
.A1(n_2854),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_2881)
);

OAI21xp33_ASAP7_75t_L g2882 ( 
.A1(n_2852),
.A2(n_275),
.B(n_276),
.Y(n_2882)
);

NOR3xp33_ASAP7_75t_SL g2883 ( 
.A(n_2845),
.B(n_276),
.C(n_277),
.Y(n_2883)
);

NOR3xp33_ASAP7_75t_L g2884 ( 
.A(n_2854),
.B(n_278),
.C(n_279),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2853),
.B(n_278),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2856),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2843),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_2887)
);

OA211x2_ASAP7_75t_L g2888 ( 
.A1(n_2854),
.A2(n_283),
.B(n_280),
.C(n_282),
.Y(n_2888)
);

NAND4xp25_ASAP7_75t_L g2889 ( 
.A(n_2848),
.B(n_284),
.C(n_282),
.D(n_283),
.Y(n_2889)
);

NOR3x1_ASAP7_75t_L g2890 ( 
.A(n_2837),
.B(n_285),
.C(n_286),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2856),
.Y(n_2891)
);

NAND4xp25_ASAP7_75t_L g2892 ( 
.A(n_2848),
.B(n_288),
.C(n_286),
.D(n_287),
.Y(n_2892)
);

O2A1O1Ixp33_ASAP7_75t_SL g2893 ( 
.A1(n_2854),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_2893)
);

BUFx2_ASAP7_75t_L g2894 ( 
.A(n_2878),
.Y(n_2894)
);

OAI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2857),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2888),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_2886),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2891),
.Y(n_2898)
);

AOI21xp33_ASAP7_75t_L g2899 ( 
.A1(n_2871),
.A2(n_290),
.B(n_292),
.Y(n_2899)
);

NAND3xp33_ASAP7_75t_L g2900 ( 
.A(n_2861),
.B(n_293),
.C(n_294),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2858),
.B(n_294),
.Y(n_2901)
);

NOR2x1_ASAP7_75t_L g2902 ( 
.A(n_2875),
.B(n_293),
.Y(n_2902)
);

INVxp67_ASAP7_75t_L g2903 ( 
.A(n_2864),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2869),
.B(n_296),
.Y(n_2904)
);

AOI221xp5_ASAP7_75t_L g2905 ( 
.A1(n_2885),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_298),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2859),
.A2(n_300),
.B1(n_295),
.B2(n_299),
.Y(n_2906)
);

AOI211xp5_ASAP7_75t_L g2907 ( 
.A1(n_2862),
.A2(n_300),
.B(n_301),
.C(n_348),
.Y(n_2907)
);

NOR2x1_ASAP7_75t_L g2908 ( 
.A(n_2889),
.B(n_301),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2860),
.B(n_350),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2883),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2893),
.B(n_352),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2890),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2867),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2882),
.A2(n_353),
.B(n_354),
.Y(n_2914)
);

OAI21xp5_ASAP7_75t_SL g2915 ( 
.A1(n_2887),
.A2(n_2892),
.B(n_2877),
.Y(n_2915)
);

AOI221xp5_ASAP7_75t_L g2916 ( 
.A1(n_2874),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.C(n_362),
.Y(n_2916)
);

INVxp67_ASAP7_75t_SL g2917 ( 
.A(n_2876),
.Y(n_2917)
);

AOI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2873),
.A2(n_366),
.B1(n_363),
.B2(n_364),
.Y(n_2918)
);

AO22x2_ASAP7_75t_L g2919 ( 
.A1(n_2866),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2919)
);

AOI221xp5_ASAP7_75t_L g2920 ( 
.A1(n_2872),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.C(n_373),
.Y(n_2920)
);

AOI21xp33_ASAP7_75t_L g2921 ( 
.A1(n_2881),
.A2(n_376),
.B(n_377),
.Y(n_2921)
);

NAND5xp2_ASAP7_75t_SL g2922 ( 
.A(n_2865),
.B(n_381),
.C(n_378),
.D(n_379),
.E(n_382),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2868),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_2923)
);

NOR2x1_ASAP7_75t_L g2924 ( 
.A(n_2880),
.B(n_2870),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2863),
.B(n_388),
.Y(n_2925)
);

BUFx2_ASAP7_75t_L g2926 ( 
.A(n_2879),
.Y(n_2926)
);

OAI211xp5_ASAP7_75t_L g2927 ( 
.A1(n_2884),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2888),
.Y(n_2928)
);

OAI221xp5_ASAP7_75t_L g2929 ( 
.A1(n_2878),
.A2(n_397),
.B1(n_394),
.B2(n_395),
.C(n_399),
.Y(n_2929)
);

OAI21xp5_ASAP7_75t_SL g2930 ( 
.A1(n_2859),
.A2(n_844),
.B(n_841),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2888),
.Y(n_2931)
);

OR2x2_ASAP7_75t_L g2932 ( 
.A(n_2896),
.B(n_402),
.Y(n_2932)
);

NOR3xp33_ASAP7_75t_L g2933 ( 
.A(n_2894),
.B(n_2897),
.C(n_2898),
.Y(n_2933)
);

OR2x2_ASAP7_75t_L g2934 ( 
.A(n_2928),
.B(n_404),
.Y(n_2934)
);

NAND4xp25_ASAP7_75t_L g2935 ( 
.A(n_2931),
.B(n_412),
.C(n_421),
.D(n_401),
.Y(n_2935)
);

NOR2x1_ASAP7_75t_L g2936 ( 
.A(n_2895),
.B(n_405),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2904),
.Y(n_2937)
);

AND2x2_ASAP7_75t_SL g2938 ( 
.A(n_2912),
.B(n_406),
.Y(n_2938)
);

NOR3xp33_ASAP7_75t_L g2939 ( 
.A(n_2913),
.B(n_407),
.C(n_408),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2924),
.B(n_409),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2910),
.B(n_410),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2925),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2902),
.B(n_411),
.Y(n_2943)
);

NAND4xp75_ASAP7_75t_L g2944 ( 
.A(n_2899),
.B(n_416),
.C(n_413),
.D(n_415),
.Y(n_2944)
);

NOR2xp67_ASAP7_75t_L g2945 ( 
.A(n_2906),
.B(n_417),
.Y(n_2945)
);

NOR2xp67_ASAP7_75t_SL g2946 ( 
.A(n_2911),
.B(n_2929),
.Y(n_2946)
);

NOR2xp67_ASAP7_75t_L g2947 ( 
.A(n_2901),
.B(n_418),
.Y(n_2947)
);

OAI211xp5_ASAP7_75t_L g2948 ( 
.A1(n_2930),
.A2(n_422),
.B(n_419),
.C(n_420),
.Y(n_2948)
);

NOR4xp25_ASAP7_75t_L g2949 ( 
.A(n_2903),
.B(n_427),
.C(n_424),
.D(n_425),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2908),
.Y(n_2950)
);

NAND4xp75_ASAP7_75t_L g2951 ( 
.A(n_2909),
.B(n_431),
.C(n_428),
.D(n_429),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2900),
.Y(n_2952)
);

HB1xp67_ASAP7_75t_L g2953 ( 
.A(n_2922),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2917),
.Y(n_2954)
);

AOI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2915),
.A2(n_437),
.B1(n_432),
.B2(n_436),
.Y(n_2955)
);

INVx3_ASAP7_75t_SL g2956 ( 
.A(n_2919),
.Y(n_2956)
);

NOR2xp67_ASAP7_75t_L g2957 ( 
.A(n_2927),
.B(n_438),
.Y(n_2957)
);

NAND4xp75_ASAP7_75t_L g2958 ( 
.A(n_2905),
.B(n_444),
.C(n_440),
.D(n_442),
.Y(n_2958)
);

NOR2x1_ASAP7_75t_L g2959 ( 
.A(n_2926),
.B(n_445),
.Y(n_2959)
);

OAI21xp33_ASAP7_75t_SL g2960 ( 
.A1(n_2921),
.A2(n_446),
.B(n_447),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2907),
.B(n_448),
.Y(n_2961)
);

NOR3xp33_ASAP7_75t_L g2962 ( 
.A(n_2916),
.B(n_2920),
.C(n_2918),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2923),
.B(n_450),
.Y(n_2963)
);

NOR3x1_ASAP7_75t_L g2964 ( 
.A(n_2914),
.B(n_454),
.C(n_453),
.Y(n_2964)
);

INVxp67_ASAP7_75t_L g2965 ( 
.A(n_2919),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2894),
.Y(n_2966)
);

NOR3xp33_ASAP7_75t_L g2967 ( 
.A(n_2894),
.B(n_451),
.C(n_456),
.Y(n_2967)
);

OAI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2894),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.Y(n_2968)
);

AND2x4_ASAP7_75t_L g2969 ( 
.A(n_2897),
.B(n_460),
.Y(n_2969)
);

NAND3xp33_ASAP7_75t_L g2970 ( 
.A(n_2894),
.B(n_461),
.C(n_462),
.Y(n_2970)
);

OAI21xp33_ASAP7_75t_L g2971 ( 
.A1(n_2896),
.A2(n_463),
.B(n_464),
.Y(n_2971)
);

NOR3xp33_ASAP7_75t_L g2972 ( 
.A(n_2894),
.B(n_466),
.C(n_467),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2894),
.Y(n_2973)
);

NOR2x1_ASAP7_75t_L g2974 ( 
.A(n_2894),
.B(n_468),
.Y(n_2974)
);

NAND4xp75_ASAP7_75t_L g2975 ( 
.A(n_2924),
.B(n_473),
.C(n_469),
.D(n_470),
.Y(n_2975)
);

HB1xp67_ASAP7_75t_L g2976 ( 
.A(n_2896),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2966),
.Y(n_2977)
);

OR2x2_ASAP7_75t_L g2978 ( 
.A(n_2973),
.B(n_474),
.Y(n_2978)
);

NOR2xp67_ASAP7_75t_L g2979 ( 
.A(n_2976),
.B(n_475),
.Y(n_2979)
);

OAI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2933),
.A2(n_476),
.B(n_479),
.Y(n_2980)
);

NOR2xp67_ASAP7_75t_L g2981 ( 
.A(n_2954),
.B(n_481),
.Y(n_2981)
);

NAND4xp75_ASAP7_75t_L g2982 ( 
.A(n_2940),
.B(n_485),
.C(n_482),
.D(n_483),
.Y(n_2982)
);

NOR3xp33_ASAP7_75t_L g2983 ( 
.A(n_2937),
.B(n_486),
.C(n_488),
.Y(n_2983)
);

AOI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2953),
.A2(n_489),
.B(n_490),
.Y(n_2984)
);

O2A1O1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2950),
.A2(n_495),
.B(n_491),
.C(n_494),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2943),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2956),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_L g2988 ( 
.A(n_2965),
.B(n_496),
.Y(n_2988)
);

BUFx2_ASAP7_75t_L g2989 ( 
.A(n_2969),
.Y(n_2989)
);

NAND3xp33_ASAP7_75t_SL g2990 ( 
.A(n_2942),
.B(n_499),
.C(n_498),
.Y(n_2990)
);

OAI22xp5_ASAP7_75t_L g2991 ( 
.A1(n_2952),
.A2(n_501),
.B1(n_497),
.B2(n_500),
.Y(n_2991)
);

AOI21xp33_ASAP7_75t_L g2992 ( 
.A1(n_2974),
.A2(n_503),
.B(n_505),
.Y(n_2992)
);

OAI221xp5_ASAP7_75t_L g2993 ( 
.A1(n_2957),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.C(n_509),
.Y(n_2993)
);

NOR3xp33_ASAP7_75t_L g2994 ( 
.A(n_2941),
.B(n_510),
.C(n_511),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2961),
.B(n_513),
.Y(n_2995)
);

INVxp33_ASAP7_75t_L g2996 ( 
.A(n_2959),
.Y(n_2996)
);

INVx3_ASAP7_75t_L g2997 ( 
.A(n_2969),
.Y(n_2997)
);

INVxp67_ASAP7_75t_L g2998 ( 
.A(n_2938),
.Y(n_2998)
);

NOR2xp33_ASAP7_75t_L g2999 ( 
.A(n_2960),
.B(n_514),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2932),
.Y(n_3000)
);

NAND4xp25_ASAP7_75t_SL g3001 ( 
.A(n_2936),
.B(n_519),
.C(n_517),
.D(n_518),
.Y(n_3001)
);

OAI211xp5_ASAP7_75t_L g3002 ( 
.A1(n_2971),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2934),
.Y(n_3003)
);

INVxp67_ASAP7_75t_SL g3004 ( 
.A(n_2947),
.Y(n_3004)
);

AO22x2_ASAP7_75t_L g3005 ( 
.A1(n_2975),
.A2(n_2944),
.B1(n_2958),
.B2(n_2970),
.Y(n_3005)
);

INVxp67_ASAP7_75t_L g3006 ( 
.A(n_2946),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2964),
.Y(n_3007)
);

OR5x1_ASAP7_75t_L g3008 ( 
.A(n_2948),
.B(n_527),
.C(n_523),
.D(n_525),
.E(n_528),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2963),
.B(n_529),
.Y(n_3009)
);

OAI21xp33_ASAP7_75t_L g3010 ( 
.A1(n_2962),
.A2(n_530),
.B(n_531),
.Y(n_3010)
);

NOR2x1_ASAP7_75t_L g3011 ( 
.A(n_2935),
.B(n_532),
.Y(n_3011)
);

AOI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2945),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_3012)
);

NOR4xp75_ASAP7_75t_SL g3013 ( 
.A(n_2968),
.B(n_538),
.C(n_536),
.D(n_537),
.Y(n_3013)
);

INVx4_ASAP7_75t_L g3014 ( 
.A(n_2987),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_3007),
.A2(n_2967),
.B1(n_2972),
.B2(n_2939),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2977),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2989),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2997),
.Y(n_3018)
);

OAI22xp5_ASAP7_75t_SL g3019 ( 
.A1(n_3006),
.A2(n_2949),
.B1(n_2955),
.B2(n_2951),
.Y(n_3019)
);

OAI211xp5_ASAP7_75t_L g3020 ( 
.A1(n_2980),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_3020)
);

INVxp67_ASAP7_75t_L g3021 ( 
.A(n_2997),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_3004),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2981),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2999),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2979),
.B(n_545),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2978),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2998),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_3000),
.Y(n_3028)
);

INVx5_ASAP7_75t_L g3029 ( 
.A(n_2995),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_3003),
.Y(n_3030)
);

INVxp33_ASAP7_75t_L g3031 ( 
.A(n_3009),
.Y(n_3031)
);

AOI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2986),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_3032)
);

AND2x4_ASAP7_75t_L g3033 ( 
.A(n_3011),
.B(n_2988),
.Y(n_3033)
);

OAI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2996),
.A2(n_2993),
.B1(n_3005),
.B2(n_3012),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_3005),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_3013),
.B(n_549),
.Y(n_3036)
);

XOR2x1_ASAP7_75t_L g3037 ( 
.A(n_2991),
.B(n_551),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_3008),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2994),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2984),
.B(n_3010),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2982),
.Y(n_3041)
);

NOR3xp33_ASAP7_75t_L g3042 ( 
.A(n_2992),
.B(n_555),
.C(n_556),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_3001),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_3029),
.B(n_2983),
.Y(n_3044)
);

AND2x4_ASAP7_75t_L g3045 ( 
.A(n_3016),
.B(n_2990),
.Y(n_3045)
);

OR2x2_ASAP7_75t_L g3046 ( 
.A(n_3014),
.B(n_3002),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_SL g3047 ( 
.A1(n_3022),
.A2(n_2985),
.B(n_557),
.Y(n_3047)
);

HB1xp67_ASAP7_75t_L g3048 ( 
.A(n_3029),
.Y(n_3048)
);

NAND2x1_ASAP7_75t_L g3049 ( 
.A(n_3035),
.B(n_558),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_3021),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.Y(n_3050)
);

AOI22xp5_ASAP7_75t_L g3051 ( 
.A1(n_3027),
.A2(n_3017),
.B1(n_3018),
.B2(n_3028),
.Y(n_3051)
);

AO22x2_ASAP7_75t_L g3052 ( 
.A1(n_3030),
.A2(n_565),
.B1(n_562),
.B2(n_564),
.Y(n_3052)
);

AND3x4_ASAP7_75t_L g3053 ( 
.A(n_3038),
.B(n_567),
.C(n_568),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_3033),
.A2(n_3019),
.B1(n_3034),
.B2(n_3031),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3037),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_3036),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_3026),
.Y(n_3057)
);

OAI22xp33_ASAP7_75t_SL g3058 ( 
.A1(n_3023),
.A2(n_3025),
.B1(n_3040),
.B2(n_3043),
.Y(n_3058)
);

OAI22xp5_ASAP7_75t_L g3059 ( 
.A1(n_3015),
.A2(n_3024),
.B1(n_3041),
.B2(n_3039),
.Y(n_3059)
);

AOI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_3042),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3060)
);

NAND5xp2_ASAP7_75t_L g3061 ( 
.A(n_3020),
.B(n_575),
.C(n_572),
.D(n_573),
.E(n_576),
.Y(n_3061)
);

XNOR2xp5_ASAP7_75t_L g3062 ( 
.A(n_3032),
.B(n_577),
.Y(n_3062)
);

AOI21xp33_ASAP7_75t_L g3063 ( 
.A1(n_3016),
.A2(n_578),
.B(n_579),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_3016),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_3029),
.B(n_580),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_3053),
.Y(n_3066)
);

AND2x4_ASAP7_75t_L g3067 ( 
.A(n_3056),
.B(n_581),
.Y(n_3067)
);

OR3x1_ASAP7_75t_L g3068 ( 
.A(n_3064),
.B(n_584),
.C(n_585),
.Y(n_3068)
);

AOI221xp5_ASAP7_75t_L g3069 ( 
.A1(n_3048),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.C(n_591),
.Y(n_3069)
);

OA22x2_ASAP7_75t_L g3070 ( 
.A1(n_3054),
.A2(n_596),
.B1(n_593),
.B2(n_595),
.Y(n_3070)
);

OA22x2_ASAP7_75t_L g3071 ( 
.A1(n_3051),
.A2(n_601),
.B1(n_597),
.B2(n_600),
.Y(n_3071)
);

AOI22x1_ASAP7_75t_L g3072 ( 
.A1(n_3046),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_3072)
);

OAI221xp5_ASAP7_75t_L g3073 ( 
.A1(n_3057),
.A2(n_612),
.B1(n_606),
.B2(n_609),
.C(n_614),
.Y(n_3073)
);

OA22x2_ASAP7_75t_L g3074 ( 
.A1(n_3045),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_3074)
);

AOI221xp5_ASAP7_75t_L g3075 ( 
.A1(n_3058),
.A2(n_621),
.B1(n_618),
.B2(n_619),
.C(n_622),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_SL g3076 ( 
.A1(n_3055),
.A2(n_627),
.B1(n_623),
.B2(n_624),
.Y(n_3076)
);

XNOR2xp5_ASAP7_75t_L g3077 ( 
.A(n_3068),
.B(n_3049),
.Y(n_3077)
);

OR5x1_ASAP7_75t_L g3078 ( 
.A(n_3066),
.B(n_3047),
.C(n_3059),
.D(n_3044),
.E(n_3062),
.Y(n_3078)
);

NOR3xp33_ASAP7_75t_L g3079 ( 
.A(n_3075),
.B(n_3065),
.C(n_3063),
.Y(n_3079)
);

NOR3xp33_ASAP7_75t_L g3080 ( 
.A(n_3076),
.B(n_3061),
.C(n_3050),
.Y(n_3080)
);

NAND3xp33_ASAP7_75t_SL g3081 ( 
.A(n_3069),
.B(n_3060),
.C(n_3052),
.Y(n_3081)
);

AOI211xp5_ASAP7_75t_L g3082 ( 
.A1(n_3073),
.A2(n_3052),
.B(n_631),
.C(n_629),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3067),
.B(n_630),
.Y(n_3083)
);

NOR3xp33_ASAP7_75t_L g3084 ( 
.A(n_3070),
.B(n_632),
.C(n_633),
.Y(n_3084)
);

AOI211xp5_ASAP7_75t_L g3085 ( 
.A1(n_3074),
.A2(n_639),
.B(n_635),
.C(n_637),
.Y(n_3085)
);

OAI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_3077),
.A2(n_3071),
.B(n_3072),
.Y(n_3086)
);

AOI22xp33_ASAP7_75t_L g3087 ( 
.A1(n_3080),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_3087)
);

OAI22x1_ASAP7_75t_L g3088 ( 
.A1(n_3083),
.A2(n_645),
.B1(n_643),
.B2(n_644),
.Y(n_3088)
);

AOI21x1_ASAP7_75t_L g3089 ( 
.A1(n_3078),
.A2(n_646),
.B(n_647),
.Y(n_3089)
);

AOI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_3079),
.A2(n_652),
.B1(n_649),
.B2(n_651),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_3082),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_3084),
.B(n_659),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3089),
.Y(n_3093)
);

XNOR2xp5_ASAP7_75t_L g3094 ( 
.A(n_3086),
.B(n_3081),
.Y(n_3094)
);

XNOR2xp5_ASAP7_75t_L g3095 ( 
.A(n_3091),
.B(n_3085),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3092),
.B(n_660),
.Y(n_3096)
);

AOI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_3087),
.A2(n_851),
.B1(n_663),
.B2(n_661),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_3090),
.A2(n_665),
.B1(n_662),
.B2(n_664),
.Y(n_3098)
);

NOR3xp33_ASAP7_75t_L g3099 ( 
.A(n_3088),
.B(n_666),
.C(n_668),
.Y(n_3099)
);

CKINVDCx20_ASAP7_75t_R g3100 ( 
.A(n_3094),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3093),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3096),
.Y(n_3102)
);

AOI22xp5_ASAP7_75t_SL g3103 ( 
.A1(n_3095),
.A2(n_850),
.B1(n_673),
.B2(n_670),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3099),
.Y(n_3104)
);

AOI22xp33_ASAP7_75t_SL g3105 ( 
.A1(n_3100),
.A2(n_3098),
.B1(n_3097),
.B2(n_679),
.Y(n_3105)
);

AO21x2_ASAP7_75t_L g3106 ( 
.A1(n_3101),
.A2(n_672),
.B(n_676),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_3102),
.A2(n_682),
.B(n_683),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_3106),
.A2(n_3104),
.B1(n_3103),
.B2(n_687),
.Y(n_3108)
);

NOR2xp33_ASAP7_75t_L g3109 ( 
.A(n_3105),
.B(n_684),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_3109),
.Y(n_3110)
);

OR2x6_ASAP7_75t_L g3111 ( 
.A(n_3110),
.B(n_3107),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_3111),
.A2(n_3108),
.B1(n_690),
.B2(n_685),
.Y(n_3112)
);

AOI211xp5_ASAP7_75t_L g3113 ( 
.A1(n_3112),
.A2(n_692),
.B(n_689),
.C(n_691),
.Y(n_3113)
);


endmodule