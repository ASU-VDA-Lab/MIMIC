module fake_jpeg_19548_n_189 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_30),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_23),
.B1(n_20),
.B2(n_29),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_59),
.B1(n_77),
.B2(n_22),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_41),
.B1(n_35),
.B2(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_60),
.B1(n_72),
.B2(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_20),
.B1(n_29),
.B2(n_36),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_41),
.B1(n_46),
.B2(n_54),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_38),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_32),
.B(n_37),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_38),
.B1(n_29),
.B2(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_21),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_26),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_82),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_99),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_21),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_95),
.C(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_97),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_67),
.B(n_75),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_15),
.C(n_16),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_17),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_17),
.B1(n_26),
.B2(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_86),
.A3(n_99),
.B1(n_87),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_119),
.B(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_120),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_95),
.Y(n_128)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_113),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_1),
.B(n_2),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_72),
.B1(n_69),
.B2(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_122),
.B1(n_82),
.B2(n_90),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_15),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_79),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_63),
.B1(n_67),
.B2(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_135),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_84),
.C(n_118),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.C(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_126),
.B1(n_132),
.B2(n_138),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_84),
.B1(n_91),
.B2(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_133),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_80),
.C(n_82),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_92),
.B1(n_64),
.B2(n_71),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_92),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_74),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_106),
.B(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_64),
.B1(n_73),
.B2(n_15),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_128),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_114),
.A3(n_129),
.B1(n_110),
.B2(n_130),
.C(n_137),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_132),
.B1(n_133),
.B2(n_125),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_115),
.B(n_122),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_131),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_145),
.C(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_157),
.C(n_102),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_151),
.B(n_111),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_134),
.C(n_130),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_147),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_140),
.C(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_162),
.B1(n_140),
.B2(n_136),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_108),
.B1(n_107),
.B2(n_119),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_166),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_165),
.B1(n_170),
.B2(n_153),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_136),
.B1(n_113),
.B2(n_102),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_15),
.C(n_73),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_136),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_15),
.C(n_21),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_2),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_177),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.C(n_184),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_3),
.B1(n_7),
.B2(n_9),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_183),
.B(n_11),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_13),
.B(n_9),
.C(n_12),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_12),
.B(n_13),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);


endmodule