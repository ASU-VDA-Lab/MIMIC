module real_jpeg_33320_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_633, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_633;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_620;
wire n_332;
wire n_456;
wire n_578;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_0),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_0),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_0),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_1),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_1),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_1),
.A2(n_149),
.B1(n_209),
.B2(n_214),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_1),
.A2(n_149),
.B1(n_366),
.B2(n_370),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g620 ( 
.A1(n_1),
.A2(n_149),
.B1(n_621),
.B2(n_623),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_3),
.A2(n_100),
.B1(n_265),
.B2(n_269),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_3),
.A2(n_100),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_3),
.A2(n_100),
.B1(n_238),
.B2(n_479),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_134),
.B1(n_139),
.B2(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_4),
.A2(n_139),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_4),
.A2(n_139),
.B1(n_423),
.B2(n_425),
.Y(n_422)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_5),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_6),
.B(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_6),
.A2(n_189),
.B(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_R g300 ( 
.A(n_6),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_6),
.A2(n_300),
.B1(n_495),
.B2(n_497),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_6),
.B(n_83),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_6),
.A2(n_159),
.B1(n_567),
.B2(n_571),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_7),
.A2(n_326),
.B1(n_327),
.B2(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_7),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_7),
.A2(n_326),
.B1(n_414),
.B2(n_418),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_11),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_11),
.Y(n_242)
);

AOI22x1_ASAP7_75t_L g391 ( 
.A1(n_11),
.A2(n_242),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_11),
.A2(n_242),
.B1(n_342),
.B2(n_613),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_106),
.B1(n_112),
.B2(n_116),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_12),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_12),
.A2(n_116),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_12),
.A2(n_116),
.B1(n_458),
.B2(n_463),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_12),
.A2(n_116),
.B1(n_508),
.B2(n_510),
.Y(n_507)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_13),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_14),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_14),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_14),
.A2(n_232),
.B1(n_293),
.B2(n_297),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_14),
.A2(n_232),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_14),
.A2(n_48),
.B1(n_232),
.B2(n_433),
.Y(n_432)
);

AOI22x1_ASAP7_75t_SL g46 ( 
.A1(n_15),
.A2(n_47),
.B1(n_54),
.B2(n_60),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_15),
.A2(n_60),
.B1(n_251),
.B2(n_256),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_15),
.A2(n_60),
.B1(n_214),
.B2(n_489),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_15),
.A2(n_60),
.B1(n_559),
.B2(n_561),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_21),
.B(n_630),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_16),
.B(n_631),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_17),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_17),
.A2(n_66),
.B1(n_282),
.B2(n_288),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_17),
.A2(n_66),
.B1(n_229),
.B2(n_516),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_17),
.A2(n_66),
.B1(n_568),
.B2(n_570),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_18),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_18),
.Y(n_491)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_19),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_R g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_595),
.B2(n_629),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_447),
.B(n_590),
.Y(n_24)
);

NAND4xp25_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_303),
.C(n_401),
.D(n_439),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_273),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_27),
.B(n_273),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_192),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_28),
.A2(n_441),
.B(n_442),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_129),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_81),
.Y(n_29)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_30),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_44),
.B(n_61),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22x1_ASAP7_75t_L g431 ( 
.A1(n_32),
.A2(n_70),
.B1(n_376),
.B2(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_32),
.A2(n_432),
.B1(n_619),
.B2(n_620),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_33),
.A2(n_63),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

NOR2x1_ASAP7_75t_R g299 ( 
.A(n_33),
.B(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_33),
.A2(n_46),
.B1(n_260),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_33),
.A2(n_260),
.B1(n_348),
.B2(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_35)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_36),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_39),
.Y(n_183)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_41),
.Y(n_616)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_53),
.Y(n_174)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_53),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_53),
.Y(n_435)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_57),
.Y(n_191)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_58),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_59),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_72),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_77),
.Y(n_378)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_77),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_77),
.Y(n_624)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_81),
.B(n_129),
.C(n_306),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_96),
.B1(n_105),
.B2(n_117),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_82),
.A2(n_105),
.B1(n_117),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_82),
.A2(n_250),
.B(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_82),
.A2(n_96),
.B1(n_117),
.B2(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_82),
.A2(n_117),
.B1(n_281),
.B2(n_494),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_82),
.A2(n_117),
.B1(n_611),
.B2(n_612),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22x1_ASAP7_75t_SL g363 ( 
.A1(n_83),
.A2(n_279),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_83),
.A2(n_279),
.B1(n_365),
.B2(n_422),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AO21x2_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_118),
.B(n_123),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_89),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_89),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_90),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_90),
.Y(n_317)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_90),
.Y(n_417)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_94),
.B(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_94),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_95),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_95),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_99),
.Y(n_426)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_104),
.Y(n_258)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_114),
.Y(n_424)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_115),
.Y(n_498)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_117),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_123),
.A2(n_468),
.B(n_473),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_125),
.Y(n_288)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_165),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_130),
.A2(n_131),
.B1(n_165),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_142),
.B1(n_148),
.B2(n_158),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_133),
.A2(n_159),
.B1(n_236),
.B2(n_245),
.Y(n_235)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_138),
.Y(n_509)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

BUFx2_ASAP7_75t_SL g298 ( 
.A(n_141),
.Y(n_298)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_143),
.B(n_300),
.Y(n_573)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_147),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_147),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_148),
.A2(n_158),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_154),
.Y(n_540)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g477 ( 
.A1(n_158),
.A2(n_292),
.B1(n_478),
.B2(n_482),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_158),
.A2(n_320),
.B1(n_556),
.B2(n_557),
.Y(n_555)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_159),
.A2(n_236),
.B(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_159),
.A2(n_325),
.B(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_159),
.A2(n_503),
.B1(n_506),
.B2(n_507),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_159),
.A2(n_503),
.B1(n_558),
.B2(n_567),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_162),
.Y(n_562)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_163),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_164),
.Y(n_482)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_164),
.Y(n_571)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_165),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_175),
.B1(n_178),
.B2(n_188),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_187),
.Y(n_372)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_248),
.B1(n_271),
.B2(n_272),
.Y(n_192)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_235),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_194),
.B(n_235),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_208),
.B1(n_217),
.B2(n_228),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_195),
.A2(n_208),
.B1(n_217),
.B2(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_195),
.A2(n_217),
.B1(n_488),
.B2(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AO21x2_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_218),
.B(n_224),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_201),
.Y(n_542)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_217),
.A2(n_228),
.B1(n_264),
.B2(n_270),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_217),
.A2(n_270),
.B1(n_310),
.B2(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_217),
.Y(n_411)
);

AOI21xp33_ASAP7_75t_SL g608 ( 
.A1(n_217),
.A2(n_270),
.B(n_413),
.Y(n_608)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_217),
.A2(n_270),
.B(n_413),
.Y(n_617)
);

NAND2xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_222),
.Y(n_464)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_222),
.Y(n_533)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_223),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_223),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_224),
.Y(n_546)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_231),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_241),
.Y(n_332)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_241),
.Y(n_481)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_241),
.Y(n_576)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_243),
.Y(n_510)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_245),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.C(n_263),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_263),
.Y(n_275)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_255),
.Y(n_496)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_260),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_264),
.A2(n_270),
.B1(n_456),
.B2(n_465),
.Y(n_455)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_270),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_270),
.B(n_300),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_271),
.B(n_272),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_R g442 ( 
.A(n_271),
.B(n_272),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.C(n_301),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_274),
.B(n_587),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_276),
.B(n_301),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_289),
.C(n_299),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_277),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_284),
.Y(n_476)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_289),
.A2(n_290),
.B1(n_299),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_299),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_300),
.B(n_469),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_300),
.B(n_474),
.C(n_476),
.Y(n_473)
);

OAI21xp33_ASAP7_75t_SL g527 ( 
.A1(n_300),
.A2(n_528),
.B(n_530),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_300),
.B(n_531),
.Y(n_530)
);

A2O1A1O1Ixp25_ASAP7_75t_L g590 ( 
.A1(n_303),
.A2(n_401),
.B(n_591),
.C(n_593),
.D(n_594),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_357),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_304),
.B(n_357),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_333),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_305),
.B(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_308),
.A2(n_334),
.B1(n_335),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_308),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_318),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_309),
.B(n_318),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_328),
.Y(n_545)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_332),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_356),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_338),
.C(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_336),
.B(n_445),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_346),
.B(n_355),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_346),
.Y(n_355)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_383),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_384),
.C(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_381),
.B2(n_382),
.Y(n_359)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_373),
.B2(n_374),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_382),
.C(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_399),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_389),
.B(n_398),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_390),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_385),
.A2(n_386),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_386),
.B(n_390),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_386),
.Y(n_605)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_391),
.Y(n_410)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx2_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_399),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_402),
.B(n_404),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_405),
.B(n_438),
.C(n_626),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_428),
.B1(n_437),
.B2(n_438),
.Y(n_407)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_421),
.B(n_427),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_421),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_420),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

AOI22x1_ASAP7_75t_L g486 ( 
.A1(n_411),
.A2(n_420),
.B1(n_457),
.B2(n_487),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_411),
.A2(n_420),
.B1(n_515),
.B2(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_422),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx8_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_427),
.Y(n_601)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_428),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_436),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_431),
.Y(n_604)
);

INVx8_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_436),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_440),
.B(n_443),
.C(n_592),
.Y(n_591)
);

AOI21x1_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_585),
.B(n_589),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_499),
.B(n_584),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_483),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_450),
.B(n_483),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_451),
.B(n_455),
.C(n_466),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_466),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_477),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_467),
.B(n_477),
.Y(n_484)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_472),
.Y(n_475)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_478),
.Y(n_506)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_481),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.C(n_492),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_484),
.B(n_519),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_486),
.A2(n_492),
.B(n_520),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

AOI31xp67_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_522),
.A3(n_550),
.B(n_583),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_518),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_501),
.B(n_518),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_511),
.C(n_512),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_507),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_509),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_511),
.B(n_513),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_549),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_547),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_547),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_525),
.B(n_534),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_525),
.B(n_535),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_525),
.A2(n_535),
.B(n_554),
.Y(n_582)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_526),
.B(n_534),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_529),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_543),
.B1(n_544),
.B2(n_546),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_537),
.B(n_541),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_551),
.C(n_563),
.Y(n_550)
);

AO21x1_ASAP7_75t_L g551 ( 
.A1(n_552),
.A2(n_553),
.B(n_555),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_582),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_581),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_577),
.B(n_580),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_566),
.B(n_572),
.Y(n_565)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_573),
.B(n_574),
.Y(n_572)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

BUFx12f_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_579),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_578),
.B(n_579),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_586),
.B(n_588),
.Y(n_585)
);

NOR2x1_ASAP7_75t_L g589 ( 
.A(n_586),
.B(n_588),
.Y(n_589)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_595),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_627),
.Y(n_595)
);

INVxp33_ASAP7_75t_SL g596 ( 
.A(n_597),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_625),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_625),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_606),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_601),
.B(n_602),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_603),
.A2(n_604),
.B1(n_605),
.B2(n_633),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_618),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_608),
.A2(n_609),
.B1(n_610),
.B2(n_617),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_610),
.Y(n_609)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);


endmodule