module real_aes_7287_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_1170;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1175;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_905;
wire n_518;
wire n_792;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_1034;
wire n_923;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1160;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_1078;
wire n_495;
wire n_892;
wire n_994;
wire n_1072;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_1053;
wire n_872;
wire n_906;
wire n_477;
wire n_1182;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1189;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_1168;
wire n_755;
wire n_1025;
wire n_1148;
wire n_409;
wire n_781;
wire n_860;
wire n_909;
wire n_523;
wire n_748;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1081;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_1198;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_812;
wire n_534;
wire n_925;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1196;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_1174;
wire n_1100;
wire n_1167;
wire n_1193;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_1179;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1157;
wire n_1158;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_1187;
wire n_727;
wire n_1083;
wire n_749;
wire n_663;
wire n_1056;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_1162;
wire n_861;
wire n_705;
wire n_1191;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_1190;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_719;
wire n_566;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1156;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_1185;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1101;
wire n_447;
wire n_1102;
wire n_1173;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_1119;
wire n_802;
wire n_868;
wire n_877;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_0), .A2(n_185), .B1(n_934), .B2(n_935), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_1), .B(n_471), .Y(n_508) );
XOR2x2_ASAP7_75t_L g414 ( .A(n_2), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_3), .A2(n_316), .B1(n_606), .B2(n_871), .Y(n_870) );
OA22x2_ASAP7_75t_L g883 ( .A1(n_4), .A2(n_884), .B1(n_885), .B2(n_910), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_4), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_5), .A2(n_176), .B1(n_470), .B2(n_663), .C(n_664), .Y(n_662) );
OA22x2_ASAP7_75t_L g852 ( .A1(n_6), .A2(n_853), .B1(n_854), .B2(n_878), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_6), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g1144 ( .A(n_7), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_8), .A2(n_97), .B1(n_749), .B2(n_874), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_9), .A2(n_301), .B1(n_545), .B2(n_639), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_10), .A2(n_365), .B1(n_625), .B2(n_626), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_11), .Y(n_695) );
AO22x2_ASAP7_75t_L g433 ( .A1(n_12), .A2(n_231), .B1(n_424), .B2(n_429), .Y(n_433) );
INVx1_ASAP7_75t_L g1130 ( .A(n_12), .Y(n_1130) );
AOI22xp5_ASAP7_75t_SL g1066 ( .A1(n_13), .A2(n_395), .B1(n_705), .B2(n_935), .Y(n_1066) );
AOI222xp33_ASAP7_75t_L g996 ( .A1(n_14), .A2(n_63), .B1(n_339), .B2(n_642), .C1(n_669), .C2(n_997), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_15), .A2(n_317), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_16), .A2(n_70), .B1(n_591), .B2(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_SL g1061 ( .A1(n_17), .A2(n_257), .B1(n_701), .B2(n_1062), .Y(n_1061) );
AO22x1_ASAP7_75t_L g943 ( .A1(n_18), .A2(n_944), .B1(n_967), .B2(n_968), .Y(n_943) );
INVx1_ASAP7_75t_L g967 ( .A(n_18), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_19), .A2(n_113), .B1(n_629), .B2(n_699), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_20), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_21), .A2(n_25), .B1(n_637), .B2(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_22), .A2(n_390), .B1(n_894), .B2(n_961), .Y(n_960) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_23), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_24), .A2(n_386), .B1(n_451), .B2(n_453), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_26), .A2(n_277), .B1(n_514), .B2(n_516), .Y(n_816) );
INVx1_ASAP7_75t_L g484 ( .A(n_27), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_28), .A2(n_259), .B1(n_470), .B2(n_990), .C(n_991), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_29), .A2(n_378), .B1(n_451), .B2(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_30), .A2(n_186), .B1(n_473), .B2(n_1059), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_31), .A2(n_355), .B1(n_524), .B2(n_525), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_32), .A2(n_106), .B1(n_486), .B2(n_490), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_33), .A2(n_974), .B1(n_998), .B2(n_999), .Y(n_973) );
INVx1_ASAP7_75t_L g998 ( .A(n_33), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_34), .A2(n_59), .B1(n_622), .B2(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_35), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_36), .A2(n_266), .B1(n_477), .B2(n_637), .Y(n_1174) );
AO22x2_ASAP7_75t_L g431 ( .A1(n_37), .A2(n_119), .B1(n_424), .B2(n_425), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_38), .A2(n_272), .B1(n_560), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_39), .A2(n_206), .B1(n_562), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_40), .A2(n_331), .B1(n_514), .B2(n_1189), .Y(n_1188) );
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_41), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_42), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_43), .A2(n_267), .B1(n_633), .B2(n_790), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g1085 ( .A(n_44), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_45), .A2(n_348), .B1(n_504), .B2(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_46), .A2(n_343), .B1(n_565), .B2(n_753), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_47), .A2(n_237), .B1(n_620), .B2(n_732), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_48), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_49), .B(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_50), .A2(n_288), .B1(n_420), .B2(n_605), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_51), .A2(n_241), .B1(n_620), .B2(n_626), .Y(n_966) );
AOI222xp33_ASAP7_75t_L g1159 ( .A1(n_52), .A2(n_158), .B1(n_311), .B2(n_642), .C1(n_902), .C2(n_1160), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_53), .A2(n_281), .B1(n_543), .B2(n_544), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_54), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_55), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_56), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_57), .A2(n_203), .B1(n_544), .B2(n_671), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_58), .A2(n_154), .B1(n_444), .B2(n_701), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_60), .B(n_482), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_61), .A2(n_220), .B1(n_333), .B2(n_590), .C1(n_669), .C2(n_671), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_62), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_64), .A2(n_380), .B1(n_567), .B2(n_622), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_65), .A2(n_223), .B1(n_462), .B2(n_876), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_66), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_67), .A2(n_197), .B1(n_841), .B2(n_894), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_68), .Y(n_1099) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_69), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_71), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_72), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_73), .A2(n_379), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_74), .A2(n_313), .B1(n_513), .B2(n_514), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_75), .A2(n_342), .B1(n_625), .B2(n_965), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_76), .A2(n_213), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_77), .A2(n_115), .B1(n_604), .B2(n_661), .Y(n_962) );
INVx1_ASAP7_75t_L g1068 ( .A(n_78), .Y(n_1068) );
AOI222xp33_ASAP7_75t_L g1040 ( .A1(n_79), .A2(n_211), .B1(n_251), .B2(n_723), .C1(n_724), .C2(n_769), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1081 ( .A(n_80), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g1102 ( .A1(n_81), .A2(n_214), .B1(n_477), .B2(n_637), .Y(n_1102) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_82), .A2(n_86), .B1(n_843), .B2(n_845), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_83), .A2(n_294), .B1(n_609), .B2(n_798), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_84), .A2(n_111), .B1(n_630), .B2(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_85), .A2(n_283), .B1(n_453), .B2(n_630), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_87), .A2(n_157), .B1(n_418), .B2(n_513), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_88), .A2(n_268), .B1(n_474), .B2(n_487), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_89), .A2(n_245), .B1(n_699), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_90), .A2(n_253), .B1(n_707), .B2(n_841), .Y(n_840) );
AOI22xp5_ASAP7_75t_SL g1063 ( .A1(n_91), .A2(n_264), .B1(n_444), .B2(n_1064), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_92), .A2(n_238), .B1(n_486), .B2(n_763), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_93), .Y(n_581) );
OA22x2_ASAP7_75t_L g825 ( .A1(n_94), .A2(n_826), .B1(n_827), .B2(n_850), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_94), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_95), .A2(n_261), .B1(n_453), .B2(n_573), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_96), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_98), .A2(n_293), .B1(n_513), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_99), .A2(n_226), .B1(n_565), .B2(n_567), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_100), .A2(n_126), .B1(n_701), .B2(n_798), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_101), .Y(n_808) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_102), .A2(n_271), .B1(n_424), .B2(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g1127 ( .A(n_102), .Y(n_1127) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_103), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_104), .A2(n_108), .B1(n_560), .B2(n_562), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_105), .A2(n_192), .B1(n_639), .B2(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_107), .Y(n_1148) );
AOI22xp5_ASAP7_75t_SL g1067 ( .A1(n_109), .A2(n_217), .B1(n_609), .B2(n_630), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_110), .A2(n_315), .B1(n_622), .B2(n_734), .Y(n_1039) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_112), .A2(n_1168), .B1(n_1190), .B2(n_1191), .Y(n_1167) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_112), .Y(n_1190) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_114), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_116), .A2(n_207), .B1(n_634), .B2(n_909), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g1001 ( .A1(n_117), .A2(n_1002), .B1(n_1022), .B2(n_1023), .Y(n_1001) );
INVx1_ASAP7_75t_L g1022 ( .A(n_117), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_118), .A2(n_125), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g1131 ( .A(n_119), .Y(n_1131) );
CKINVDCx20_ASAP7_75t_R g1154 ( .A(n_120), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_121), .B(n_772), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g1076 ( .A(n_122), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_123), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_124), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_127), .A2(n_349), .B1(n_474), .B2(n_639), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_128), .A2(n_371), .B1(n_625), .B2(n_707), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_129), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_130), .A2(n_205), .B1(n_613), .B2(n_939), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_131), .B(n_633), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_132), .A2(n_346), .B1(n_513), .B2(n_602), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g928 ( .A1(n_133), .A2(n_216), .B1(n_929), .B2(n_930), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_134), .A2(n_375), .B1(n_560), .B2(n_610), .Y(n_1109) );
AOI22xp33_ASAP7_75t_SL g847 ( .A1(n_135), .A2(n_286), .B1(n_514), .B2(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g1139 ( .A(n_136), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_137), .A2(n_151), .B1(n_503), .B2(n_543), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_138), .A2(n_194), .B1(n_434), .B2(n_602), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_139), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g1172 ( .A(n_140), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_141), .A2(n_351), .B1(n_606), .B2(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_142), .A2(n_254), .B1(n_474), .B2(n_486), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_143), .A2(n_260), .B1(n_504), .B2(n_837), .Y(n_907) );
AOI22xp33_ASAP7_75t_SL g1053 ( .A1(n_144), .A2(n_360), .B1(n_503), .B2(n_671), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_145), .A2(n_212), .B1(n_567), .B2(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_146), .A2(n_165), .B1(n_699), .B2(n_756), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_147), .A2(n_199), .B1(n_633), .B2(n_634), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_148), .A2(n_376), .B1(n_610), .B2(n_626), .Y(n_1092) );
XNOR2x2_ASAP7_75t_L g616 ( .A(n_149), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_150), .A2(n_163), .B1(n_732), .B2(n_756), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_152), .A2(n_222), .B1(n_560), .B2(n_976), .C(n_978), .Y(n_975) );
INVx1_ASAP7_75t_L g527 ( .A(n_153), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_155), .B(n_471), .Y(n_812) );
AND2x6_ASAP7_75t_L g401 ( .A(n_156), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_156), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_159), .A2(n_385), .B1(n_462), .B2(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_160), .A2(n_196), .B1(n_521), .B2(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g927 ( .A(n_161), .B(n_663), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_162), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_164), .A2(n_367), .B1(n_453), .B2(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_166), .A2(n_200), .B1(n_418), .B2(n_434), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g926 ( .A(n_167), .B(n_790), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g1100 ( .A1(n_168), .A2(n_280), .B1(n_590), .B2(n_641), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_169), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g1137 ( .A(n_170), .Y(n_1137) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_171), .A2(n_644), .B1(n_673), .B2(n_674), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_171), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_172), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_173), .B(n_507), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_174), .Y(n_1150) );
AOI222xp33_ASAP7_75t_L g640 ( .A1(n_175), .A2(n_215), .B1(n_356), .B2(n_482), .C1(n_641), .C2(n_642), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_177), .A2(n_320), .B1(n_732), .B2(n_965), .Y(n_964) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_178), .A2(n_262), .B1(n_424), .B2(n_425), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g1128 ( .A(n_178), .B(n_1129), .Y(n_1128) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_179), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_180), .Y(n_900) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_181), .A2(n_306), .B1(n_455), .B2(n_614), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_182), .A2(n_204), .B1(n_418), .B2(n_562), .C(n_984), .Y(n_983) );
AOI22xp33_ASAP7_75t_SL g1088 ( .A1(n_183), .A2(n_190), .B1(n_573), .B2(n_625), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_184), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_187), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_188), .A2(n_210), .B1(n_453), .B2(n_521), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_189), .A2(n_198), .B1(n_634), .B2(n_909), .Y(n_1103) );
AOI22xp33_ASAP7_75t_SL g1089 ( .A1(n_191), .A2(n_341), .B1(n_753), .B2(n_896), .Y(n_1089) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_193), .A2(n_208), .B1(n_451), .B2(n_562), .C(n_646), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_195), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_201), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_202), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g1184 ( .A(n_209), .Y(n_1184) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_218), .A2(n_399), .B(n_407), .C(n_1132), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_219), .A2(n_252), .B1(n_699), .B2(n_701), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_221), .A2(n_244), .B1(n_444), .B2(n_522), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_224), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_225), .A2(n_249), .B1(n_462), .B2(n_654), .C(n_655), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_227), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_228), .A2(n_353), .B1(n_752), .B2(n_753), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_229), .A2(n_250), .B1(n_459), .B2(n_462), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_230), .A2(n_357), .B1(n_661), .B2(n_1010), .Y(n_1009) );
NAND2xp5_ASAP7_75t_SL g1057 ( .A(n_232), .B(n_663), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_233), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g986 ( .A(n_234), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_235), .A2(n_276), .B1(n_524), .B2(n_525), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_236), .A2(n_289), .B1(n_766), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_239), .A2(n_323), .B1(n_604), .B2(n_606), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_240), .Y(n_592) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_242), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_242), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_243), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_246), .A2(n_265), .B1(n_513), .B2(n_1032), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g1158 ( .A(n_247), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_248), .A2(n_344), .B1(n_562), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g1084 ( .A(n_255), .Y(n_1084) );
CKINVDCx20_ASAP7_75t_R g1052 ( .A(n_256), .Y(n_1052) );
INVx2_ASAP7_75t_L g406 ( .A(n_258), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g1176 ( .A(n_263), .Y(n_1176) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_269), .Y(n_690) );
XNOR2x1_ASAP7_75t_L g780 ( .A(n_270), .B(n_781), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_273), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_274), .A2(n_744), .B1(n_774), .B2(n_775), .Y(n_743) );
INVx1_ASAP7_75t_L g774 ( .A(n_274), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_275), .Y(n_948) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_278), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_279), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_282), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g1178 ( .A(n_284), .Y(n_1178) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_285), .Y(n_761) );
OA22x2_ASAP7_75t_L g1093 ( .A1(n_287), .A2(n_1094), .B1(n_1095), .B2(n_1111), .Y(n_1093) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_287), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_290), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_291), .A2(n_310), .B1(n_517), .B2(n_749), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_292), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_295), .Y(n_595) );
OA22x2_ASAP7_75t_L g709 ( .A1(n_296), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_296), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_297), .B(n_663), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_298), .A2(n_368), .B1(n_441), .B2(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g424 ( .A(n_299), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_299), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g1082 ( .A(n_300), .Y(n_1082) );
CKINVDCx20_ASAP7_75t_R g1183 ( .A(n_302), .Y(n_1183) );
CKINVDCx20_ASAP7_75t_R g1173 ( .A(n_303), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_304), .A2(n_354), .B1(n_604), .B2(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_305), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g1155 ( .A1(n_307), .A2(n_396), .B1(n_634), .B2(n_663), .C(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_308), .A2(n_345), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_309), .A2(n_383), .B1(n_570), .B2(n_613), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g1133 ( .A1(n_312), .A2(n_1134), .B1(n_1161), .B2(n_1162), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_312), .Y(n_1161) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_314), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_318), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_319), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_321), .Y(n_947) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_322), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_324), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_325), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_326), .A2(n_918), .B1(n_919), .B2(n_941), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_326), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_327), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_328), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_329), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_330), .A2(n_374), .B1(n_473), .B2(n_477), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_332), .Y(n_1020) );
INVx1_ASAP7_75t_L g405 ( .A(n_334), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_335), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_336), .Y(n_588) );
INVx1_ASAP7_75t_L g402 ( .A(n_337), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_338), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_340), .Y(n_532) );
XOR2x2_ASAP7_75t_L g577 ( .A(n_347), .B(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_350), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g1180 ( .A(n_352), .Y(n_1180) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_358), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g1152 ( .A(n_359), .Y(n_1152) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_361), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_362), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_363), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_364), .A2(n_397), .B1(n_467), .B2(n_470), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_366), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_369), .A2(n_377), .B1(n_629), .B2(n_630), .Y(n_628) );
XNOR2x1_ASAP7_75t_L g528 ( .A(n_370), .B(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_372), .A2(n_392), .B1(n_622), .B2(n_753), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_373), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_381), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g1157 ( .A(n_382), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_384), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_387), .B(n_543), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_388), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_389), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_391), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_393), .B(n_1056), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_394), .Y(n_956) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_402), .Y(n_1123) );
OA21x2_ASAP7_75t_L g1197 ( .A1(n_403), .A2(n_1122), .B(n_1198), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_970), .B1(n_1117), .B2(n_1118), .C(n_1119), .Y(n_407) );
INVx1_ASAP7_75t_L g1118 ( .A(n_408), .Y(n_1118) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_677), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_574), .B1(n_675), .B2(n_676), .Y(n_409) );
INVx1_ASAP7_75t_L g676 ( .A(n_410), .Y(n_676) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AO22x1_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_492), .B2(n_493), .Y(n_412) );
AO22x1_ASAP7_75t_L g915 ( .A1(n_413), .A2(n_414), .B1(n_916), .B2(n_917), .Y(n_915) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
NOR4xp75_ASAP7_75t_L g415 ( .A(n_416), .B(n_449), .C(n_465), .D(n_480), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_417), .B(n_440), .Y(n_416) );
INVx2_ASAP7_75t_L g648 ( .A(n_418), .Y(n_648) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g630 ( .A(n_419), .Y(n_630) );
INVx3_ASAP7_75t_L g798 ( .A(n_419), .Y(n_798) );
INVx2_ASAP7_75t_L g965 ( .A(n_419), .Y(n_965) );
INVx6_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g521 ( .A(n_420), .Y(n_521) );
BUFx3_ASAP7_75t_L g573 ( .A(n_420), .Y(n_573) );
BUFx3_ASAP7_75t_L g707 ( .A(n_420), .Y(n_707) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_430), .Y(n_420) );
AND2x2_ASAP7_75t_L g452 ( .A(n_421), .B(n_438), .Y(n_452) );
AND2x6_ASAP7_75t_L g455 ( .A(n_421), .B(n_456), .Y(n_455) );
AND2x6_ASAP7_75t_L g483 ( .A(n_421), .B(n_479), .Y(n_483) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g461 ( .A(n_422), .B(n_428), .Y(n_461) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g436 ( .A(n_423), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_423), .B(n_428), .Y(n_448) );
AND2x2_ASAP7_75t_L g476 ( .A(n_423), .B(n_433), .Y(n_476) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_426), .Y(n_429) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g437 ( .A(n_428), .Y(n_437) );
INVx1_ASAP7_75t_L g489 ( .A(n_428), .Y(n_489) );
AND2x2_ASAP7_75t_L g443 ( .A(n_430), .B(n_436), .Y(n_443) );
AND2x6_ASAP7_75t_L g471 ( .A(n_430), .B(n_461), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_430), .B(n_461), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_430), .B(n_436), .Y(n_658) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx2_ASAP7_75t_L g439 ( .A(n_431), .Y(n_439) );
INVx1_ASAP7_75t_L g447 ( .A(n_431), .Y(n_447) );
OR2x2_ASAP7_75t_L g457 ( .A(n_431), .B(n_432), .Y(n_457) );
AND2x2_ASAP7_75t_L g479 ( .A(n_431), .B(n_433), .Y(n_479) );
AND2x2_ASAP7_75t_L g438 ( .A(n_432), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g841 ( .A(n_434), .Y(n_841) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g513 ( .A(n_435), .Y(n_513) );
BUFx3_ASAP7_75t_L g614 ( .A(n_435), .Y(n_614) );
BUFx3_ASAP7_75t_L g705 ( .A(n_435), .Y(n_705) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_436), .B(n_438), .Y(n_652) );
INVx1_ASAP7_75t_L g478 ( .A(n_437), .Y(n_478) );
AND2x4_ASAP7_75t_L g460 ( .A(n_438), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g463 ( .A(n_438), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g526 ( .A(n_439), .Y(n_526) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_441), .Y(n_752) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx5_ASAP7_75t_L g522 ( .A(n_442), .Y(n_522) );
BUFx3_ASAP7_75t_L g566 ( .A(n_442), .Y(n_566) );
INVx4_ASAP7_75t_L g605 ( .A(n_442), .Y(n_605) );
INVx3_ASAP7_75t_L g622 ( .A(n_442), .Y(n_622) );
INVx1_ASAP7_75t_L g844 ( .A(n_442), .Y(n_844) );
INVx8_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx4f_ASAP7_75t_SL g661 ( .A(n_445), .Y(n_661) );
BUFx2_ASAP7_75t_L g734 ( .A(n_445), .Y(n_734) );
BUFx2_ASAP7_75t_L g845 ( .A(n_445), .Y(n_845) );
BUFx2_ASAP7_75t_L g988 ( .A(n_445), .Y(n_988) );
INVx6_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g567 ( .A(n_446), .Y(n_567) );
INVx1_ASAP7_75t_L g606 ( .A(n_446), .Y(n_606) );
INVx1_ASAP7_75t_SL g753 ( .A(n_446), .Y(n_753) );
OR2x6_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g475 ( .A(n_447), .Y(n_475) );
INVx1_ASAP7_75t_L g464 ( .A(n_448), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_450), .B(n_458), .Y(n_449) );
INVx1_ASAP7_75t_L g1153 ( .A(n_451), .Y(n_1153) );
BUFx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
INVx2_ASAP7_75t_L g700 ( .A(n_452), .Y(n_700) );
BUFx2_ASAP7_75t_SL g1062 ( .A(n_452), .Y(n_1062) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_SL g609 ( .A(n_454), .Y(n_609) );
INVx3_ASAP7_75t_L g654 ( .A(n_454), .Y(n_654) );
INVx4_ASAP7_75t_L g874 ( .A(n_454), .Y(n_874) );
INVx11_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx11_ASAP7_75t_L g518 ( .A(n_455), .Y(n_518) );
AND2x4_ASAP7_75t_L g469 ( .A(n_456), .B(n_461), .Y(n_469) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g534 ( .A(n_457), .B(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g756 ( .A(n_459), .Y(n_756) );
BUFx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_460), .Y(n_524) );
BUFx3_ASAP7_75t_L g611 ( .A(n_460), .Y(n_611) );
BUFx3_ASAP7_75t_L g701 ( .A(n_460), .Y(n_701) );
INVx2_ASAP7_75t_L g877 ( .A(n_460), .Y(n_877) );
INVx1_ASAP7_75t_L g535 ( .A(n_461), .Y(n_535) );
INVx1_ASAP7_75t_L g982 ( .A(n_462), .Y(n_982) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g514 ( .A(n_463), .Y(n_514) );
INVx1_ASAP7_75t_L g571 ( .A(n_463), .Y(n_571) );
BUFx2_ASAP7_75t_SL g602 ( .A(n_463), .Y(n_602) );
BUFx3_ASAP7_75t_L g620 ( .A(n_463), .Y(n_620) );
BUFx2_ASAP7_75t_SL g749 ( .A(n_463), .Y(n_749) );
BUFx2_ASAP7_75t_L g935 ( .A(n_463), .Y(n_935) );
BUFx3_ASAP7_75t_L g1141 ( .A(n_463), .Y(n_1141) );
AND2x2_ASAP7_75t_L g525 ( .A(n_464), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_472), .Y(n_465) );
BUFx2_ASAP7_75t_L g990 ( .A(n_467), .Y(n_990) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g507 ( .A(n_468), .Y(n_507) );
INVx5_ASAP7_75t_L g633 ( .A(n_468), .Y(n_633) );
INVx2_ASAP7_75t_L g909 ( .A(n_468), .Y(n_909) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g635 ( .A(n_471), .Y(n_635) );
BUFx2_ASAP7_75t_L g790 ( .A(n_471), .Y(n_790) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g638 ( .A(n_474), .Y(n_638) );
BUFx2_ASAP7_75t_L g763 ( .A(n_474), .Y(n_763) );
BUFx2_ASAP7_75t_L g837 ( .A(n_474), .Y(n_837) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x4_ASAP7_75t_L g487 ( .A(n_476), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g490 ( .A(n_476), .B(n_491), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_476), .B(n_526), .Y(n_550) );
BUFx3_ASAP7_75t_L g504 ( .A(n_477), .Y(n_504) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_477), .Y(n_639) );
BUFx2_ASAP7_75t_SL g786 ( .A(n_477), .Y(n_786) );
BUFx2_ASAP7_75t_SL g1059 ( .A(n_477), .Y(n_1059) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
INVx1_ASAP7_75t_L g555 ( .A(n_479), .Y(n_555) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_484), .B(n_485), .Y(n_480) );
OAI21xp33_ASAP7_75t_SL g720 ( .A1(n_481), .A2(n_721), .B(n_722), .Y(n_720) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g501 ( .A(n_483), .Y(n_501) );
INVx4_ASAP7_75t_L g670 ( .A(n_483), .Y(n_670) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_483), .Y(n_769) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_483), .Y(n_1080) );
INVx2_ASAP7_75t_L g1098 ( .A(n_483), .Y(n_1098) );
BUFx6f_ASAP7_75t_L g997 ( .A(n_486), .Y(n_997) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
BUFx2_ASAP7_75t_L g641 ( .A(n_487), .Y(n_641) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_487), .Y(n_766) );
BUFx4f_ASAP7_75t_SL g902 ( .A(n_487), .Y(n_902) );
INVx1_ASAP7_75t_L g491 ( .A(n_489), .Y(n_491) );
BUFx12f_ASAP7_75t_L g503 ( .A(n_490), .Y(n_503) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_490), .Y(n_545) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_490), .Y(n_591) );
INVx1_ASAP7_75t_L g904 ( .A(n_490), .Y(n_904) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
XNOR2x1_ASAP7_75t_SL g493 ( .A(n_494), .B(n_528), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_527), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_498), .B(n_510), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_502), .Y(n_499) );
OAI21xp33_ASAP7_75t_SL g540 ( .A1(n_501), .A2(n_541), .B(n_542), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_501), .A2(n_588), .B1(n_589), .B2(n_592), .C(n_593), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g859 ( .A1(n_501), .A2(n_860), .B(n_861), .Y(n_859) );
BUFx4f_ASAP7_75t_SL g642 ( .A(n_503), .Y(n_642) );
INVx2_ASAP7_75t_L g725 ( .A(n_503), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .C(n_509), .Y(n_505) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx3_ASAP7_75t_L g561 ( .A(n_516), .Y(n_561) );
BUFx3_ASAP7_75t_L g625 ( .A(n_516), .Y(n_625) );
BUFx3_ASAP7_75t_L g894 ( .A(n_516), .Y(n_894) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_516), .Y(n_939) );
INVx1_ASAP7_75t_L g891 ( .A(n_517), .Y(n_891) );
INVx5_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g629 ( .A(n_518), .Y(n_629) );
INVx2_ASAP7_75t_L g732 ( .A(n_518), .Y(n_732) );
INVx1_ASAP7_75t_L g848 ( .A(n_518), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
BUFx2_ASAP7_75t_L g871 ( .A(n_522), .Y(n_871) );
BUFx6f_ASAP7_75t_L g1010 ( .A(n_522), .Y(n_1010) );
INVx4_ASAP7_75t_L g563 ( .A(n_524), .Y(n_563) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_557), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .C(n_546), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_536), .B2(n_537), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_533), .A2(n_538), .B1(n_689), .B2(n_690), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_533), .A2(n_949), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g583 ( .A(n_534), .Y(n_583) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_534), .Y(n_717) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_537), .A2(n_715), .B1(n_718), .B2(n_719), .Y(n_714) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g586 ( .A(n_538), .Y(n_586) );
OAI22xp5_ASAP7_75t_SL g1074 ( .A1(n_538), .A2(n_717), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g868 ( .A(n_539), .Y(n_868) );
INVx4_ASAP7_75t_L g672 ( .A(n_543), .Y(n_672) );
BUFx2_ASAP7_75t_L g723 ( .A(n_543), .Y(n_723) );
INVx1_ASAP7_75t_L g833 ( .A(n_544), .Y(n_833) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_551), .B2(n_552), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_548), .A2(n_598), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVx3_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g993 ( .A(n_549), .Y(n_993) );
INVx4_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_550), .Y(n_596) );
BUFx3_ASAP7_75t_L g666 ( .A(n_550), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_550), .A2(n_554), .B1(n_695), .B2(n_696), .Y(n_694) );
OAI22xp33_ASAP7_75t_SL g726 ( .A1(n_550), .A2(n_598), .B1(n_727), .B2(n_728), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_550), .A2(n_552), .B1(n_857), .B2(n_858), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_552), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_664) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g598 ( .A(n_553), .Y(n_598) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g995 ( .A(n_554), .Y(n_995) );
OR2x6_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_568), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .Y(n_558) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g934 ( .A(n_563), .Y(n_934) );
OAI221xp5_ASAP7_75t_SL g1182 ( .A1(n_563), .A2(n_980), .B1(n_1183), .B2(n_1184), .C(n_1185), .Y(n_1182) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_571), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g675 ( .A(n_574), .Y(n_675) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_643), .Y(n_574) );
OAI22xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_577), .B1(n_615), .B2(n_616), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_599), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_587), .C(n_594), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_584), .B2(n_585), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_582), .A2(n_947), .B1(n_948), .B2(n_949), .Y(n_946) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g1171 ( .A(n_583), .Y(n_1171) );
OAI221xp5_ASAP7_75t_SL g759 ( .A1(n_585), .A2(n_717), .B1(n_760), .B2(n_761), .C(n_762), .Y(n_759) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g950 ( .A1(n_589), .A2(n_768), .B1(n_951), .B2(n_952), .C1(n_953), .C2(n_954), .Y(n_950) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx2_ASAP7_75t_L g772 ( .A(n_591), .Y(n_772) );
INVx2_ASAP7_75t_L g863 ( .A(n_591), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_598), .A2(n_666), .B1(n_956), .B2(n_957), .Y(n_955) );
OAI22xp5_ASAP7_75t_SL g1083 ( .A1(n_598), .A2(n_666), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_607), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g897 ( .A(n_605), .Y(n_897) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_605), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .Y(n_607) );
INVx1_ASAP7_75t_L g1149 ( .A(n_609), .Y(n_1149) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx4f_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g627 ( .A(n_614), .Y(n_627) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND4xp75_ASAP7_75t_L g617 ( .A(n_618), .B(n_623), .C(n_631), .D(n_640), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g980 ( .A(n_629), .Y(n_980) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_632), .B(n_636), .Y(n_631) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_633), .Y(n_663) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_635), .Y(n_1056) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g929 ( .A(n_638), .Y(n_929) );
INVx1_ASAP7_75t_SL g931 ( .A(n_639), .Y(n_931) );
INVx1_ASAP7_75t_L g951 ( .A(n_641), .Y(n_951) );
INVx1_ASAP7_75t_L g1179 ( .A(n_642), .Y(n_1179) );
INVx1_ASAP7_75t_L g674 ( .A(n_644), .Y(n_674) );
AND4x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_653), .C(n_662), .D(n_668), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_648), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_648), .A2(n_1148), .B1(n_1149), .B2(n_1150), .Y(n_1147) );
OAI221xp5_ASAP7_75t_SL g746 ( .A1(n_650), .A2(n_747), .B1(n_748), .B2(n_750), .C(n_751), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_650), .A2(n_1152), .B1(n_1153), .B2(n_1154), .Y(n_1151) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g738 ( .A(n_651), .Y(n_738) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_657), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_657), .A2(n_1143), .B1(n_1144), .B2(n_1145), .Y(n_1142) );
BUFx2_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g1177 ( .A(n_669), .Y(n_1177) );
INVx4_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g783 ( .A1(n_670), .A2(n_784), .B(n_785), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_670), .A2(n_808), .B(n_809), .Y(n_807) );
BUFx2_ASAP7_75t_L g830 ( .A(n_670), .Y(n_830) );
OAI21xp5_ASAP7_75t_SL g1051 ( .A1(n_670), .A2(n_1052), .B(n_1053), .Y(n_1051) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_820), .Y(n_677) );
OAI22xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_777), .B1(n_778), .B2(n_819), .Y(n_678) );
INVx2_ASAP7_75t_L g819 ( .A(n_679), .Y(n_819) );
AO22x2_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B1(n_743), .B2(n_776), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_708), .B2(n_709), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND3x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_697), .C(n_703), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .C(n_694), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_702), .Y(n_697) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g1032 ( .A(n_700), .Y(n_1032) );
INVx1_ASAP7_75t_L g741 ( .A(n_701), .Y(n_741) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g977 ( .A(n_705), .Y(n_977) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_705), .Y(n_1189) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
XNOR2x2_ASAP7_75t_L g778 ( .A(n_709), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_729), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_720), .C(n_726), .Y(n_713) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_717), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
INVx3_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_735), .C(n_739), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx2_ASAP7_75t_L g776 ( .A(n_743), .Y(n_776) );
INVx1_ASAP7_75t_L g775 ( .A(n_744), .Y(n_775) );
AND2x2_ASAP7_75t_SL g744 ( .A(n_745), .B(n_758), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_754), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g1138 ( .A(n_756), .Y(n_1138) );
NOR2xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_764), .Y(n_758) );
OAI222xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B1(n_768), .B2(n_770), .C1(n_771), .C2(n_773), .Y(n_764) );
OAI222xp33_ASAP7_75t_L g829 ( .A1(n_765), .A2(n_830), .B1(n_831), .B2(n_832), .C1(n_833), .C2(n_834), .Y(n_829) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_765), .A2(n_830), .B1(n_1016), .B2(n_1017), .C(n_1018), .Y(n_1015) );
OAI222xp33_ASAP7_75t_L g1175 ( .A1(n_765), .A2(n_1176), .B1(n_1177), .B2(n_1178), .C1(n_1179), .C2(n_1180), .Y(n_1175) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
OAI222xp33_ASAP7_75t_L g899 ( .A1(n_768), .A2(n_900), .B1(n_901), .B2(n_903), .C1(n_904), .C2(n_905), .Y(n_899) );
INVx2_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g922 ( .A(n_769), .Y(n_922) );
INVxp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI22x1_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_800), .B1(n_801), .B2(n_818), .Y(n_779) );
INVx2_ASAP7_75t_L g818 ( .A(n_780), .Y(n_818) );
AND2x4_ASAP7_75t_L g781 ( .A(n_782), .B(n_792), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .C(n_791), .Y(n_787) );
NOR2x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_796), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_800), .A2(n_801), .B1(n_882), .B2(n_883), .Y(n_881) );
INVx3_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
XOR2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_817), .Y(n_801) );
NAND3x1_ASAP7_75t_SL g802 ( .A(n_803), .B(n_806), .C(n_814), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
NOR2x1_ASAP7_75t_L g806 ( .A(n_807), .B(n_810), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .C(n_813), .Y(n_810) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_911), .B1(n_912), .B2(n_969), .Y(n_820) );
INVx1_ASAP7_75t_L g969 ( .A(n_821), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .B1(n_879), .B2(n_880), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B1(n_851), .B2(n_852), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g850 ( .A(n_827), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_839), .C(n_846), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_835), .Y(n_828) );
INVx1_ASAP7_75t_L g1160 ( .A(n_830), .Y(n_1160) );
OAI222xp33_ASAP7_75t_L g1077 ( .A1(n_833), .A2(n_1078), .B1(n_1079), .B2(n_1080), .C1(n_1081), .C2(n_1082), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_838), .Y(n_835) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_842), .Y(n_839) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVxp67_ASAP7_75t_L g1145 ( .A(n_845), .Y(n_1145) );
AND2x2_ASAP7_75t_L g846 ( .A(n_847), .B(n_849), .Y(n_846) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g878 ( .A(n_854), .Y(n_878) );
NAND2x1_ASAP7_75t_L g854 ( .A(n_855), .B(n_869), .Y(n_854) );
NOR3xp33_ASAP7_75t_SL g855 ( .A(n_856), .B(n_859), .C(n_864), .Y(n_855) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
OA211x2_ASAP7_75t_L g1033 ( .A1(n_867), .A2(n_1034), .B(n_1035), .C(n_1036), .Y(n_1033) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g949 ( .A(n_868), .Y(n_949) );
AND4x1_ASAP7_75t_L g869 ( .A(n_870), .B(n_872), .C(n_873), .D(n_875), .Y(n_869) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g961 ( .A(n_877), .Y(n_961) );
INVx1_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g910 ( .A(n_885), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_898), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_892), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_895), .Y(n_892) );
INVx3_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_906), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
BUFx3_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_942), .B2(n_943), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g941 ( .A(n_919), .Y(n_941) );
NAND3x1_ASAP7_75t_L g919 ( .A(n_920), .B(n_932), .C(n_937), .Y(n_919) );
NOR2x1_ASAP7_75t_L g920 ( .A(n_921), .B(n_925), .Y(n_920) );
OAI21xp5_ASAP7_75t_SL g921 ( .A1(n_922), .A2(n_923), .B(n_924), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .C(n_928), .Y(n_925) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
AND2x2_ASAP7_75t_L g932 ( .A(n_933), .B(n_936), .Y(n_932) );
AND2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_940), .Y(n_937) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_SL g968 ( .A(n_944), .Y(n_968) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_958), .Y(n_944) );
NOR3xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_950), .C(n_955), .Y(n_945) );
OAI221xp5_ASAP7_75t_SL g1170 ( .A1(n_949), .A2(n_1171), .B1(n_1172), .B2(n_1173), .C(n_1174), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_963), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_960), .B(n_962), .Y(n_959) );
NAND2xp5_ASAP7_75t_SL g963 ( .A(n_964), .B(n_966), .Y(n_963) );
INVx1_ASAP7_75t_L g1117 ( .A(n_970), .Y(n_1117) );
AOI22xp5_ASAP7_75t_SL g970 ( .A1(n_971), .A2(n_972), .B1(n_1045), .B2(n_1116), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_1000), .B1(n_1043), .B2(n_1044), .Y(n_972) );
INVx1_ASAP7_75t_L g1043 ( .A(n_973), .Y(n_1043) );
INVx1_ASAP7_75t_L g999 ( .A(n_974), .Y(n_999) );
AND4x2_ASAP7_75t_L g974 ( .A(n_975), .B(n_983), .C(n_989), .D(n_996), .Y(n_974) );
INVx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_980), .B1(n_981), .B2(n_982), .Y(n_978) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_993), .A2(n_995), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
INVx2_ASAP7_75t_SL g1078 ( .A(n_997), .Y(n_1078) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1000), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1024), .B1(n_1025), .B2(n_1042), .Y(n_1000) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1001), .Y(n_1042) );
INVx1_ASAP7_75t_SL g1023 ( .A(n_1002), .Y(n_1023) );
AND2x2_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1011), .Y(n_1002) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
NOR3xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1015), .C(n_1019), .Y(n_1011) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
XOR2x2_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1041), .Y(n_1027) );
NAND4xp75_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1033), .C(n_1037), .D(n_1040), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1045), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1069), .B1(n_1114), .B2(n_1115), .Y(n_1046) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1047), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
XOR2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1068), .Y(n_1048) );
NAND3x1_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1060), .C(n_1065), .Y(n_1049) );
NOR2x1_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1054), .Y(n_1050) );
NAND3xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1057), .C(n_1058), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1063), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1069), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1093), .B1(n_1112), .B2(n_1113), .Y(n_1069) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1070), .Y(n_1112) );
XNOR2x2_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1086), .Y(n_1072) );
NOR3xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1077), .C(n_1083), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1090), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1092), .Y(n_1090) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1093), .Y(n_1113) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1095), .Y(n_1111) );
NAND2x1_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1104), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1101), .Y(n_1096) );
OAI21xp5_ASAP7_75t_SL g1097 ( .A1(n_1098), .A2(n_1099), .B(n_1100), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1103), .Y(n_1101) );
NOR2x1_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1108), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
INVx1_ASAP7_75t_SL g1119 ( .A(n_1120), .Y(n_1119) );
NOR2x1_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1125), .Y(n_1120) );
OR2x2_ASAP7_75t_SL g1194 ( .A(n_1121), .B(n_1126), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1124), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1122), .B(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1123), .B(n_1164), .Y(n_1198) );
CKINVDCx16_ASAP7_75t_R g1164 ( .A(n_1124), .Y(n_1164) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_1126), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1128), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1131), .Y(n_1129) );
OAI222xp33_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1163), .B1(n_1165), .B2(n_1190), .C1(n_1192), .C2(n_1195), .Y(n_1132) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1134), .Y(n_1162) );
AND4x1_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1146), .C(n_1155), .D(n_1159), .Y(n_1134) );
NOR2xp33_ASAP7_75t_SL g1135 ( .A(n_1136), .B(n_1142), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1138), .B1(n_1139), .B2(n_1140), .Y(n_1136) );
INVxp67_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1151), .Y(n_1146) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_SL g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1168), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1181), .Y(n_1168) );
NOR2xp33_ASAP7_75t_SL g1169 ( .A(n_1170), .B(n_1175), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1186), .Y(n_1181) );
NAND2xp33_ASAP7_75t_SL g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
CKINVDCx20_ASAP7_75t_R g1192 ( .A(n_1193), .Y(n_1192) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
CKINVDCx20_ASAP7_75t_R g1196 ( .A(n_1197), .Y(n_1196) );
endmodule