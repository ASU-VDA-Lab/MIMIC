module fake_jpeg_4302_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_26),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_13),
.B1(n_19),
.B2(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_13),
.B1(n_25),
.B2(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_11),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_17),
.C(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_33),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_43),
.B1(n_14),
.B2(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_13),
.B1(n_19),
.B2(n_18),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_18),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_16),
.C(n_12),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_48),
.B1(n_44),
.B2(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_51),
.B1(n_41),
.B2(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_50),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_9),
.B2(n_8),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_36),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_58),
.B(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_57),
.B1(n_8),
.B2(n_9),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_65),
.B1(n_56),
.B2(n_53),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.C(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_52),
.C(n_44),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_2),
.C(n_3),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_68),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_63),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_55),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_61),
.C(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_69),
.B(n_3),
.C(n_4),
.Y(n_74)
);

OAI31xp33_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_2),
.A3(n_4),
.B(n_5),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_70),
.B(n_4),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_6),
.Y(n_78)
);


endmodule