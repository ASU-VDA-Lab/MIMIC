module fake_ariane_1409_n_1909 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1909);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1909;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_24),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_19),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_98),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_20),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_83),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_14),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_73),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_29),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_174),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_58),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_18),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_31),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_80),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_173),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_77),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_107),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_132),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_122),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_32),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_187),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_139),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_118),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_45),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_87),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_11),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_127),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_91),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_167),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_59),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_30),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_33),
.Y(n_246)
);

BUFx2_ASAP7_75t_SL g247 ( 
.A(n_6),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_119),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_46),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_48),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_143),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_35),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_144),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_33),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_56),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_185),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_178),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_181),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_53),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_89),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_147),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_94),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_166),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_61),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_76),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_161),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_70),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_123),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_146),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_153),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_141),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_138),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_192),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_114),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_97),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_115),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_51),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_110),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_4),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_60),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_67),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_47),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_5),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_164),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_68),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_101),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_9),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_95),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_102),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_75),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_99),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_177),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_112),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_84),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_191),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_85),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_96),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_42),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_176),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_50),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_186),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_162),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_39),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_105),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_46),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_142),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_19),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_180),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_3),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_184),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_109),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_92),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_134),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_74),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_44),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_125),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_128),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_18),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_2),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_108),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_182),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_106),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_15),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_57),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_64),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_39),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_169),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_163),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_155),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_21),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_78),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_121),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_21),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_158),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_5),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_23),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_154),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_50),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_103),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_11),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_15),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_10),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_28),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_145),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_40),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_100),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_3),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_63),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_34),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_159),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_27),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_71),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_47),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_62),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_7),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_10),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_25),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_129),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_130),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_82),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_41),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_148),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_41),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_117),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_9),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_120),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_43),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_382),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_216),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_243),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_243),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_200),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_379),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_193),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_379),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_209),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_211),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_253),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_222),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_258),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_262),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_263),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_273),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_297),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_303),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_276),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_194),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_367),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_247),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_371),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_207),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_228),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_358),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_223),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_227),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_193),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_228),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_206),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_206),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_287),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_194),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_309),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_276),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_206),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_374),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_383),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_246),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_246),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_219),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_269),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_269),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_276),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_219),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_276),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_195),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_346),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_197),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_195),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_219),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_276),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_288),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_236),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_354),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_288),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_288),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_199),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_288),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_366),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_238),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_236),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_288),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_236),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_316),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_316),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_240),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_316),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_245),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_197),
.Y(n_466)
);

BUFx2_ASAP7_75t_SL g467 ( 
.A(n_218),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_218),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_369),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_196),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_198),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_204),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_199),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_210),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_310),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_214),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_231),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_198),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_239),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_201),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_390),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_412),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_298),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_413),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_310),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_202),
.B1(n_381),
.B2(n_230),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_456),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g497 ( 
.A1(n_451),
.A2(n_244),
.B(n_241),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_439),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_452),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_454),
.Y(n_501)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_458),
.A2(n_264),
.B(n_252),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_473),
.B(n_315),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_475),
.B(n_315),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_446),
.A2(n_271),
.B(n_268),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_468),
.B(n_477),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_372),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_447),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_416),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_480),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_417),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_426),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_468),
.B(n_278),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_419),
.B(n_228),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_431),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_419),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_476),
.B(n_372),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_434),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_419),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_393),
.B(n_280),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_442),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_421),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_387),
.Y(n_533)
);

OAI21xp33_ASAP7_75t_L g534 ( 
.A1(n_394),
.A2(n_397),
.B(n_395),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_388),
.B(n_330),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_462),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_445),
.B(n_250),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_406),
.B(n_250),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_399),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_389),
.B(n_330),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_391),
.B(n_201),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_400),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_444),
.B(n_281),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_449),
.B(n_289),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_402),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_403),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_405),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_410),
.B(n_414),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_415),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_387),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_R g561 ( 
.A(n_484),
.B(n_422),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_559),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_493),
.A2(n_386),
.B1(n_418),
.B2(n_392),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_520),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_460),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_559),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_517),
.B(n_406),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_R g570 ( 
.A(n_516),
.B(n_424),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_528),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_486),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_517),
.B(n_482),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_508),
.A2(n_362),
.B(n_320),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_500),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_498),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_538),
.B(n_423),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_484),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_498),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_506),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_538),
.B(n_423),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_485),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_539),
.A2(n_392),
.B1(n_418),
.B2(n_453),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_504),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_499),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_538),
.B(n_443),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_536),
.B(n_463),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_499),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_501),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_552),
.B(n_466),
.C(n_443),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_536),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_539),
.B(n_466),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_490),
.B(n_465),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_500),
.Y(n_598)
);

OAI21xp33_ASAP7_75t_SL g599 ( 
.A1(n_542),
.A2(n_453),
.B(n_469),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_507),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_506),
.B(n_472),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_538),
.B(n_472),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_515),
.B(n_470),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_523),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_552),
.B(n_479),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_537),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_542),
.A2(n_386),
.B1(n_479),
.B2(n_481),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_537),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_535),
.A2(n_360),
.B1(n_248),
.B2(n_481),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_507),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_540),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_536),
.B(n_409),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_540),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_509),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_506),
.B(n_224),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_530),
.B(n_320),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_540),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_535),
.A2(n_461),
.B1(n_459),
.B2(n_457),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_543),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_543),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_512),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_542),
.A2(n_212),
.B1(n_203),
.B2(n_202),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_512),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_506),
.B(n_235),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g630 ( 
.A1(n_508),
.A2(n_384),
.B(n_362),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_513),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_511),
.A2(n_275),
.B1(n_270),
.B2(n_267),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_501),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_513),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_528),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_545),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_545),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_528),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_528),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_523),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_528),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_528),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_545),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_485),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_528),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_488),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_506),
.B(n_259),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_545),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_488),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_547),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_545),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_547),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_488),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_489),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_523),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_489),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_558),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_514),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_558),
.Y(n_662)
);

BUFx6f_ASAP7_75t_SL g663 ( 
.A(n_511),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_496),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_547),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_496),
.B(n_441),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_558),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_557),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_493),
.A2(n_348),
.B1(n_342),
.B2(n_291),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_492),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_384),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_487),
.B(n_455),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_511),
.A2(n_327),
.B1(n_257),
.B2(n_255),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_548),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_557),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_489),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_532),
.B(n_203),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_494),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_487),
.B(n_284),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_396),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_532),
.A2(n_291),
.B1(n_230),
.B2(n_221),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_511),
.B(n_286),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_515),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_530),
.B(n_420),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_492),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_557),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_494),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_557),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_520),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_515),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_547),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_547),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_547),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_524),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_547),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_524),
.B(n_420),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_524),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_550),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_550),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_550),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_524),
.B(n_427),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_524),
.B(n_427),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_490),
.B(n_212),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_494),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_503),
.B(n_296),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_495),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_548),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_535),
.A2(n_461),
.B1(n_459),
.B2(n_457),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_495),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_522),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_503),
.B(n_302),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_550),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_679),
.B(n_503),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_563),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_684),
.B(n_433),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_564),
.Y(n_717)
);

AND2x6_ASAP7_75t_SL g718 ( 
.A(n_591),
.B(n_544),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_L g719 ( 
.A1(n_599),
.A2(n_534),
.B1(n_556),
.B2(n_555),
.C(n_553),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_595),
.B(n_551),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_595),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_577),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_573),
.B(n_672),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_694),
.B(n_505),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_618),
.A2(n_497),
.B1(n_502),
.B2(n_535),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_688),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_570),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_664),
.B(n_586),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_694),
.B(n_505),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_583),
.B(n_550),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_569),
.B(n_550),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_596),
.B(n_550),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_564),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_583),
.B(n_560),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_664),
.B(n_551),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_580),
.B(n_433),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_601),
.B(n_705),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_572),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_583),
.B(n_560),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_711),
.B(n_535),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_585),
.B(n_438),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_577),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_688),
.B(n_560),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_645),
.B(n_492),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_590),
.B(n_438),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_578),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_572),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_582),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_582),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_683),
.B(n_549),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_683),
.A2(n_534),
.B(n_556),
.C(n_555),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_579),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

AND3x1_ASAP7_75t_L g755 ( 
.A(n_587),
.B(n_551),
.C(n_546),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_617),
.B(n_549),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_591),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_688),
.B(n_560),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_584),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_581),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_636),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_448),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_614),
.B(n_448),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_697),
.B(n_636),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_629),
.B(n_553),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_SL g767 ( 
.A(n_653),
.B(n_533),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_697),
.B(n_560),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_697),
.B(n_560),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_637),
.B(n_560),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_SL g771 ( 
.A(n_608),
.B(n_342),
.C(n_221),
.Y(n_771)
);

O2A1O1Ixp5_ASAP7_75t_L g772 ( 
.A1(n_637),
.A2(n_546),
.B(n_544),
.C(n_519),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_584),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_648),
.B(n_541),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_588),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_690),
.B(n_541),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_644),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_644),
.B(n_560),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_618),
.A2(n_347),
.B1(n_510),
.B2(n_350),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_618),
.B(n_541),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_670),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_588),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_649),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_618),
.B(n_510),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_600),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_649),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_671),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_671),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_696),
.B(n_353),
.C(n_348),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_674),
.B(n_519),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_574),
.B(n_605),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_652),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_707),
.B(n_521),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_652),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_606),
.B(n_396),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_600),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_562),
.B(n_521),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_654),
.B(n_205),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_654),
.B(n_205),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_685),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_591),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_568),
.B(n_682),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_525),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_701),
.B(n_408),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_703),
.B(n_525),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_651),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_668),
.A2(n_375),
.B1(n_373),
.B2(n_365),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_703),
.B(n_526),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_675),
.B(n_208),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_611),
.Y(n_810)
);

INVx8_ASAP7_75t_L g811 ( 
.A(n_671),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_567),
.B(n_526),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_675),
.B(n_208),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_567),
.B(n_529),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_686),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_702),
.B(n_408),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_686),
.B(n_213),
.Y(n_817)
);

BUFx12f_ASAP7_75t_L g818 ( 
.A(n_581),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_591),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_597),
.B(n_529),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_578),
.B(n_598),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_589),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_597),
.B(n_531),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_611),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_613),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_574),
.B(n_605),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_668),
.B(n_531),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_598),
.B(n_213),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_671),
.B(n_497),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_626),
.B(n_215),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_661),
.B(n_554),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_594),
.B(n_411),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_626),
.B(n_215),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_671),
.B(n_497),
.Y(n_834)
);

BUFx6f_ASAP7_75t_SL g835 ( 
.A(n_604),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_671),
.B(n_497),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_651),
.B(n_217),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_677),
.B(n_411),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_680),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_602),
.B(n_497),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_607),
.B(n_502),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_613),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_565),
.A2(n_353),
.B1(n_361),
.B2(n_365),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_589),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_632),
.A2(n_361),
.B1(n_373),
.B2(n_375),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_592),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_609),
.A2(n_381),
.B(n_313),
.C(n_317),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_592),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_677),
.B(n_554),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_604),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_616),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_561),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_651),
.B(n_217),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_604),
.B(n_251),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_610),
.A2(n_502),
.B1(n_508),
.B2(n_370),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_612),
.B(n_502),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_666),
.B(n_279),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_616),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_681),
.B(n_293),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_627),
.B(n_299),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_615),
.B(n_502),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_651),
.B(n_220),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_651),
.B(n_220),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_673),
.B(n_304),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_619),
.B(n_225),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_621),
.B(n_225),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_593),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_574),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_625),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_669),
.B(n_318),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_593),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_663),
.B(n_321),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_633),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_693),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_633),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_623),
.B(n_226),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_663),
.B(n_323),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_624),
.B(n_226),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_660),
.A2(n_508),
.B1(n_334),
.B2(n_312),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_662),
.B(n_229),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_667),
.B(n_229),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_710),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_818),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_822),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_787),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_728),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_605),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_713),
.B(n_640),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_818),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_715),
.B(n_708),
.C(n_620),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_722),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_737),
.B(n_663),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_864),
.A2(n_631),
.B1(n_625),
.B2(n_628),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_852),
.Y(n_894)
);

INVx4_ASAP7_75t_SL g895 ( 
.A(n_806),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_844),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_736),
.B(n_741),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_846),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_848),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_735),
.B(n_628),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_806),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_772),
.A2(n_692),
.B(n_691),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_755),
.A2(n_658),
.B1(n_640),
.B2(n_641),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_791),
.A2(n_641),
.B(n_640),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_867),
.Y(n_906)
);

CKINVDCx8_ASAP7_75t_R g907 ( 
.A(n_718),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_774),
.B(n_658),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_802),
.B(n_658),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_742),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_749),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_871),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_839),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_756),
.B(n_631),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_726),
.B(n_655),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_721),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_870),
.A2(n_712),
.B1(n_695),
.B2(n_700),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_873),
.A2(n_634),
.B1(n_508),
.B2(n_693),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_745),
.B(n_710),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_766),
.B(n_634),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_757),
.B(n_710),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_724),
.B(n_691),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_801),
.B(n_638),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_SL g924 ( 
.A1(n_839),
.A2(n_816),
.B1(n_804),
.B2(n_795),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_729),
.B(n_692),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_859),
.A2(n_712),
.B1(n_700),
.B2(n_699),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_748),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_740),
.B(n_695),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_763),
.B(n_699),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_790),
.B(n_805),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_875),
.Y(n_931)
);

O2A1O1Ixp5_ASAP7_75t_L g932 ( 
.A1(n_837),
.A2(n_862),
.B(n_863),
.C(n_853),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_761),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_808),
.B(n_638),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_749),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_714),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_776),
.B(n_639),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_776),
.B(n_639),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_819),
.A2(n_698),
.B1(n_665),
.B2(n_655),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_849),
.B(n_325),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_800),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_776),
.B(n_642),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_751),
.B(n_642),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_744),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_750),
.Y(n_945)
);

BUFx4f_ASAP7_75t_SL g946 ( 
.A(n_761),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_726),
.B(n_655),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_771),
.A2(n_698),
.B1(n_665),
.B2(n_655),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_789),
.B(n_758),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_716),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_717),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_733),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_803),
.B(n_643),
.Y(n_953)
);

INVx8_ASAP7_75t_L g954 ( 
.A(n_811),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_850),
.A2(n_698),
.B1(n_665),
.B2(n_655),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_860),
.A2(n_646),
.B1(n_643),
.B2(n_704),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_727),
.B(n_665),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_812),
.B(n_646),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_855),
.A2(n_709),
.B1(n_706),
.B2(n_704),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_R g960 ( 
.A(n_744),
.B(n_647),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_760),
.A2(n_678),
.B1(n_706),
.B2(n_647),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_787),
.B(n_665),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_814),
.B(n_698),
.Y(n_963)
);

NAND2x1_ASAP7_75t_L g964 ( 
.A(n_787),
.B(n_698),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_820),
.B(n_571),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_720),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_788),
.B(n_868),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_823),
.B(n_571),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_788),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_760),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_835),
.A2(n_571),
.B1(n_635),
.B2(n_352),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_788),
.B(n_868),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_738),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_SL g974 ( 
.A(n_727),
.B(n_566),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_747),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_780),
.B(n_784),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_753),
.B(n_571),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_754),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_762),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_777),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_868),
.B(n_571),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_793),
.B(n_635),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_783),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_773),
.A2(n_709),
.B1(n_650),
.B2(n_687),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_744),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_797),
.B(n_635),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_781),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_826),
.A2(n_635),
.B(n_687),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_874),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_806),
.B(n_635),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_786),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_792),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_746),
.B(n_650),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_806),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_794),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_835),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_773),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_775),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_767),
.B(n_575),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_872),
.B(n_656),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_779),
.A2(n_832),
.B1(n_843),
.B2(n_877),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_815),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_775),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_782),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_854),
.B(n_656),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_764),
.B(n_657),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_811),
.B(n_575),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_838),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_811),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_730),
.A2(n_739),
.B(n_734),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_730),
.A2(n_678),
.B(n_676),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_782),
.B(n_657),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_857),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_765),
.B(n_659),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_785),
.B(n_659),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_785),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_828),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_796),
.B(n_676),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_828),
.B(n_333),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_874),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_796),
.B(n_336),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_765),
.B(n_343),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_830),
.B(n_341),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_810),
.B(n_343),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_732),
.B(n_882),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_810),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_752),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_811),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_830),
.A2(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_824),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_833),
.A2(n_378),
.B1(n_355),
.B2(n_357),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_824),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_821),
.B(n_630),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_825),
.B(n_345),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_825),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_842),
.B(n_345),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_833),
.B(n_630),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_842),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_851),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_851),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_734),
.A2(n_522),
.B(n_355),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_858),
.A2(n_364),
.B1(n_295),
.B2(n_301),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_858),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_869),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_719),
.B(n_308),
.C(n_335),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_869),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_827),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_752),
.B(n_349),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_840),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_831),
.B(n_357),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_798),
.A2(n_368),
.B1(n_376),
.B2(n_378),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_841),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_821),
.B(n_368),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_847),
.B(n_376),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_725),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_856),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_768),
.B(n_566),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_731),
.A2(n_380),
.B(n_326),
.Y(n_1058)
);

NOR2xp67_ASAP7_75t_L g1059 ( 
.A(n_807),
.B(n_566),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_829),
.B(n_377),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_865),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_866),
.B(n_876),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_861),
.A2(n_522),
.B(n_495),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_834),
.B(n_522),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_836),
.B(n_522),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_798),
.B(n_0),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_878),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_847),
.B(n_232),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_799),
.B(n_233),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_768),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_845),
.A2(n_689),
.B1(n_622),
.B2(n_576),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_884),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_896),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_898),
.A2(n_731),
.B(n_799),
.C(n_809),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_898),
.B(n_809),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_892),
.B(n_880),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_892),
.B(n_881),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_894),
.B(n_883),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_930),
.A2(n_813),
.B1(n_817),
.B2(n_862),
.Y(n_1079)
);

CKINVDCx10_ASAP7_75t_R g1080 ( 
.A(n_913),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_941),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_899),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_886),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_887),
.A2(n_739),
.B(n_759),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1001),
.A2(n_813),
.B1(n_817),
.B2(n_853),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_960),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_900),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1055),
.A2(n_863),
.B1(n_837),
.B2(n_879),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1008),
.B(n_778),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1055),
.A2(n_769),
.B1(n_770),
.B2(n_778),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_891),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_902),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_905),
.A2(n_759),
.B(n_743),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_933),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_909),
.A2(n_743),
.B(n_769),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_944),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_901),
.B(n_770),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_1066),
.A2(n_339),
.B(n_305),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_890),
.A2(n_338),
.B1(n_292),
.B2(n_285),
.C(n_283),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_902),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_982),
.A2(n_306),
.B(n_234),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_966),
.B(n_0),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_954),
.B(n_228),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1028),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_SL g1105 ( 
.A(n_949),
.B(n_266),
.C(n_265),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1066),
.A2(n_518),
.B(n_527),
.C(n_12),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_966),
.B(n_929),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_949),
.B(n_924),
.C(n_1019),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_910),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_986),
.A2(n_311),
.B(n_237),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_987),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_929),
.B(n_4),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_1009),
.B(n_566),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1050),
.B(n_7),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_954),
.B(n_228),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_916),
.A2(n_319),
.B1(n_249),
.B2(n_254),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_906),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_916),
.B(n_242),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1013),
.B(n_256),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_919),
.B(n_12),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_R g1121 ( 
.A(n_927),
.B(n_260),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1055),
.A2(n_274),
.B1(n_272),
.B2(n_261),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_996),
.B(n_277),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_967),
.A2(n_329),
.B(n_294),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_967),
.A2(n_331),
.B(n_300),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_911),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1055),
.A2(n_282),
.B1(n_340),
.B2(n_307),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_935),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1061),
.B(n_314),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_972),
.A2(n_324),
.B(n_328),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_912),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1025),
.A2(n_527),
.B(n_518),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_919),
.B(n_976),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_1019),
.A2(n_322),
.B(n_332),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_L g1135 ( 
.A1(n_932),
.A2(n_518),
.B(n_527),
.C(n_17),
.Y(n_1135)
);

BUFx4_ASAP7_75t_SL g1136 ( 
.A(n_883),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_902),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_972),
.A2(n_689),
.B(n_622),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_889),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1023),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1045),
.A2(n_689),
.B1(n_622),
.B2(n_576),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_928),
.A2(n_689),
.B(n_622),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1067),
.B(n_13),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_945),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_963),
.A2(n_689),
.B(n_622),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1023),
.A2(n_290),
.B(n_566),
.C(n_576),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1017),
.B(n_985),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_981),
.A2(n_16),
.B(n_22),
.C(n_24),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_931),
.A2(n_290),
.B1(n_25),
.B2(n_26),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_970),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_965),
.A2(n_576),
.B(n_290),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_946),
.B(n_576),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_997),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1045),
.A2(n_1062),
.B(n_1027),
.C(n_932),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_968),
.A2(n_290),
.B(n_491),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_936),
.B(n_22),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_950),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_998),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_960),
.A2(n_921),
.B1(n_1020),
.B2(n_1022),
.Y(n_1159)
);

CKINVDCx11_ASAP7_75t_R g1160 ( 
.A(n_907),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_904),
.A2(n_491),
.B(n_27),
.C(n_28),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1004),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_940),
.B(n_26),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_946),
.B(n_1070),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_897),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_888),
.A2(n_491),
.B(n_66),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_908),
.A2(n_491),
.B(n_72),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_951),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_958),
.A2(n_491),
.B(n_65),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_952),
.B(n_31),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_897),
.B(n_1005),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_973),
.B(n_36),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1052),
.B(n_36),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1070),
.B(n_491),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1070),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1037),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_914),
.A2(n_81),
.B(n_175),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_920),
.A2(n_79),
.B(n_170),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1022),
.A2(n_37),
.B(n_38),
.C(n_42),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1026),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_975),
.B(n_43),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_981),
.A2(n_88),
.B(n_156),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_921),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_978),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_902),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1043),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_979),
.B(n_52),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_980),
.B(n_52),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1070),
.B(n_53),
.Y(n_1189)
);

BUFx8_ASAP7_75t_L g1190 ( 
.A(n_1028),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_983),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1044),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_999),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1010),
.A2(n_113),
.B(n_151),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1037),
.A2(n_54),
.B(n_55),
.C(n_57),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1049),
.B(n_520),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_954),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1021),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1056),
.B(n_520),
.Y(n_1199)
);

NOR3xp33_ASAP7_75t_L g1200 ( 
.A(n_1053),
.B(n_520),
.C(n_90),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1009),
.B(n_520),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1046),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_999),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1038),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_990),
.A2(n_86),
.B(n_111),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_989),
.B(n_971),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_991),
.B(n_520),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_1028),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_SL g1209 ( 
.A(n_1028),
.B(n_520),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_992),
.B(n_126),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_995),
.A2(n_135),
.B1(n_136),
.B2(n_1002),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_990),
.A2(n_934),
.B(n_1025),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_988),
.A2(n_947),
.B(n_915),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1006),
.B(n_1042),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1003),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_915),
.A2(n_947),
.B(n_977),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1042),
.B(n_1029),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_943),
.A2(n_903),
.B(n_925),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1011),
.A2(n_1063),
.B(n_922),
.Y(n_1219)
);

NOR3xp33_ASAP7_75t_SL g1220 ( 
.A(n_1069),
.B(n_1053),
.C(n_1054),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1031),
.B(n_1051),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1047),
.B(n_1000),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1016),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_937),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1047),
.B(n_893),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_994),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_938),
.B(n_942),
.Y(n_1227)
);

CKINVDCx6p67_ASAP7_75t_R g1228 ( 
.A(n_994),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_923),
.A2(n_957),
.B1(n_926),
.B2(n_917),
.Y(n_1229)
);

AND3x2_ASAP7_75t_L g1230 ( 
.A(n_974),
.B(n_1068),
.C(n_923),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1228),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1075),
.B(n_989),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1133),
.A2(n_962),
.B(n_1007),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1197),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1072),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1213),
.A2(n_1065),
.B(n_1064),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1218),
.A2(n_962),
.B(n_1007),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1217),
.A2(n_893),
.B1(n_956),
.B2(n_1048),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1184),
.A2(n_948),
.B(n_1071),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1088),
.A2(n_1058),
.A3(n_1039),
.B(n_953),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1135),
.A2(n_1014),
.B(n_1065),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1183),
.B(n_895),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1083),
.B(n_1035),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1222),
.B(n_1035),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1108),
.B(n_956),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1132),
.A2(n_1064),
.B(n_1014),
.Y(n_1246)
);

AO32x2_ASAP7_75t_L g1247 ( 
.A1(n_1085),
.A2(n_1033),
.A3(n_918),
.B1(n_1060),
.B2(n_959),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1208),
.B(n_1040),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1221),
.A2(n_1036),
.B1(n_1034),
.B2(n_1024),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1112),
.A2(n_1059),
.B(n_885),
.C(n_969),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1219),
.A2(n_1007),
.B(n_885),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1089),
.B(n_1040),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1219),
.A2(n_1012),
.B(n_1018),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1076),
.A2(n_969),
.B(n_1060),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1171),
.B(n_1032),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1212),
.A2(n_1033),
.B(n_1015),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1077),
.A2(n_1033),
.B(n_964),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1091),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1088),
.A2(n_993),
.A3(n_1041),
.B(n_918),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1114),
.B(n_1111),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1085),
.A2(n_1032),
.B1(n_1030),
.B2(n_939),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1093),
.A2(n_955),
.B(n_1030),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1074),
.A2(n_959),
.B(n_961),
.Y(n_1263)
);

O2A1O1Ixp5_ASAP7_75t_L g1264 ( 
.A1(n_1120),
.A2(n_1079),
.B(n_1167),
.C(n_1166),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1073),
.Y(n_1265)
);

AOI211x1_ASAP7_75t_L g1266 ( 
.A1(n_1184),
.A2(n_895),
.B(n_984),
.C(n_1071),
.Y(n_1266)
);

INVx5_ASAP7_75t_L g1267 ( 
.A(n_1103),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1081),
.B(n_895),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1109),
.Y(n_1269)
);

BUFx2_ASAP7_75t_R g1270 ( 
.A(n_1139),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1160),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1084),
.A2(n_1057),
.B(n_1095),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_SL g1273 ( 
.A1(n_1176),
.A2(n_1057),
.B(n_1195),
.C(n_1161),
.Y(n_1273)
);

O2A1O1Ixp5_ASAP7_75t_SL g1274 ( 
.A1(n_1149),
.A2(n_1174),
.B(n_1193),
.C(n_1079),
.Y(n_1274)
);

NOR4xp25_ASAP7_75t_L g1275 ( 
.A(n_1140),
.B(n_1191),
.C(n_1149),
.D(n_1179),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_SL g1276 ( 
.A(n_1197),
.B(n_1208),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_SL g1277 ( 
.A(n_1121),
.B(n_1134),
.C(n_1099),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1126),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1154),
.A2(n_1169),
.B(n_1216),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1155),
.A2(n_1090),
.A3(n_1225),
.B(n_1151),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1164),
.B(n_1086),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1194),
.A2(n_1210),
.B(n_1211),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1204),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_SL g1284 ( 
.A(n_1098),
.B(n_1123),
.C(n_1105),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1196),
.A2(n_1199),
.B(n_1182),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1196),
.A2(n_1199),
.B(n_1177),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1090),
.A2(n_1211),
.A3(n_1146),
.B(n_1173),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1178),
.A2(n_1229),
.B(n_1173),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1082),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1220),
.A2(n_1215),
.B(n_1223),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1205),
.A2(n_1206),
.B(n_1207),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1096),
.B(n_1119),
.Y(n_1292)
);

AND2x6_ASAP7_75t_SL g1293 ( 
.A(n_1189),
.B(n_1129),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1102),
.B(n_1163),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1224),
.B(n_1198),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1106),
.A2(n_1191),
.B(n_1172),
.C(n_1181),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1087),
.B(n_1168),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1203),
.A2(n_1187),
.B1(n_1170),
.B2(n_1156),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1117),
.B(n_1131),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1128),
.A2(n_1153),
.A3(n_1202),
.B(n_1192),
.Y(n_1300)
);

NOR2xp67_ASAP7_75t_L g1301 ( 
.A(n_1208),
.B(n_1226),
.Y(n_1301)
);

AOI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1157),
.A2(n_1143),
.B1(n_1188),
.B2(n_1127),
.C(n_1122),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1113),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1145),
.A2(n_1138),
.B(n_1142),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1097),
.A2(n_1200),
.B(n_1130),
.Y(n_1305)
);

AND3x4_ASAP7_75t_L g1306 ( 
.A(n_1078),
.B(n_1080),
.C(n_1136),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1159),
.B(n_1147),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1092),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1214),
.B(n_1165),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1175),
.B(n_1208),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1144),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1113),
.A2(n_1127),
.B(n_1122),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_1227),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1124),
.A2(n_1125),
.B(n_1201),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1148),
.B(n_1116),
.C(n_1227),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1190),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1150),
.B(n_1162),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1092),
.Y(n_1318)
);

NAND2xp33_ASAP7_75t_R g1319 ( 
.A(n_1230),
.B(n_1103),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1141),
.A2(n_1227),
.B(n_1226),
.Y(n_1320)
);

O2A1O1Ixp5_ASAP7_75t_L g1321 ( 
.A1(n_1118),
.A2(n_1104),
.B(n_1152),
.C(n_1158),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1092),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1104),
.A2(n_1186),
.B(n_1180),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1115),
.A2(n_1100),
.B(n_1137),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1115),
.A2(n_1100),
.B(n_1137),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1190),
.Y(n_1326)
);

AOI221x1_ASAP7_75t_L g1327 ( 
.A1(n_1185),
.A2(n_1045),
.B1(n_898),
.B2(n_1085),
.C(n_1149),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1209),
.B(n_728),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1107),
.B(n_898),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1085),
.A2(n_898),
.B(n_715),
.Y(n_1330)
);

AO32x2_ASAP7_75t_L g1331 ( 
.A1(n_1085),
.A2(n_1149),
.A3(n_1079),
.B1(n_1191),
.B2(n_1184),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1132),
.A2(n_1213),
.B(n_1218),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1107),
.B(n_898),
.Y(n_1333)
);

NOR2x1_ASAP7_75t_SL g1334 ( 
.A(n_1103),
.B(n_1115),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1107),
.B(n_898),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1213),
.A2(n_1132),
.B(n_1219),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_SL g1337 ( 
.A(n_1081),
.Y(n_1337)
);

INVx3_ASAP7_75t_SL g1338 ( 
.A(n_1094),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1108),
.B(n_728),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1081),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1075),
.A2(n_1135),
.B(n_1133),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1111),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1075),
.B(n_715),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1108),
.B(n_728),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1107),
.B(n_898),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1111),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1072),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_SL g1348 ( 
.A1(n_1112),
.A2(n_1074),
.B(n_1120),
.C(n_1133),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1219),
.A2(n_1213),
.B(n_1135),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1088),
.A2(n_1058),
.A3(n_1154),
.B(n_1218),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1136),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1075),
.B(n_898),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1107),
.B(n_898),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1213),
.A2(n_1132),
.B(n_1219),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1107),
.B(n_898),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1133),
.A2(n_1218),
.B(n_887),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1133),
.A2(n_1218),
.B(n_887),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1075),
.B(n_715),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1107),
.B(n_898),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1160),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1107),
.B(n_898),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1075),
.B(n_715),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1072),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1107),
.B(n_898),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1213),
.A2(n_1132),
.B(n_1219),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1107),
.B(n_898),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1213),
.A2(n_1132),
.B(n_1219),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1075),
.B(n_898),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1213),
.A2(n_1132),
.B(n_1219),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1094),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1075),
.B(n_715),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1133),
.A2(n_1218),
.B(n_887),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1075),
.A2(n_898),
.B(n_715),
.C(n_1001),
.Y(n_1373)
);

AO31x2_ASAP7_75t_L g1374 ( 
.A1(n_1088),
.A2(n_1058),
.A3(n_1154),
.B(n_1218),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1111),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1083),
.B(n_886),
.Y(n_1376)
);

AOI221x1_ASAP7_75t_L g1377 ( 
.A1(n_1085),
.A2(n_1045),
.B1(n_898),
.B2(n_1149),
.C(n_1176),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1197),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1091),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1075),
.B(n_715),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1219),
.A2(n_1213),
.B(n_1135),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1075),
.A2(n_898),
.B(n_715),
.C(n_1001),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1111),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1072),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1213),
.A2(n_1132),
.B(n_1219),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1072),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1133),
.A2(n_1218),
.B(n_887),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1088),
.A2(n_1058),
.A3(n_1154),
.B(n_1218),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1365),
.A2(n_1369),
.B(n_1367),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1282),
.A2(n_1279),
.B(n_1356),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1297),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1385),
.A2(n_1304),
.B(n_1256),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1272),
.A2(n_1286),
.B(n_1285),
.Y(n_1394)
);

BUFx2_ASAP7_75t_SL g1395 ( 
.A(n_1360),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1237),
.A2(n_1236),
.B(n_1251),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1373),
.A2(n_1382),
.B(n_1330),
.C(n_1371),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1299),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1290),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1246),
.A2(n_1262),
.B(n_1253),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1309),
.B(n_1294),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1377),
.A2(n_1330),
.B1(n_1327),
.B2(n_1343),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1288),
.A2(n_1372),
.B(n_1357),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1300),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1264),
.A2(n_1291),
.B(n_1257),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1358),
.A2(n_1362),
.B(n_1380),
.C(n_1296),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1300),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1387),
.A2(n_1241),
.B(n_1233),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1245),
.A2(n_1298),
.B1(n_1312),
.B2(n_1359),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1241),
.A2(n_1263),
.B(n_1381),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1349),
.A2(n_1381),
.B(n_1323),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1349),
.A2(n_1303),
.B(n_1274),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1352),
.A2(n_1368),
.B1(n_1366),
.B2(n_1364),
.Y(n_1413)
);

AOI21xp33_ASAP7_75t_L g1414 ( 
.A1(n_1298),
.A2(n_1249),
.B(n_1302),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1348),
.A2(n_1250),
.B(n_1239),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1320),
.A2(n_1254),
.B(n_1314),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1239),
.A2(n_1341),
.B(n_1273),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1277),
.A2(n_1238),
.B1(n_1345),
.B2(n_1361),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1341),
.A2(n_1334),
.B(n_1305),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1271),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1335),
.A2(n_1353),
.B1(n_1355),
.B2(n_1339),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1320),
.A2(n_1314),
.B(n_1305),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1300),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1261),
.A2(n_1238),
.B(n_1249),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1275),
.B(n_1315),
.C(n_1344),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1338),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_SL g1427 ( 
.A1(n_1252),
.A2(n_1324),
.B(n_1325),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1261),
.A2(n_1315),
.B(n_1244),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1275),
.A2(n_1321),
.B(n_1232),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_SL g1430 ( 
.A1(n_1255),
.A2(n_1307),
.B(n_1363),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1370),
.B(n_1316),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1235),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1293),
.B(n_1328),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1342),
.A2(n_1375),
.B1(n_1383),
.B2(n_1346),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1265),
.B(n_1386),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1289),
.A2(n_1384),
.B(n_1347),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1331),
.A2(n_1267),
.B1(n_1295),
.B2(n_1319),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1317),
.A2(n_1311),
.B(n_1247),
.Y(n_1438)
);

INVx3_ASAP7_75t_SL g1439 ( 
.A(n_1351),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1284),
.A2(n_1292),
.B(n_1260),
.C(n_1243),
.Y(n_1440)
);

NAND2x1p5_ASAP7_75t_L g1441 ( 
.A(n_1276),
.B(n_1310),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1268),
.B(n_1242),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1313),
.A2(n_1301),
.B(n_1234),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1331),
.A2(n_1370),
.B(n_1293),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1301),
.A2(n_1378),
.B(n_1234),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1231),
.Y(n_1446)
);

AOI221x1_ASAP7_75t_L g1447 ( 
.A1(n_1281),
.A2(n_1331),
.B1(n_1379),
.B2(n_1278),
.C(n_1269),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1266),
.B(n_1281),
.C(n_1322),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1337),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1248),
.A2(n_1247),
.B(n_1287),
.Y(n_1450)
);

OAI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1326),
.A2(n_1340),
.B1(n_1283),
.B2(n_1316),
.C(n_1376),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1280),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1248),
.A2(n_1287),
.B(n_1318),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1378),
.A2(n_1280),
.B(n_1350),
.Y(n_1454)
);

INVx3_ASAP7_75t_SL g1455 ( 
.A(n_1231),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1280),
.A2(n_1388),
.B(n_1374),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1231),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1350),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1270),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1310),
.B(n_1308),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1350),
.A2(n_1388),
.B(n_1374),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1318),
.B(n_1266),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1287),
.A2(n_1374),
.B(n_1388),
.C(n_1240),
.Y(n_1463)
);

BUFx4f_ASAP7_75t_SL g1464 ( 
.A(n_1318),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1306),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1259),
.B(n_1329),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1259),
.A2(n_890),
.B1(n_715),
.B2(n_924),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1336),
.A2(n_1365),
.B(n_1354),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1300),
.Y(n_1469)
);

AOI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1343),
.A2(n_1358),
.B1(n_1380),
.B2(n_1371),
.C(n_1362),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1350),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1231),
.Y(n_1472)
);

AOI21xp33_ASAP7_75t_L g1473 ( 
.A1(n_1296),
.A2(n_715),
.B(n_898),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1343),
.A2(n_1362),
.B(n_1358),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1258),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1297),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1282),
.A2(n_1279),
.B(n_1356),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1260),
.B(n_1343),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1343),
.A2(n_890),
.B1(n_1362),
.B2(n_1358),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_SL g1481 ( 
.A(n_1316),
.B(n_818),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1343),
.A2(n_1362),
.B(n_1358),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1343),
.A2(n_1362),
.B1(n_1371),
.B2(n_1358),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1343),
.B(n_1358),
.Y(n_1485)
);

NOR2x1_ASAP7_75t_L g1486 ( 
.A(n_1284),
.B(n_1277),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1490)
);

AO31x2_ASAP7_75t_L g1491 ( 
.A1(n_1327),
.A2(n_1377),
.A3(n_1288),
.B(n_1282),
.Y(n_1491)
);

BUFx8_ASAP7_75t_SL g1492 ( 
.A(n_1360),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1493)
);

BUFx12f_ASAP7_75t_L g1494 ( 
.A(n_1271),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_SL g1495 ( 
.A(n_1270),
.B(n_852),
.Y(n_1495)
);

OAI211xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1343),
.A2(n_1362),
.B(n_1371),
.C(n_1358),
.Y(n_1496)
);

AO31x2_ASAP7_75t_L g1497 ( 
.A1(n_1327),
.A2(n_1377),
.A3(n_1288),
.B(n_1282),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1332),
.A2(n_1354),
.B(n_1336),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1313),
.B(n_1320),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1343),
.A2(n_1362),
.B1(n_1371),
.B2(n_1358),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1336),
.A2(n_1365),
.B(n_1354),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1350),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1297),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1271),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1282),
.A2(n_1279),
.B(n_1356),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1349),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1336),
.A2(n_1365),
.B(n_1354),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1260),
.B(n_1343),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1268),
.B(n_1242),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1268),
.B(n_1242),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_SL g1513 ( 
.A(n_1267),
.B(n_1103),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1514)
);

CKINVDCx14_ASAP7_75t_R g1515 ( 
.A(n_1506),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1412),
.A2(n_1456),
.B(n_1463),
.Y(n_1516)
);

CKINVDCx16_ASAP7_75t_R g1517 ( 
.A(n_1506),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1433),
.B(n_1409),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1466),
.B(n_1418),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1401),
.B(n_1435),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1433),
.B(n_1409),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1479),
.A2(n_1406),
.B1(n_1470),
.B2(n_1485),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1463),
.A2(n_1477),
.B(n_1391),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1434),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1418),
.B(n_1470),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1474),
.B(n_1482),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_1485),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1507),
.A2(n_1447),
.B(n_1461),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1392),
.B(n_1398),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1484),
.A2(n_1501),
.B(n_1473),
.C(n_1496),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1397),
.A2(n_1402),
.B(n_1417),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1440),
.A2(n_1513),
.B(n_1402),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1432),
.B(n_1436),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1405),
.A2(n_1393),
.B(n_1399),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1500),
.B(n_1442),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1421),
.B(n_1476),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

O2A1O1Ixp5_ASAP7_75t_L g1538 ( 
.A1(n_1414),
.A2(n_1417),
.B(n_1415),
.C(n_1429),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1496),
.A2(n_1413),
.B(n_1444),
.C(n_1425),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1421),
.B(n_1504),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1475),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1437),
.B(n_1424),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1438),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1438),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1443),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1489),
.A2(n_1505),
.B(n_1499),
.C(n_1451),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1419),
.A2(n_1430),
.B(n_1437),
.C(n_1439),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1424),
.B(n_1428),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1467),
.B(n_1455),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1467),
.B(n_1455),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1424),
.B(n_1491),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1448),
.B(n_1422),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1465),
.A2(n_1431),
.B1(n_1457),
.B2(n_1439),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1465),
.A2(n_1457),
.B1(n_1464),
.B2(n_1459),
.Y(n_1554)
);

BUFx2_ASAP7_75t_R g1555 ( 
.A(n_1492),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1464),
.A2(n_1462),
.B1(n_1441),
.B2(n_1446),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1491),
.B(n_1497),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1458),
.B(n_1471),
.Y(n_1558)
);

AOI211xp5_ASAP7_75t_L g1559 ( 
.A1(n_1450),
.A2(n_1399),
.B(n_1481),
.C(n_1495),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1394),
.A2(n_1411),
.B(n_1410),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1491),
.B(n_1497),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1441),
.A2(n_1446),
.B1(n_1450),
.B2(n_1472),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1458),
.A2(n_1503),
.B(n_1471),
.C(n_1427),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1494),
.A2(n_1420),
.B1(n_1395),
.B2(n_1449),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1503),
.A2(n_1416),
.B(n_1453),
.C(n_1408),
.Y(n_1565)
);

NOR2xp67_ASAP7_75t_L g1566 ( 
.A(n_1426),
.B(n_1452),
.Y(n_1566)
);

O2A1O1Ixp5_ASAP7_75t_L g1567 ( 
.A1(n_1403),
.A2(n_1508),
.B(n_1512),
.C(n_1511),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1446),
.A2(n_1460),
.B1(n_1497),
.B2(n_1509),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1445),
.B(n_1454),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1509),
.A2(n_1502),
.B1(n_1468),
.B2(n_1469),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_1404),
.B(n_1469),
.Y(n_1571)
);

AND2x2_ASAP7_75t_SL g1572 ( 
.A(n_1404),
.B(n_1407),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1396),
.B(n_1509),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1502),
.A2(n_1468),
.B1(n_1423),
.B2(n_1400),
.Y(n_1574)
);

AOI221x1_ASAP7_75t_SL g1575 ( 
.A1(n_1468),
.A2(n_1502),
.B1(n_1389),
.B2(n_1480),
.C(n_1483),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1390),
.A2(n_1487),
.B1(n_1488),
.B2(n_1490),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1493),
.B(n_1498),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1464),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1406),
.A2(n_1373),
.B(n_1382),
.C(n_1330),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1492),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1401),
.B(n_1435),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1401),
.B(n_1435),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1414),
.A2(n_1330),
.B1(n_1358),
.B2(n_1362),
.C(n_1343),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1479),
.A2(n_1406),
.B1(n_1470),
.B2(n_1485),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1492),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1412),
.A2(n_1456),
.B(n_1463),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1466),
.B(n_1418),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1466),
.B(n_1418),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1492),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1466),
.B(n_1418),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1479),
.A2(n_1406),
.B1(n_1470),
.B2(n_1485),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1466),
.B(n_1418),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1569),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1533),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1523),
.B(n_1551),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1531),
.A2(n_1570),
.B(n_1561),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1523),
.B(n_1551),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1543),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1544),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1524),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1573),
.B(n_1557),
.Y(n_1606)
);

INVx4_ASAP7_75t_SL g1607 ( 
.A(n_1535),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1528),
.B(n_1516),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1545),
.B(n_1577),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1570),
.A2(n_1576),
.B(n_1574),
.Y(n_1610)
);

AOI221x1_ASAP7_75t_SL g1611 ( 
.A1(n_1522),
.A2(n_1596),
.B1(n_1586),
.B2(n_1527),
.C(n_1525),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1534),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1574),
.A2(n_1542),
.B(n_1565),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1528),
.B(n_1516),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1552),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1589),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1589),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1560),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1522),
.B(n_1586),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1596),
.B(n_1527),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1542),
.A2(n_1593),
.B(n_1597),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1568),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1519),
.A2(n_1590),
.B(n_1593),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1529),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1548),
.B(n_1560),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1529),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1558),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1519),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1575),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1590),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1591),
.B(n_1597),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1514),
.B(n_1582),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1588),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1575),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1576),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1520),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1584),
.A2(n_1525),
.B(n_1579),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1563),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1571),
.A2(n_1532),
.B(n_1518),
.Y(n_1640)
);

AO21x2_ASAP7_75t_L g1641 ( 
.A1(n_1521),
.A2(n_1540),
.B(n_1536),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1584),
.B(n_1530),
.C(n_1539),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1567),
.Y(n_1643)
);

NAND2x1_ASAP7_75t_L g1644 ( 
.A(n_1562),
.B(n_1556),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1566),
.B(n_1556),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1643),
.B(n_1547),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1606),
.B(n_1625),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1631),
.B(n_1628),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1611),
.A2(n_1546),
.B1(n_1538),
.B2(n_1526),
.C(n_1537),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1606),
.B(n_1550),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1606),
.B(n_1549),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1603),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1612),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1600),
.B(n_1572),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1583),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1607),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1644),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1602),
.B(n_1581),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1629),
.A2(n_1562),
.B(n_1541),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1604),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1605),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1602),
.B(n_1559),
.Y(n_1662)
);

OAI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1611),
.A2(n_1638),
.B1(n_1619),
.B2(n_1642),
.C(n_1620),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1644),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1553),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1628),
.B(n_1553),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1598),
.B(n_1554),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1598),
.B(n_1554),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1663),
.A2(n_1638),
.B1(n_1642),
.B2(n_1620),
.C(n_1619),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1656),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_SL g1671 ( 
.A(n_1657),
.B(n_1664),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1663),
.B(n_1629),
.C(n_1634),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1649),
.A2(n_1634),
.B1(n_1630),
.B2(n_1622),
.C(n_1643),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1657),
.B(n_1612),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1652),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1662),
.A2(n_1641),
.B1(n_1640),
.B2(n_1623),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1660),
.Y(n_1678)
);

AOI222xp33_ASAP7_75t_L g1679 ( 
.A1(n_1649),
.A2(n_1631),
.B1(n_1630),
.B2(n_1639),
.C1(n_1622),
.C2(n_1608),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1646),
.A2(n_1515),
.B(n_1636),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1656),
.B(n_1607),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1656),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1639),
.C(n_1636),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1662),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1662),
.B(n_1608),
.C(n_1614),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1623),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1653),
.A2(n_1615),
.B(n_1614),
.C(n_1608),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1657),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1657),
.B(n_1645),
.Y(n_1689)
);

AOI222xp33_ASAP7_75t_L g1690 ( 
.A1(n_1654),
.A2(n_1622),
.B1(n_1614),
.B2(n_1599),
.C1(n_1641),
.C2(n_1616),
.Y(n_1690)
);

OAI31xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1667),
.A2(n_1632),
.A3(n_1635),
.B(n_1633),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1664),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1648),
.B(n_1637),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1665),
.A2(n_1517),
.B(n_1587),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1659),
.A2(n_1641),
.B1(n_1640),
.B2(n_1623),
.Y(n_1695)
);

CKINVDCx6p67_ASAP7_75t_R g1696 ( 
.A(n_1664),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_R g1697 ( 
.A(n_1668),
.B(n_1580),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1659),
.A2(n_1641),
.B1(n_1640),
.B2(n_1623),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1656),
.Y(n_1699)
);

OAI31xp33_ASAP7_75t_L g1700 ( 
.A1(n_1666),
.A2(n_1617),
.A3(n_1616),
.B(n_1637),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1659),
.A2(n_1610),
.B(n_1613),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1659),
.A2(n_1621),
.B1(n_1601),
.B2(n_1624),
.C(n_1626),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1681),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1674),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1684),
.B(n_1648),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1681),
.Y(n_1706)
);

INVx4_ASAP7_75t_SL g1707 ( 
.A(n_1689),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1674),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1676),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1669),
.A2(n_1661),
.B(n_1665),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1683),
.B(n_1655),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1681),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1676),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1701),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1688),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1678),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1683),
.B(n_1658),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1701),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1701),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1688),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1691),
.B(n_1647),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1670),
.B(n_1647),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1678),
.Y(n_1723)
);

INVx4_ASAP7_75t_R g1724 ( 
.A(n_1688),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1671),
.B(n_1681),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1672),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1692),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1702),
.A2(n_1610),
.B(n_1618),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1692),
.Y(n_1729)
);

NOR3xp33_ASAP7_75t_L g1730 ( 
.A(n_1726),
.B(n_1672),
.C(n_1673),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1728),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1725),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1721),
.B(n_1671),
.Y(n_1733)
);

INVx4_ASAP7_75t_L g1734 ( 
.A(n_1725),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1725),
.B(n_1706),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1725),
.B(n_1689),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1728),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_L g1738 ( 
.A(n_1710),
.B(n_1685),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1704),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1726),
.B(n_1679),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1728),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1724),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1705),
.B(n_1685),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1721),
.B(n_1682),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1704),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1710),
.B(n_1700),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1708),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1725),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1728),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1708),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1709),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1721),
.B(n_1706),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1705),
.B(n_1700),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1706),
.B(n_1682),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1709),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_SL g1756 ( 
.A(n_1711),
.B(n_1697),
.C(n_1680),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1728),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1706),
.B(n_1689),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1712),
.B(n_1699),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1711),
.B(n_1693),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1717),
.B(n_1713),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1717),
.B(n_1686),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1715),
.B(n_1555),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1712),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1689),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1703),
.B(n_1696),
.Y(n_1767)
);

NAND4xp25_ASAP7_75t_L g1768 ( 
.A(n_1715),
.B(n_1680),
.C(n_1694),
.D(n_1687),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1703),
.B(n_1722),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1716),
.B(n_1693),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1703),
.B(n_1696),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1739),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1733),
.B(n_1720),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.Y(n_1774)
);

OA21x2_ASAP7_75t_L g1775 ( 
.A1(n_1731),
.A2(n_1741),
.B(n_1737),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1730),
.B(n_1690),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1740),
.B(n_1555),
.Y(n_1777)
);

NOR4xp25_ASAP7_75t_L g1778 ( 
.A(n_1740),
.B(n_1720),
.C(n_1729),
.D(n_1719),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1739),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1730),
.B(n_1650),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1738),
.A2(n_1677),
.B1(n_1694),
.B2(n_1692),
.Y(n_1781)
);

INVxp33_ASAP7_75t_L g1782 ( 
.A(n_1764),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1761),
.B(n_1729),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1733),
.B(n_1727),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1761),
.B(n_1716),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1745),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1738),
.B(n_1650),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1742),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1746),
.B(n_1650),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1746),
.B(n_1753),
.Y(n_1790)
);

NAND2x2_ASAP7_75t_L g1791 ( 
.A(n_1742),
.B(n_1727),
.Y(n_1791)
);

NAND2x1_ASAP7_75t_L g1792 ( 
.A(n_1734),
.B(n_1724),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1735),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1770),
.B(n_1723),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1727),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1748),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1735),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1745),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1752),
.B(n_1722),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1747),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1747),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1756),
.A2(n_1695),
.B(n_1698),
.C(n_1675),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1731),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1753),
.B(n_1651),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1744),
.B(n_1722),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1806)
);

NAND2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1748),
.B(n_1675),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1770),
.B(n_1723),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1788),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1778),
.B(n_1769),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1782),
.B(n_1592),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1790),
.B(n_1769),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1767),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1795),
.B(n_1767),
.Y(n_1814)
);

INVxp67_ASAP7_75t_L g1815 ( 
.A(n_1777),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1796),
.B(n_1762),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1777),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1804),
.B(n_1762),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1776),
.B(n_1744),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1788),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1805),
.B(n_1793),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1773),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1805),
.B(n_1771),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1793),
.B(n_1736),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1781),
.A2(n_1749),
.B1(n_1757),
.B2(n_1737),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1782),
.B(n_1768),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1793),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1802),
.A2(n_1743),
.B1(n_1736),
.B2(n_1734),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1780),
.B(n_1743),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1773),
.B(n_1784),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1785),
.B(n_1763),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1783),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1772),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1819),
.A2(n_1741),
.B1(n_1749),
.B2(n_1757),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1822),
.B(n_1799),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1826),
.A2(n_1741),
.B1(n_1749),
.B2(n_1757),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1810),
.A2(n_1802),
.B(n_1787),
.C(n_1737),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1833),
.B(n_1820),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1827),
.A2(n_1791),
.B1(n_1789),
.B2(n_1797),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_L g1841 ( 
.A(n_1829),
.B(n_1728),
.C(n_1774),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1811),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1809),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1834),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1834),
.Y(n_1845)
);

OAI21xp33_ASAP7_75t_L g1846 ( 
.A1(n_1830),
.A2(n_1784),
.B(n_1768),
.Y(n_1846)
);

XNOR2xp5_ASAP7_75t_L g1847 ( 
.A(n_1831),
.B(n_1825),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_L g1848 ( 
.A(n_1809),
.B(n_1792),
.Y(n_1848)
);

NOR2xp67_ASAP7_75t_L g1849 ( 
.A(n_1828),
.B(n_1797),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1820),
.B(n_1799),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1815),
.A2(n_1791),
.B1(n_1734),
.B2(n_1807),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1828),
.B(n_1735),
.Y(n_1852)
);

OAI21xp33_ASAP7_75t_L g1853 ( 
.A1(n_1817),
.A2(n_1785),
.B(n_1763),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1824),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1839),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1843),
.B(n_1812),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1853),
.B(n_1831),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1847),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1850),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1852),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1836),
.B(n_1821),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1852),
.B(n_1825),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1849),
.B(n_1821),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_SL g1864 ( 
.A(n_1842),
.B(n_1564),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1848),
.B(n_1825),
.Y(n_1865)
);

OAI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1864),
.A2(n_1846),
.B(n_1814),
.Y(n_1866)
);

AOI311xp33_ASAP7_75t_L g1867 ( 
.A1(n_1855),
.A2(n_1840),
.A3(n_1854),
.B(n_1824),
.C(n_1851),
.Y(n_1867)
);

OAI21xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1862),
.A2(n_1823),
.B(n_1734),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1865),
.Y(n_1869)
);

AOI21xp33_ASAP7_75t_L g1870 ( 
.A1(n_1858),
.A2(n_1838),
.B(n_1841),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1863),
.A2(n_1835),
.B(n_1837),
.Y(n_1871)
);

NOR3xp33_ASAP7_75t_L g1872 ( 
.A(n_1859),
.B(n_1816),
.C(n_1844),
.Y(n_1872)
);

AOI222xp33_ASAP7_75t_L g1873 ( 
.A1(n_1857),
.A2(n_1845),
.B1(n_1774),
.B2(n_1803),
.C1(n_1719),
.C2(n_1714),
.Y(n_1873)
);

NAND4xp25_ASAP7_75t_L g1874 ( 
.A(n_1864),
.B(n_1825),
.C(n_1814),
.D(n_1813),
.Y(n_1874)
);

AOI21xp33_ASAP7_75t_L g1875 ( 
.A1(n_1860),
.A2(n_1832),
.B(n_1803),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1870),
.A2(n_1865),
.B1(n_1861),
.B2(n_1775),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1869),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1871),
.A2(n_1856),
.B(n_1832),
.C(n_1818),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1866),
.B(n_1823),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1872),
.B(n_1813),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1873),
.A2(n_1775),
.B1(n_1806),
.B2(n_1818),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_SL g1882 ( 
.A(n_1877),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1880),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1879),
.B(n_1867),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1878),
.B(n_1868),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1876),
.A2(n_1875),
.B(n_1874),
.Y(n_1886)
);

NAND2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1881),
.B(n_1771),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1877),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1886),
.A2(n_1884),
.B(n_1887),
.Y(n_1889)
);

NOR2x1_ASAP7_75t_L g1890 ( 
.A(n_1888),
.B(n_1779),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1883),
.A2(n_1775),
.B1(n_1806),
.B2(n_1801),
.Y(n_1891)
);

NOR3xp33_ASAP7_75t_L g1892 ( 
.A(n_1886),
.B(n_1806),
.C(n_1798),
.Y(n_1892)
);

OAI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1885),
.A2(n_1732),
.B(n_1765),
.C(n_1786),
.Y(n_1893)
);

OAI321xp33_ASAP7_75t_L g1894 ( 
.A1(n_1891),
.A2(n_1882),
.A3(n_1807),
.B1(n_1714),
.B2(n_1718),
.C(n_1719),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1890),
.Y(n_1895)
);

AOI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1889),
.A2(n_1808),
.B(n_1794),
.C(n_1732),
.Y(n_1896)
);

NAND4xp25_ASAP7_75t_L g1897 ( 
.A(n_1895),
.B(n_1892),
.C(n_1893),
.D(n_1732),
.Y(n_1897)
);

AOI322xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1894),
.A3(n_1896),
.B1(n_1719),
.B2(n_1718),
.C1(n_1714),
.C2(n_1732),
.Y(n_1898)
);

AOI222xp33_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1714),
.B1(n_1718),
.B2(n_1760),
.C1(n_1751),
.C2(n_1755),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_SL g1900 ( 
.A1(n_1898),
.A2(n_1751),
.B(n_1750),
.Y(n_1900)
);

OAI22x1_ASAP7_75t_L g1901 ( 
.A1(n_1899),
.A2(n_1735),
.B1(n_1765),
.B2(n_1758),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1900),
.Y(n_1902)
);

OAI22xp5_ASAP7_75t_SL g1903 ( 
.A1(n_1902),
.A2(n_1765),
.B1(n_1578),
.B2(n_1766),
.Y(n_1903)
);

OAI22x1_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1901),
.B1(n_1765),
.B2(n_1766),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1718),
.B(n_1750),
.Y(n_1905)
);

NAND2xp33_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1755),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1760),
.B(n_1758),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1907),
.A2(n_1766),
.B1(n_1758),
.B2(n_1754),
.C(n_1759),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1766),
.B(n_1758),
.C(n_1754),
.Y(n_1909)
);


endmodule