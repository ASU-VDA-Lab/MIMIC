module fake_jpeg_30426_n_510 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_9),
.B(n_3),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_69),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_80),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_28),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_15),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_25),
.Y(n_135)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_33),
.B1(n_31),
.B2(n_34),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_103),
.A2(n_88),
.B1(n_74),
.B2(n_68),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_51),
.B(n_32),
.C(n_42),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_17),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_39),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_96),
.B1(n_94),
.B2(n_65),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_121),
.A2(n_85),
.B1(n_81),
.B2(n_27),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_126),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_42),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_71),
.B(n_51),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_47),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_78),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_101),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_161),
.B(n_163),
.Y(n_237)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_106),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_165),
.B(n_168),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_167),
.B1(n_184),
.B2(n_206),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_93),
.B1(n_61),
.B2(n_67),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_39),
.Y(n_168)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_169),
.Y(n_229)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_170),
.Y(n_241)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_171),
.Y(n_224)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_13),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_66),
.C(n_73),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_177),
.B(n_131),
.Y(n_247)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_17),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_180),
.B(n_181),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_35),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_115),
.A2(n_87),
.B1(n_84),
.B2(n_75),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_182),
.A2(n_185),
.B1(n_213),
.B2(n_100),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_108),
.B(n_35),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_191),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_98),
.B1(n_53),
.B2(n_56),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_113),
.A2(n_62),
.B1(n_99),
.B2(n_97),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_47),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_26),
.Y(n_191)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_192),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_122),
.B(n_26),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_30),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_144),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_197),
.Y(n_257)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

BUFx4f_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_200),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_203),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

CKINVDCx12_ASAP7_75t_R g205 ( 
.A(n_125),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_205),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_136),
.B(n_24),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_210),
.Y(n_234)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_209),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_141),
.B(n_24),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_131),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_110),
.B(n_19),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_110),
.B(n_135),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_158),
.A2(n_37),
.B1(n_31),
.B2(n_33),
.Y(n_213)
);

AOI22x1_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_107),
.B1(n_145),
.B2(n_126),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g270 ( 
.A1(n_215),
.A2(n_245),
.B1(n_127),
.B2(n_137),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_125),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_216),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_220),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_177),
.A2(n_156),
.B(n_109),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_222),
.A2(n_228),
.B(n_239),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_103),
.B1(n_121),
.B2(n_155),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_225),
.B1(n_244),
.B2(n_25),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_37),
.B1(n_34),
.B2(n_138),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_140),
.B(n_129),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_238),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_172),
.A2(n_159),
.B(n_116),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_133),
.B1(n_142),
.B2(n_111),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_178),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_185),
.B(n_20),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_253),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_20),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_246),
.Y(n_328)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_245),
.A2(n_182),
.B1(n_213),
.B2(n_167),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_265),
.A2(n_267),
.B1(n_272),
.B2(n_276),
.Y(n_300)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_184),
.B1(n_174),
.B2(n_192),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_258),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_281),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_195),
.B1(n_204),
.B2(n_203),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_171),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_278),
.Y(n_301)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

BUFx24_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

INVx13_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_215),
.A2(n_198),
.B1(n_202),
.B2(n_186),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_217),
.A2(n_208),
.B1(n_200),
.B2(n_164),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_277),
.A2(n_293),
.B1(n_227),
.B2(n_236),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_223),
.A2(n_176),
.B1(n_151),
.B2(n_208),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_279),
.Y(n_312)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_215),
.A2(n_56),
.B(n_53),
.C(n_179),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_282),
.A2(n_218),
.B(n_233),
.C(n_224),
.Y(n_305)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_283),
.Y(n_317)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_41),
.B(n_40),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_222),
.A2(n_197),
.B(n_196),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_224),
.B(n_253),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_164),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_287),
.B(n_294),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_30),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_289),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_244),
.A2(n_34),
.B1(n_33),
.B2(n_196),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_235),
.B(n_179),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_240),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_252),
.Y(n_334)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_298),
.Y(n_323)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_264),
.A2(n_239),
.B(n_216),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_299),
.A2(n_322),
.B(n_332),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_264),
.A2(n_228),
.B(n_233),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_303),
.B(n_335),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_238),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_320),
.C(n_331),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_270),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_316),
.B(n_325),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_232),
.B(n_257),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_260),
.A2(n_243),
.B(n_237),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_327),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_251),
.C(n_234),
.Y(n_320)
);

AO22x1_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_250),
.B1(n_232),
.B2(n_256),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_234),
.B(n_255),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_246),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_329),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_257),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_257),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_229),
.C(n_241),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_282),
.A2(n_250),
.B(n_1),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_334),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_263),
.B(n_221),
.Y(n_335)
);

INVx4_ASAP7_75t_SL g336 ( 
.A(n_319),
.Y(n_336)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_278),
.B1(n_267),
.B2(n_265),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_338),
.A2(n_357),
.B1(n_305),
.B2(n_250),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_340),
.A2(n_316),
.B(n_332),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_333),
.B(n_325),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_341),
.B(n_364),
.Y(n_371)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_300),
.A2(n_301),
.B1(n_281),
.B2(n_311),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_351),
.B1(n_361),
.B2(n_322),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_344),
.Y(n_377)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

INVx13_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_352),
.Y(n_375)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_329),
.Y(n_350)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_300),
.A2(n_270),
.B1(n_296),
.B2(n_289),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_308),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_307),
.A2(n_270),
.B1(n_271),
.B2(n_290),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_298),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_362),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_301),
.A2(n_271),
.B1(n_261),
.B2(n_262),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_327),
.B(n_297),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_268),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_307),
.A2(n_283),
.B1(n_269),
.B2(n_285),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_266),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_366),
.B(n_367),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_304),
.B(n_292),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_311),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_368),
.B(n_321),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_328),
.C(n_331),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_388),
.C(n_392),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_385),
.B(n_340),
.Y(n_407)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_299),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_371),
.B(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_318),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_343),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_358),
.B(n_303),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_391),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_336),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_384),
.A2(n_338),
.B1(n_337),
.B2(n_350),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_359),
.A2(n_310),
.B(n_322),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_312),
.Y(n_386)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_324),
.C(n_312),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_396),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_305),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_305),
.Y(n_392)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_279),
.C(n_291),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_353),
.C(n_355),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_SL g398 ( 
.A(n_345),
.B(n_315),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_398),
.B(n_345),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_400),
.A2(n_417),
.B1(n_378),
.B2(n_390),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_375),
.B(n_422),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_402),
.B(n_413),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_412),
.C(n_414),
.Y(n_426)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_407),
.A2(n_410),
.B(n_419),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_389),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_408),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_346),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_385),
.A2(n_340),
.B(n_339),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_354),
.C(n_356),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_361),
.C(n_365),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_376),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_394),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_339),
.B1(n_357),
.B2(n_351),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_381),
.B1(n_382),
.B2(n_393),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_373),
.A2(n_359),
.B1(n_344),
.B2(n_293),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_321),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_421),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_370),
.A2(n_347),
.B(n_280),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_372),
.B(n_41),
.C(n_40),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_418),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_219),
.Y(n_421)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_391),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_437),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_407),
.A2(n_373),
.B(n_392),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_432),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_386),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_421),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_434),
.A2(n_439),
.B1(n_419),
.B2(n_410),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_397),
.C(n_396),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_404),
.C(n_400),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_440),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_411),
.A2(n_406),
.B1(n_414),
.B2(n_399),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_378),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_377),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_443),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g443 ( 
.A(n_423),
.B(n_374),
.CI(n_313),
.CON(n_443),
.SN(n_443)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_441),
.B(n_413),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_444),
.A2(n_453),
.B(n_455),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_456),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_452),
.C(n_454),
.Y(n_471)
);

BUFx4f_ASAP7_75t_SL g450 ( 
.A(n_424),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_313),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_411),
.C(n_408),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_433),
.B(n_408),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_420),
.C(n_374),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_426),
.B(n_11),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_439),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_219),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_431),
.B(n_10),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_459),
.A2(n_12),
.B1(n_10),
.B2(n_3),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_431),
.B1(n_428),
.B2(n_432),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_450),
.A2(n_440),
.B1(n_425),
.B2(n_429),
.Y(n_465)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_446),
.A2(n_443),
.B1(n_425),
.B2(n_430),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_443),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_446),
.A2(n_430),
.B1(n_293),
.B2(n_236),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_468),
.B(n_473),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_469),
.B(n_472),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_460),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_454),
.Y(n_476)
);

XOR2x2_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_275),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_475),
.B(n_12),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_477),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_467),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_452),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_482),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_448),
.B(n_450),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_0),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_274),
.C(n_1),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_474),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_487),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_489),
.A2(n_492),
.B(n_493),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_486),
.B(n_463),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_491),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_477),
.B(n_474),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_484),
.A2(n_469),
.B1(n_472),
.B2(n_465),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_479),
.C(n_485),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_495),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_490),
.A2(n_481),
.B(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_498),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_488),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_503),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_479),
.C(n_1),
.Y(n_503)
);

AOI322xp5_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_499),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_505),
.A2(n_0),
.B(n_4),
.Y(n_506)
);

OAI21x1_ASAP7_75t_SL g507 ( 
.A1(n_506),
.A2(n_504),
.B(n_6),
.Y(n_507)
);

AOI21x1_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_5),
.B(n_7),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_5),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_7),
.Y(n_510)
);


endmodule