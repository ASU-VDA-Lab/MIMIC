module fake_jpeg_899_n_685 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_685);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_685;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_61),
.B(n_69),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_64),
.Y(n_212)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_68),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_9),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_86),
.Y(n_133)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_76),
.Y(n_164)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_77),
.Y(n_183)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_79),
.Y(n_225)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_31),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_82),
.B(n_97),
.Y(n_170)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_84),
.Y(n_198)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_98),
.Y(n_157)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_91),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_9),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_100),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_30),
.B(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_106),
.Y(n_172)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_30),
.B(n_7),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_25),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_109),
.B(n_112),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_25),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_25),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_114),
.B(n_116),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_49),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g182 ( 
.A(n_128),
.Y(n_182)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_58),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_130),
.B(n_131),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_58),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_34),
.Y(n_132)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_105),
.B1(n_129),
.B2(n_107),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_81),
.A2(n_56),
.B1(n_29),
.B2(n_34),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_56),
.B1(n_39),
.B2(n_26),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_84),
.A2(n_56),
.B1(n_28),
.B2(n_39),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_145),
.B(n_202),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_28),
.B1(n_52),
.B2(n_32),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_147),
.A2(n_168),
.B1(n_184),
.B2(n_193),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_89),
.A2(n_38),
.B1(n_27),
.B2(n_51),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_150),
.A2(n_64),
.B1(n_127),
.B2(n_113),
.Y(n_239)
);

OR2x4_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_45),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_153),
.A2(n_171),
.B(n_173),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_83),
.A2(n_38),
.B1(n_59),
.B2(n_33),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_158),
.A2(n_169),
.B1(n_175),
.B2(n_176),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_92),
.A2(n_32),
.B1(n_52),
.B2(n_29),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_68),
.A2(n_38),
.B1(n_59),
.B2(n_24),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_76),
.B(n_27),
.Y(n_171)
);

NAND2x1_ASAP7_75t_L g173 ( 
.A(n_93),
.B(n_24),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_71),
.A2(n_24),
.B1(n_60),
.B2(n_43),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_67),
.A2(n_24),
.B1(n_45),
.B2(n_51),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_94),
.A2(n_24),
.B1(n_47),
.B2(n_12),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_77),
.B(n_10),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_187),
.B(n_191),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_79),
.B(n_10),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_78),
.A2(n_124),
.B1(n_126),
.B2(n_95),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_12),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_96),
.A2(n_47),
.B1(n_6),
.B2(n_13),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_205),
.A2(n_206),
.B1(n_213),
.B2(n_217),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_128),
.A2(n_47),
.B1(n_13),
.B2(n_14),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_99),
.A2(n_47),
.B(n_13),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_211),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_100),
.A2(n_115),
.B1(n_120),
.B2(n_118),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_208),
.A2(n_226),
.B1(n_117),
.B2(n_4),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_66),
.B(n_74),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_62),
.A2(n_5),
.B1(n_17),
.B2(n_15),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_72),
.A2(n_5),
.B1(n_17),
.B2(n_15),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_101),
.A2(n_4),
.B1(n_17),
.B2(n_14),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_224),
.A2(n_19),
.B(n_138),
.C(n_226),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_133),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_227),
.B(n_241),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_162),
.B(n_1),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_228),
.B(n_238),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_170),
.A2(n_103),
.B(n_123),
.C(n_64),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_230),
.A2(n_279),
.B(n_176),
.C(n_175),
.Y(n_315)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_233),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_164),
.Y(n_235)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_1),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_239),
.A2(n_251),
.B1(n_275),
.B2(n_218),
.Y(n_308)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_240),
.Y(n_342)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_134),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_242),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_244),
.Y(n_356)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_245),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_185),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_247),
.B(n_256),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_202),
.B(n_70),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_249),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_150),
.A2(n_209),
.B1(n_208),
.B2(n_196),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_252),
.A2(n_277),
.B1(n_304),
.B2(n_307),
.Y(n_350)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_140),
.B(n_3),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_255),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_220),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_143),
.B(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_260),
.Y(n_311)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_149),
.B(n_4),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_197),
.Y(n_262)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_262),
.Y(n_345)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_200),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_265),
.Y(n_316)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_136),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_17),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_267),
.Y(n_321)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_269),
.B(n_271),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_19),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_171),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_272),
.B(n_274),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_165),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_159),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_163),
.B(n_19),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_285),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_215),
.B1(n_167),
.B2(n_195),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_157),
.A2(n_19),
.B(n_173),
.C(n_181),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_188),
.B(n_194),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_281),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_160),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_144),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_161),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_283),
.B(n_288),
.Y(n_347)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_219),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_289),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_224),
.B(n_211),
.Y(n_285)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_286),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_287),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_204),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_155),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_146),
.B(n_167),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_306),
.Y(n_326)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_155),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_291),
.B(n_292),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_201),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_223),
.B(n_195),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_293),
.B(n_296),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_300),
.Y(n_336)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_135),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_141),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_297),
.B(n_299),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_141),
.B(n_222),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_298),
.Y(n_359)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_152),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_152),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_302),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_166),
.B(n_222),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_198),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_303),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_198),
.A2(n_177),
.B1(n_151),
.B2(n_156),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_135),
.B(n_190),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_305),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_166),
.B(n_203),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_151),
.A2(n_156),
.B1(n_177),
.B2(n_193),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_308),
.B(n_231),
.Y(n_390)
);

OAI21x1_ASAP7_75t_SL g375 ( 
.A1(n_315),
.A2(n_276),
.B(n_238),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_169),
.B1(n_205),
.B2(n_214),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_317),
.A2(n_249),
.B1(n_239),
.B2(n_261),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_243),
.B(n_203),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_323),
.B(n_329),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_298),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_257),
.B(n_214),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_338),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_260),
.B(n_190),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_230),
.A2(n_158),
.B(n_213),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_343),
.B(n_367),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_228),
.B(n_190),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_340),
.B(n_244),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_259),
.A2(n_217),
.B(n_206),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_250),
.A2(n_199),
.B1(n_229),
.B2(n_278),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_261),
.B1(n_290),
.B2(n_306),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_229),
.A2(n_199),
.B1(n_270),
.B2(n_268),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_360),
.A2(n_362),
.B1(n_318),
.B2(n_345),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_272),
.A2(n_199),
.B1(n_261),
.B2(n_248),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_298),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_363),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g364 ( 
.A(n_279),
.B(n_235),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_235),
.B(n_273),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_302),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_240),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_275),
.A2(n_261),
.B(n_307),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_370),
.A2(n_384),
.B1(n_387),
.B2(n_404),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_313),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_383),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_372),
.B(n_375),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_237),
.C(n_249),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_397),
.C(n_411),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_232),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_401),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_367),
.A2(n_350),
.B1(n_308),
.B2(n_315),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_380),
.A2(n_386),
.B1(n_393),
.B2(n_415),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_381),
.A2(n_391),
.B(n_402),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_234),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_382),
.A2(n_358),
.B(n_347),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_334),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_326),
.A2(n_304),
.B1(n_302),
.B2(n_301),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

AO21x2_ASAP7_75t_L g386 ( 
.A1(n_350),
.A2(n_297),
.B(n_300),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_325),
.A2(n_303),
.B1(n_233),
.B2(n_236),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_315),
.A2(n_263),
.B(n_282),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_388),
.A2(n_361),
.B(n_347),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_389),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_390),
.A2(n_359),
.B1(n_361),
.B2(n_349),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_339),
.A2(n_284),
.B(n_267),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_351),
.A2(n_289),
.B1(n_253),
.B2(n_291),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

INVx8_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_396),
.Y(n_430)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_320),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_397),
.B(n_399),
.Y(n_429)
);

BUFx24_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_398),
.Y(n_428)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_314),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_400),
.B(n_408),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_311),
.B(n_295),
.Y(n_401)
);

NAND2xp67_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_254),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_325),
.A2(n_246),
.B1(n_262),
.B2(n_269),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_405),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_334),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_406),
.B(n_414),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_317),
.A2(n_242),
.B1(n_265),
.B2(n_245),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_407),
.A2(n_349),
.B1(n_336),
.B2(n_312),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_311),
.B(n_333),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_411),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_320),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_412),
.B(n_413),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_309),
.B(n_240),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_258),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_329),
.A2(n_286),
.B1(n_296),
.B2(n_366),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_416),
.A2(n_352),
.B1(n_312),
.B2(n_345),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_417),
.A2(n_376),
.B(n_381),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_369),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_418),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_419),
.B(n_424),
.C(n_427),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_410),
.B(n_309),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_421),
.B(n_334),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_330),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_330),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_380),
.A2(n_372),
.B1(n_386),
.B2(n_376),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_432),
.A2(n_434),
.B1(n_438),
.B2(n_370),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_386),
.A2(n_343),
.B1(n_363),
.B2(n_359),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_435),
.A2(n_453),
.B(n_454),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_382),
.A2(n_335),
.B1(n_321),
.B2(n_322),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_436),
.A2(n_449),
.B1(n_407),
.B2(n_402),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_386),
.A2(n_323),
.B1(n_338),
.B2(n_335),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_373),
.B(n_341),
.C(n_316),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_442),
.B(n_447),
.C(n_451),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_386),
.A2(n_340),
.B1(n_322),
.B2(n_321),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_444),
.A2(n_382),
.B1(n_406),
.B2(n_390),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_409),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_371),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_316),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_358),
.C(n_310),
.Y(n_451)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_452),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_375),
.B(n_310),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_353),
.C(n_320),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_458),
.B(n_412),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_460),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_424),
.B(n_403),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_419),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_383),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_467),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_464),
.A2(n_485),
.B1(n_490),
.B2(n_492),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_465),
.A2(n_470),
.B1(n_478),
.B2(n_434),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_354),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g528 ( 
.A(n_466),
.Y(n_528)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_388),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_471),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_423),
.A2(n_386),
.B1(n_390),
.B2(n_393),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_430),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_430),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_481),
.Y(n_508)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_458),
.B(n_413),
.Y(n_474)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_474),
.Y(n_514)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_475),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_450),
.A2(n_391),
.B(n_408),
.Y(n_476)
);

OAI21xp33_ASAP7_75t_L g503 ( 
.A1(n_476),
.A2(n_448),
.B(n_454),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_450),
.A2(n_415),
.B1(n_384),
.B2(n_400),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_441),
.Y(n_480)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_480),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_420),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_426),
.B(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_420),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_483),
.B(n_486),
.Y(n_531)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_484),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_354),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_394),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_487),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_456),
.B(n_392),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_455),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_489),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_432),
.A2(n_404),
.B1(n_387),
.B2(n_399),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_422),
.A2(n_377),
.B1(n_349),
.B2(n_416),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_493),
.B(n_497),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_451),
.B(n_348),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_494),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_446),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_453),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_498),
.B(n_482),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_503),
.A2(n_489),
.B(n_484),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_504),
.A2(n_509),
.B1(n_515),
.B2(n_524),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_421),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_507),
.B(n_525),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_464),
.A2(n_422),
.B1(n_450),
.B2(n_423),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_447),
.C(n_442),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_511),
.C(n_516),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_443),
.C(n_429),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_513),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_469),
.A2(n_438),
.B1(n_444),
.B2(n_443),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_429),
.C(n_435),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_469),
.A2(n_457),
.B1(n_449),
.B2(n_433),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_468),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_448),
.C(n_433),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_521),
.C(n_534),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_455),
.C(n_344),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_465),
.A2(n_428),
.B1(n_439),
.B2(n_440),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_461),
.B(n_353),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_491),
.B(n_474),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_476),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_491),
.A2(n_428),
.B(n_439),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_529),
.A2(n_485),
.B(n_488),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_463),
.B(n_344),
.C(n_348),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_528),
.B(n_467),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_537),
.B(n_543),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_501),
.Y(n_538)
);

INVx13_ASAP7_75t_L g580 ( 
.A(n_538),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_518),
.B(n_460),
.Y(n_539)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_539),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_SL g587 ( 
.A(n_540),
.B(n_389),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_542),
.A2(n_563),
.B(n_368),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_512),
.B(n_483),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_507),
.B(n_481),
.C(n_471),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_546),
.C(n_561),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_499),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_545),
.A2(n_559),
.B1(n_560),
.B2(n_562),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_498),
.B(n_472),
.C(n_487),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_526),
.Y(n_547)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_547),
.Y(n_590)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_506),
.Y(n_548)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_548),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_508),
.Y(n_550)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_550),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_551),
.A2(n_524),
.B(n_505),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_510),
.Y(n_573)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_553),
.Y(n_568)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_533),
.Y(n_555)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_555),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_509),
.A2(n_492),
.B1(n_490),
.B2(n_462),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_556),
.A2(n_558),
.B1(n_567),
.B2(n_437),
.Y(n_588)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_519),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_517),
.A2(n_462),
.B1(n_470),
.B2(n_505),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_511),
.B(n_475),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_478),
.C(n_480),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_522),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_530),
.B(n_479),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_564),
.B(n_565),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_534),
.B(n_473),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_525),
.B(n_531),
.Y(n_566)
);

OAI322xp33_ASAP7_75t_L g592 ( 
.A1(n_566),
.A2(n_336),
.A3(n_437),
.B1(n_398),
.B2(n_332),
.C1(n_355),
.C2(n_357),
.Y(n_592)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

O2A1O1Ixp5_ASAP7_75t_L g569 ( 
.A1(n_546),
.A2(n_520),
.B(n_521),
.C(n_513),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_569),
.B(n_540),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_551),
.A2(n_529),
.B(n_503),
.Y(n_571)
);

XNOR2x1_ASAP7_75t_L g595 ( 
.A(n_571),
.B(n_584),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_573),
.B(n_574),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_535),
.B(n_527),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_542),
.A2(n_504),
.B1(n_515),
.B2(n_539),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_576),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_536),
.B(n_500),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_578),
.B(n_587),
.Y(n_603)
);

XOR2x2_ASAP7_75t_L g611 ( 
.A(n_581),
.B(n_589),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_535),
.B(n_500),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_591),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_561),
.C(n_544),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_592),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_563),
.A2(n_532),
.B(n_440),
.Y(n_584)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_588),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_541),
.B(n_336),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_584),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_596),
.B(n_604),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_585),
.A2(n_538),
.B1(n_564),
.B2(n_549),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_597),
.A2(n_606),
.B1(n_567),
.B2(n_558),
.Y(n_633)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_594),
.Y(n_598)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_598),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_570),
.C(n_573),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_594),
.A2(n_550),
.B1(n_548),
.B2(n_555),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_605),
.A2(n_579),
.B1(n_593),
.B2(n_590),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_589),
.A2(n_549),
.B1(n_557),
.B2(n_547),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_575),
.Y(n_607)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_607),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_578),
.B(n_536),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_609),
.B(n_610),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_552),
.Y(n_610)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_575),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_615),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_572),
.B(n_565),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_613),
.Y(n_636)
);

XOR2x2_ASAP7_75t_L g634 ( 
.A(n_614),
.B(n_591),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_574),
.B(n_556),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_579),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_553),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_572),
.B(n_554),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_617),
.Y(n_626)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_618),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_610),
.C(n_599),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_619),
.B(n_620),
.Y(n_638)
);

BUFx24_ASAP7_75t_SL g620 ( 
.A(n_601),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_606),
.A2(n_571),
.B(n_581),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_621),
.A2(n_623),
.B(n_629),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_615),
.C(n_602),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_622),
.B(n_631),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_611),
.A2(n_577),
.B(n_576),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_608),
.A2(n_568),
.B1(n_580),
.B2(n_587),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_627),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_611),
.A2(n_580),
.B(n_568),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_633),
.A2(n_595),
.B1(n_614),
.B2(n_603),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_634),
.A2(n_635),
.B(n_603),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_595),
.A2(n_600),
.B(n_597),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_624),
.B(n_622),
.Y(n_640)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_640),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_643),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_642),
.A2(n_644),
.B(n_650),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_619),
.B(n_586),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_629),
.A2(n_582),
.B(n_602),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_621),
.B(n_609),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_645),
.B(n_646),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_635),
.A2(n_395),
.B(n_389),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_374),
.C(n_324),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_647),
.B(n_649),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_623),
.A2(n_374),
.B1(n_405),
.B2(n_318),
.Y(n_649)
);

INVxp33_ASAP7_75t_SL g650 ( 
.A(n_633),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_356),
.C(n_357),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_652),
.B(n_628),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_640),
.B(n_636),
.Y(n_653)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_653),
.Y(n_665)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_654),
.Y(n_667)
);

AOI211xp5_ASAP7_75t_L g656 ( 
.A1(n_637),
.A2(n_627),
.B(n_625),
.C(n_630),
.Y(n_656)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_656),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_648),
.Y(n_657)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_657),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_638),
.A2(n_625),
.B(n_628),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_658),
.A2(n_660),
.B(n_663),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_651),
.B(n_626),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_634),
.C(n_630),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_655),
.A2(n_651),
.B(n_639),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g674 ( 
.A(n_669),
.B(n_664),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_662),
.A2(n_659),
.B(n_657),
.Y(n_670)
);

A2O1A1O1Ixp25_ASAP7_75t_L g676 ( 
.A1(n_670),
.A2(n_673),
.B(n_647),
.C(n_652),
.D(n_656),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_661),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_671),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_662),
.A2(n_663),
.B(n_645),
.Y(n_673)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_674),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_676),
.A2(n_678),
.B(n_356),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_667),
.B(n_631),
.C(n_398),
.Y(n_677)
);

MAJx2_ASAP7_75t_L g680 ( 
.A(n_677),
.B(n_332),
.C(n_355),
.Y(n_680)
);

AOI321xp33_ASAP7_75t_L g678 ( 
.A1(n_665),
.A2(n_668),
.A3(n_672),
.B1(n_666),
.B2(n_671),
.C(n_398),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_680),
.B(n_675),
.Y(n_682)
);

BUFx24_ASAP7_75t_SL g684 ( 
.A(n_682),
.Y(n_684)
);

OAI311xp33_ASAP7_75t_L g683 ( 
.A1(n_681),
.A2(n_331),
.A3(n_337),
.B1(n_346),
.C1(n_670),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_SL g685 ( 
.A1(n_684),
.A2(n_683),
.B(n_331),
.C(n_346),
.Y(n_685)
);


endmodule