module real_jpeg_26290_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_1),
.A2(n_32),
.B1(n_71),
.B2(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_2),
.A2(n_38),
.B1(n_55),
.B2(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_38),
.B1(n_71),
.B2(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_2),
.A2(n_26),
.B(n_200),
.C(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_27),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_2),
.A2(n_29),
.B(n_53),
.C(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_2),
.B(n_70),
.C(n_71),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_2),
.B(n_51),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_114),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_2),
.B(n_68),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_9),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

CKINVDCx12_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_5),
.A2(n_34),
.B1(n_50),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_5),
.A2(n_50),
.B1(n_71),
.B2(n_73),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_24),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_129),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_129),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_8),
.A2(n_71),
.B1(n_73),
.B2(n_129),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_326),
.Y(n_16)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_39),
.B1(n_43),
.B2(n_323),
.C(n_325),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_18),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_18),
.B(n_324),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_18),
.B(n_39),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_19),
.A2(n_27),
.B(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_20),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_21),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_24),
.Y(n_128)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_24),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_25),
.A2(n_29),
.B(n_38),
.Y(n_200)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_27),
.B(n_127),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_28),
.A2(n_29),
.B1(n_53),
.B2(n_58),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_36),
.B(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_38),
.A2(n_55),
.B(n_58),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_39),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_39),
.A2(n_94),
.B1(n_103),
.B2(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_42),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_40),
.A2(n_82),
.B(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_312),
.B(n_322),
.Y(n_43)
);

OAI211xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_130),
.B(n_146),
.C(n_311),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_104),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_46),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_46),
.B(n_104),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_46),
.B(n_132),
.Y(n_311)
);

FAx1_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_79),
.CI(n_93),
.CON(n_46),
.SN(n_46)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_47),
.A2(n_48),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_63),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B(n_59),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_51),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_52),
.B(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_52),
.A2(n_60),
.B(n_139),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_77)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_56),
.B(n_242),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_59),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_59),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_60),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_74),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_64),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_67),
.B(n_90),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_66),
.B(n_76),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_75),
.B(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_68),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_71),
.B(n_266),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_75),
.B(n_239),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_76),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_80),
.A2(n_91),
.B1(n_134),
.B2(n_144),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_85),
.C(n_88),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_80),
.B(n_134),
.C(n_145),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_81),
.B(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_82),
.B(n_126),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_87),
.B(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_89),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_88),
.B(n_182),
.C(n_184),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_88),
.A2(n_89),
.B1(n_184),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_89),
.B(n_137),
.C(n_140),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_99),
.B(n_103),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_94),
.A2(n_100),
.B1(n_108),
.B2(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_94),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_94),
.A2(n_108),
.B1(n_224),
.B2(n_282),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B(n_98),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_95),
.B(n_98),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_95),
.B(n_253),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_96),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_102),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_102),
.B(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_110),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_109),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.C(n_124),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_112),
.B(n_119),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_113),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_117),
.A2(n_160),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_117),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_124),
.B1(n_125),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_122),
.B(n_186),
.Y(n_279)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_147),
.C(n_148),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_145),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_138),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_141),
.Y(n_318)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_174),
.B(n_310),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_171),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_150),
.B(n_171),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_151),
.B(n_154),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_156),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_168),
.C(n_169),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_157),
.A2(n_158),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_166),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_162),
.B(n_252),
.Y(n_271)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_168),
.A2(n_169),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_168),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_168),
.A2(n_299),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_168),
.B(n_314),
.C(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_169),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_305),
.B(n_309),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_217),
.B(n_291),
.C(n_304),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_205),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_177),
.B(n_205),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_190),
.B2(n_204),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_188),
.B2(n_189),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_180),
.B(n_189),
.C(n_204),
.Y(n_292)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_183),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_187),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_198),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_192),
.B(n_197),
.C(n_198),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_212),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_207),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_215),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_215),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_216),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_290),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_233),
.B(n_289),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_220),
.B(n_230),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.C(n_226),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_221),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_226),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_224),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_284),
.B(n_288),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_275),
.B(n_283),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_256),
.B(n_274),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_237),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_238),
.A2(n_240),
.B1(n_241),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_250),
.B2(n_255),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_249),
.C(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_263),
.B(n_273),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_269),
.B(n_272),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_276),
.B(n_277),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_301),
.B2(n_302),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_302),
.C(n_303),
.Y(n_306)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_321),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_321),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_320),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_317),
.Y(n_319)
);


endmodule