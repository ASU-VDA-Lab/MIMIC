module real_jpeg_32782_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_0),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_2),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_2),
.B(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

NAND2x1_ASAP7_75t_SL g94 ( 
.A(n_4),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_4),
.B(n_129),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_6),
.B(n_123),
.Y(n_122)
);

NAND2xp67_ASAP7_75t_SL g130 ( 
.A(n_6),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_6),
.B(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_6),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_6),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_7),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_7),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_7),
.B(n_83),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_7),
.B(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_8),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_9),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_9),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_9),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_9),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_9),
.B(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_11),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_12),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_13),
.B(n_83),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_13),
.B(n_117),
.Y(n_116)
);

NAND2x1_ASAP7_75t_L g128 ( 
.A(n_13),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_13),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_14),
.B(n_83),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_14),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_15),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_15),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_15),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_15),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_15),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_15),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_15),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_15),
.B(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_209),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_208),
.Y(n_17)
);

INVxp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_162),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_20),
.B(n_162),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_106),
.C(n_138),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_22),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.Y(n_22)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_23),
.B(n_72),
.C(n_164),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.C(n_55),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_25),
.B(n_36),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_26),
.B(n_31),
.C(n_36),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_29),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_35),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_35),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_40),
.Y(n_312)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_40),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_41),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_235)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_43),
.A2(n_44),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_48),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_49),
.Y(n_231)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.C(n_66),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_57),
.A2(n_66),
.B1(n_67),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_57),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_61),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_62),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_63),
.B(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_70),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_87),
.B2(n_88),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_85),
.B2(n_86),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_84),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_77),
.B(n_84),
.C(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_157),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g286 ( 
.A1(n_82),
.A2(n_84),
.B1(n_158),
.B2(n_159),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_83),
.Y(n_265)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_83),
.Y(n_329)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_100),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_90),
.B(n_94),
.C(n_101),
.Y(n_178)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_92),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_98),
.Y(n_320)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_102),
.B(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_107),
.B(n_138),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_111),
.C(n_126),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_126),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_121),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_140),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_120),
.Y(n_284)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_134),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_203),
.C(n_204),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_141),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_142),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.C(n_156),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_143),
.A2(n_144),
.B1(n_150),
.B2(n_151),
.Y(n_347)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_156),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_188),
.B(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_189),
.B(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_202),
.B1(n_206),
.B2(n_207),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

XOR2x2_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_238),
.B(n_358),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_236),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_211),
.B(n_236),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.C(n_232),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_212),
.B(n_356),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_215),
.B(n_233),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_219),
.C(n_229),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_216),
.B(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_219),
.A2(n_229),
.B1(n_230),
.B2(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_219),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.C(n_227),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_SL g277 ( 
.A(n_220),
.B(n_227),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_SL g276 ( 
.A(n_223),
.B(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_353),
.B(n_357),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_340),
.B(n_352),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_288),
.B(n_339),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_273),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_244),
.B(n_273),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_262),
.C(n_270),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_253),
.C(n_258),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_262),
.A2(n_263),
.B1(n_270),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_267),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_276),
.C(n_278),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_286),
.C(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_304),
.B(n_338),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_301),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_301),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.C(n_297),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_291),
.A2(n_292),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_293),
.A2(n_297),
.B1(n_298),
.B2(n_336),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_293),
.Y(n_336)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_331),
.B(n_337),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_321),
.B(n_330),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_318),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_351),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_351),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_348),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_345),
.C(n_348),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_354),
.B(n_355),
.Y(n_357)
);


endmodule