module fake_jpeg_13376_n_179 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_127;
wire n_76;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_21),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_0),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_1),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_3),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_38),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_7),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_22),
.B(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_92),
.Y(n_105)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_93),
.Y(n_95)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_83),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_63),
.B1(n_71),
.B2(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_103),
.B1(n_107),
.B2(n_66),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_64),
.B1(n_67),
.B2(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_78),
.B1(n_62),
.B2(n_79),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_59),
.B1(n_61),
.B2(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_63),
.B1(n_74),
.B2(n_65),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_55),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_120),
.C(n_125),
.Y(n_128)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_119),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_86),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_68),
.B(n_80),
.C(n_5),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_127),
.B(n_109),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_69),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_132),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_131),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_26),
.B(n_52),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_136),
.B(n_10),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_89),
.B1(n_70),
.B2(n_72),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_67),
.B1(n_72),
.B2(n_70),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_138),
.B1(n_144),
.B2(n_33),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_3),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_23),
.C(n_43),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_139),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_20),
.B1(n_40),
.B2(n_37),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_19),
.C(n_36),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_14),
.B(n_16),
.C(n_25),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_27),
.C(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_138),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_161),
.B1(n_146),
.B2(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_158),
.B1(n_160),
.B2(n_155),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_46),
.B(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_162),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_149),
.B1(n_148),
.B2(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_151),
.C(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_166),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_167),
.B1(n_168),
.B2(n_171),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_167),
.B(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_172),
.B(n_163),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_165),
.B(n_170),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_178),
.Y(n_179)
);


endmodule