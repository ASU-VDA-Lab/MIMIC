module fake_jpeg_62_n_440 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_80),
.Y(n_109)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_30),
.A2(n_14),
.B(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_14),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_26),
.Y(n_60)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_76),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_34),
.A2(n_8),
.B(n_13),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_34),
.B(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_83),
.B(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_53),
.B1(n_57),
.B2(n_47),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_85),
.A2(n_88),
.B1(n_92),
.B2(n_104),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_37),
.C(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_37),
.B1(n_42),
.B2(n_40),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_20),
.B1(n_38),
.B2(n_41),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_94),
.A2(n_95),
.B1(n_113),
.B2(n_114),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_49),
.B1(n_60),
.B2(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_38),
.B1(n_41),
.B2(n_32),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_123),
.B1(n_134),
.B2(n_138),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_20),
.B1(n_46),
.B2(n_38),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_46),
.A2(n_41),
.B1(n_32),
.B2(n_39),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_48),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_115),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_135),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_52),
.A2(n_41),
.B1(n_36),
.B2(n_33),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_65),
.A2(n_33),
.B1(n_24),
.B2(n_43),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_66),
.A2(n_43),
.B1(n_24),
.B2(n_9),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_0),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_72),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_6),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_14),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_98),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_74),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_81),
.B1(n_77),
.B2(n_9),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_4),
.B1(n_9),
.B2(n_5),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_154),
.B1(n_158),
.B2(n_161),
.Y(n_200)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_141),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_142),
.B(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_73),
.B1(n_78),
.B2(n_2),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_4),
.B(n_12),
.C(n_2),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_179),
.B(n_170),
.C(n_163),
.Y(n_201)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_157),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_105),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_162),
.B(n_167),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_0),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_105),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_165),
.A2(n_175),
.B1(n_180),
.B2(n_160),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_84),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_101),
.B(n_3),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_181),
.A3(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_239)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_3),
.B1(n_88),
.B2(n_96),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_101),
.B(n_82),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_184),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_112),
.A2(n_139),
.B(n_124),
.C(n_82),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_108),
.B1(n_131),
.B2(n_106),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_131),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_108),
.B(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_119),
.B(n_122),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_128),
.B(n_132),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_128),
.B(n_133),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_111),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_111),
.B(n_122),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_100),
.B(n_107),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_193),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_100),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_152),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_175),
.B1(n_150),
.B2(n_156),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_195),
.A2(n_197),
.B1(n_227),
.B2(n_222),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_142),
.A2(n_176),
.B1(n_153),
.B2(n_150),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_196),
.A2(n_232),
.B1(n_200),
.B2(n_201),
.Y(n_254)
);

AOI22x1_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_154),
.B1(n_143),
.B2(n_181),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_160),
.A2(n_169),
.B1(n_167),
.B2(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_143),
.C(n_159),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_210),
.B(n_234),
.C(n_240),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_155),
.B(n_190),
.C(n_185),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_230),
.B(n_233),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_183),
.B1(n_191),
.B2(n_157),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_222),
.A2(n_230),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_144),
.A2(n_183),
.B1(n_160),
.B2(n_149),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_228),
.A2(n_229),
.B1(n_198),
.B2(n_218),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_182),
.B(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_164),
.A2(n_174),
.B1(n_189),
.B2(n_145),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_152),
.B(n_164),
.C(n_151),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_172),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_172),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_243),
.B(n_263),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_244),
.B(n_276),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_196),
.A2(n_172),
.B1(n_189),
.B2(n_236),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_250),
.B(n_253),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_246),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_189),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_247),
.B(n_261),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_197),
.A2(n_239),
.B1(n_220),
.B2(n_219),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_254),
.B1(n_256),
.B2(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_241),
.B1(n_217),
.B2(n_216),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_197),
.A2(n_219),
.B(n_210),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_257),
.A2(n_260),
.B(n_273),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_214),
.A2(n_224),
.B1(n_217),
.B2(n_203),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_224),
.A2(n_240),
.B(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_203),
.B(n_202),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_213),
.B1(n_202),
.B2(n_211),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_274),
.B1(n_279),
.B2(n_244),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_212),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_234),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_264),
.A2(n_255),
.B(n_259),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_209),
.B(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_266),
.B(n_282),
.Y(n_293)
);

NAND2x1_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_231),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_250),
.B(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_211),
.B1(n_233),
.B2(n_207),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_264),
.B(n_249),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_238),
.A2(n_218),
.B1(n_206),
.B2(n_205),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_256),
.B1(n_276),
.B2(n_272),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_205),
.A2(n_221),
.B1(n_237),
.B2(n_225),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_204),
.A2(n_228),
.B1(n_200),
.B2(n_148),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_248),
.B1(n_281),
.B2(n_243),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_241),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_285),
.A2(n_307),
.B(n_314),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_251),
.CI(n_258),
.CON(n_286),
.SN(n_286)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_286),
.B(n_296),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_294),
.C(n_313),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_247),
.B1(n_282),
.B2(n_245),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_306),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_261),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_304),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_253),
.B(n_249),
.Y(n_296)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_300),
.A2(n_275),
.B1(n_307),
.B2(n_312),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_263),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_SL g305 ( 
.A(n_267),
.B(n_264),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g332 ( 
.A1(n_305),
.A2(n_296),
.B(n_284),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_266),
.B(n_242),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_309),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_268),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_262),
.B(n_265),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_283),
.B(n_316),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_265),
.A2(n_270),
.B1(n_252),
.B2(n_255),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_275),
.C(n_309),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_287),
.B(n_259),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_288),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_273),
.C(n_246),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_324),
.C(n_342),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_285),
.C(n_284),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_304),
.B(n_271),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_343),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_328),
.A2(n_297),
.B1(n_315),
.B2(n_317),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_329),
.B(n_335),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_306),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_341),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_289),
.A2(n_303),
.B1(n_293),
.B2(n_291),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_311),
.B1(n_299),
.B2(n_286),
.Y(n_351)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_339),
.A2(n_298),
.B(n_288),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_302),
.B(n_313),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_340),
.B(n_302),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_293),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_289),
.C(n_303),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_295),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_346),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_286),
.C(n_292),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_315),
.C(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

XOR2x2_ASAP7_75t_SL g371 ( 
.A(n_347),
.B(n_368),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_355),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_351),
.A2(n_354),
.B1(n_364),
.B2(n_331),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_353),
.A2(n_360),
.B(n_370),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_322),
.A2(n_288),
.B1(n_298),
.B2(n_290),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_292),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_339),
.A2(n_298),
.B1(n_314),
.B2(n_290),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_329),
.B1(n_330),
.B2(n_333),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_318),
.B(n_317),
.Y(n_357)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_319),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_297),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_362),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_324),
.C(n_323),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_324),
.C(n_345),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_331),
.B1(n_336),
.B2(n_328),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_326),
.A2(n_345),
.B(n_342),
.C(n_338),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_341),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_367),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_335),
.A2(n_326),
.B(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_348),
.B(n_320),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_383),
.Y(n_391)
);

OA21x2_ASAP7_75t_SL g398 ( 
.A1(n_374),
.A2(n_347),
.B(n_351),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_381),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_377),
.B(n_384),
.Y(n_405)
);

OAI21x1_ASAP7_75t_SL g400 ( 
.A1(n_379),
.A2(n_390),
.B(n_358),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_340),
.C(n_338),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_388),
.C(n_349),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_350),
.B(n_319),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_364),
.A2(n_327),
.B1(n_333),
.B2(n_325),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_334),
.B1(n_337),
.B2(n_344),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_385),
.A2(n_359),
.B1(n_352),
.B2(n_358),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_350),
.B(n_346),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_365),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_349),
.C(n_363),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_352),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_389),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_354),
.Y(n_390)
);

AO21x1_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_353),
.B(n_370),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_381),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_379),
.A2(n_367),
.B(n_366),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_396),
.A2(n_401),
.B(n_372),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_362),
.C(n_368),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_404),
.C(n_371),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_400),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_399),
.A2(n_384),
.B1(n_390),
.B2(n_385),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_365),
.B(n_377),
.Y(n_401)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_403),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_388),
.C(n_375),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_380),
.Y(n_406)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_401),
.A2(n_390),
.B1(n_389),
.B2(n_378),
.Y(n_410)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_376),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_411),
.A2(n_414),
.B(n_398),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_413),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_391),
.A2(n_371),
.B1(n_386),
.B2(n_393),
.Y(n_417)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_417),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_420),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_SL g420 ( 
.A(n_416),
.B(n_400),
.C(n_405),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_396),
.B(n_407),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_425),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_404),
.C(n_395),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_408),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_427),
.B(n_430),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_422),
.A2(n_407),
.B1(n_416),
.B2(n_410),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_429),
.B(n_394),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_393),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_426),
.B(n_423),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_419),
.C(n_428),
.Y(n_435)
);

AOI321xp33_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_433),
.A3(n_420),
.B1(n_429),
.B2(n_392),
.C(n_412),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_436),
.A2(n_434),
.B(n_414),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_437),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_411),
.B(n_405),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_402),
.Y(n_440)
);


endmodule