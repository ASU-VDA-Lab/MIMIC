module fake_jpeg_10002_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_35),
.Y(n_43)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_21),
.B1(n_34),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_47),
.B1(n_32),
.B2(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_47)
);

AOI222xp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_18),
.B1(n_22),
.B2(n_19),
.C1(n_20),
.C2(n_16),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_24),
.C(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_35),
.B1(n_19),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_40),
.B1(n_39),
.B2(n_20),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_60),
.B1(n_40),
.B2(n_16),
.Y(n_74)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_1),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_6),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_64),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_32),
.B1(n_23),
.B2(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_42),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_16),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_81),
.B1(n_65),
.B2(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_9),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_82),
.Y(n_89)
);

OA22x2_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_33),
.C(n_30),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_95),
.C(n_80),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_79),
.B(n_71),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_93),
.B(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_30),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_64),
.C(n_63),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_8),
.C(n_11),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_12),
.C(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_101),
.Y(n_111)
);

OAI21x1_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_93),
.B(n_86),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_74),
.B1(n_81),
.B2(n_63),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_108),
.B(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_13),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_84),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_94),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_107),
.C(n_17),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_91),
.B(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_110),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_89),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_107),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C(n_3),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_118),
.C(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_14),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_119),
.B1(n_120),
.B2(n_117),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_126),
.A3(n_15),
.B1(n_55),
.B2(n_3),
.C1(n_1),
.C2(n_17),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_122),
.B(n_2),
.C(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_133),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_17),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_17),
.C(n_55),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_137),
.A2(n_135),
.B(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_138),
.Y(n_140)
);


endmodule