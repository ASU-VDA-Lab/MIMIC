module fake_netlist_5_2118_n_633 (n_137, n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_633);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_633;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_611;
wire n_444;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_174;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_64),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_18),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_14),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_50),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_62),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_58),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_4),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_84),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_98),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_2),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_29),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_40),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_88),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_83),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_21),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_102),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_33),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_32),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_82),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_6),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_17),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_103),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_85),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_9),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_67),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_23),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_46),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_9),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_51),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_97),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_53),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_75),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_41),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_14),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_61),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_39),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_74),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_48),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_1),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_52),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_0),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_87),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_204),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_180),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_0),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

BUFx6f_ASAP7_75t_SL g214 ( 
.A(n_152),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_141),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_145),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_146),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_187),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_169),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_152),
.B(n_170),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_175),
.B(n_1),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_199),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_155),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_156),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_197),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_211),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_213),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_157),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_157),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_152),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_159),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_228),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_243),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

NAND2x1p5_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_164),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_247),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_206),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_214),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_214),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_246),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_207),
.B(n_160),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_205),
.B(n_167),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_208),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_157),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_224),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

AO22x2_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_202),
.B1(n_151),
.B2(n_143),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_171),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_226),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_242),
.B1(n_237),
.B2(n_226),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_287),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_295),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_196),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_262),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_161),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_284),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_254),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_162),
.Y(n_319)
);

BUFx4f_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_19),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_289),
.B(n_163),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_283),
.B(n_165),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_166),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_237),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g331 ( 
.A(n_267),
.B(n_242),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_168),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_254),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_290),
.A2(n_272),
.B1(n_249),
.B2(n_250),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_255),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_203),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_272),
.A2(n_198),
.B1(n_195),
.B2(n_192),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_260),
.B(n_264),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

OR2x6_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_2),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_274),
.B(n_173),
.Y(n_347)
);

BUFx4f_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

INVx4_ASAP7_75t_SL g349 ( 
.A(n_260),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_251),
.B(n_191),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_260),
.B(n_174),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_265),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_268),
.A2(n_186),
.B1(n_185),
.B2(n_184),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_276),
.B(n_176),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_280),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_270),
.B(n_181),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_266),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_271),
.B(n_178),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_277),
.C(n_298),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_279),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_285),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_302),
.B(n_285),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_311),
.A2(n_297),
.B1(n_291),
.B2(n_5),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_313),
.B(n_291),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_20),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_22),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_314),
.B(n_326),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_320),
.B(n_3),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

BUFx8_ASAP7_75t_L g378 ( 
.A(n_315),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_4),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_320),
.B(n_5),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_24),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_306),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_385)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_L g387 ( 
.A1(n_319),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_357),
.B(n_10),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_357),
.B(n_11),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_342),
.Y(n_391)
);

AND2x6_ASAP7_75t_SL g392 ( 
.A(n_346),
.B(n_13),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_25),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_26),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_335),
.B(n_15),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_27),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_305),
.B(n_28),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_323),
.B(n_30),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_328),
.B(n_89),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_15),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_16),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_336),
.B(n_90),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_300),
.B(n_91),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_354),
.B(n_16),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_300),
.B(n_31),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_324),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_304),
.B(n_37),
.Y(n_408)
);

NOR3xp33_ASAP7_75t_SL g409 ( 
.A(n_350),
.B(n_38),
.C(n_42),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_304),
.B(n_43),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_303),
.B(n_44),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_45),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_47),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_316),
.B(n_49),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_316),
.B(n_55),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_347),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_310),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_348),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_316),
.B(n_56),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_301),
.B(n_57),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_317),
.B(n_59),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_368),
.B(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_401),
.A2(n_322),
.B1(n_301),
.B2(n_346),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_368),
.B(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_382),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_391),
.B(n_317),
.Y(n_433)
);

AO22x1_ASAP7_75t_L g434 ( 
.A1(n_420),
.A2(n_322),
.B1(n_331),
.B2(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_365),
.B(n_366),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_365),
.B(n_317),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_379),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_377),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_405),
.A2(n_345),
.B1(n_344),
.B2(n_348),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_375),
.B(n_325),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_418),
.B(n_345),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_299),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_366),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_R g448 ( 
.A(n_424),
.B(n_307),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

BUFx4_ASAP7_75t_SL g450 ( 
.A(n_392),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_364),
.B(n_321),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

BUFx12f_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_371),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_413),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_412),
.B(n_338),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_321),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_349),
.Y(n_462)
);

BUFx4f_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_460),
.A2(n_421),
.B(n_404),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_431),
.A2(n_439),
.B1(n_429),
.B2(n_466),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_436),
.A2(n_421),
.B(n_394),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_381),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_431),
.A2(n_373),
.B1(n_397),
.B2(n_400),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_431),
.A2(n_373),
.B1(n_397),
.B2(n_400),
.Y(n_472)
);

AO31x2_ASAP7_75t_L g473 ( 
.A1(n_426),
.A2(n_393),
.A3(n_394),
.B(n_396),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_419),
.B(n_415),
.Y(n_474)
);

AND2x6_ASAP7_75t_SL g475 ( 
.A(n_461),
.B(n_398),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_407),
.B1(n_403),
.B2(n_370),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_376),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_386),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_443),
.A2(n_372),
.B(n_396),
.C(n_390),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_439),
.B(n_386),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_448),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_444),
.A2(n_414),
.B(n_410),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_446),
.A2(n_408),
.B(n_406),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_439),
.B(n_427),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_307),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_457),
.A2(n_338),
.B(n_332),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_442),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_489)
);

NOR2x1_ASAP7_75t_SL g490 ( 
.A(n_447),
.B(n_386),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_438),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_464),
.A2(n_386),
.B(n_349),
.Y(n_492)
);

AO31x2_ASAP7_75t_L g493 ( 
.A1(n_465),
.A2(n_386),
.A3(n_389),
.B(n_308),
.Y(n_493)
);

A2O1A1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_386),
.B(n_308),
.C(n_363),
.Y(n_494)
);

NOR2x1_ASAP7_75t_SL g495 ( 
.A(n_447),
.B(n_308),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_432),
.B(n_363),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_437),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_428),
.B1(n_459),
.B2(n_456),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_442),
.B(n_453),
.Y(n_499)
);

A2O1A1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_428),
.B(n_487),
.C(n_476),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_487),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_483),
.A2(n_440),
.B(n_441),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_474),
.A2(n_452),
.B(n_434),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_469),
.A2(n_492),
.B(n_467),
.Y(n_504)
);

OAI221xp5_ASAP7_75t_L g505 ( 
.A1(n_486),
.A2(n_455),
.B1(n_463),
.B2(n_451),
.C(n_448),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_468),
.A2(n_447),
.B(n_463),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_470),
.B(n_462),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_471),
.A2(n_447),
.B(n_451),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

O2A1O1Ixp33_ASAP7_75t_SL g510 ( 
.A1(n_494),
.A2(n_451),
.B(n_462),
.C(n_68),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_470),
.B(n_445),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_445),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_451),
.B(n_363),
.C(n_69),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_472),
.A2(n_63),
.B(n_66),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_484),
.A2(n_70),
.B(n_71),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_496),
.A2(n_72),
.B(n_73),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_76),
.B(n_79),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_454),
.Y(n_519)
);

BUFx4f_ASAP7_75t_L g520 ( 
.A(n_481),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_495),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_475),
.A2(n_80),
.B(n_81),
.C(n_86),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_501),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_490),
.B(n_473),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_512),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_502),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_482),
.Y(n_529)
);

INVx3_ASAP7_75t_SL g530 ( 
.A(n_512),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_497),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_498),
.A2(n_481),
.B1(n_493),
.B2(n_473),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_503),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_503),
.Y(n_534)
);

OAI211xp5_ASAP7_75t_L g535 ( 
.A1(n_522),
.A2(n_450),
.B(n_493),
.C(n_94),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_522),
.B(n_513),
.C(n_520),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_512),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_92),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_519),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_500),
.A2(n_505),
.B1(n_511),
.B2(n_513),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_507),
.B(n_138),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_499),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g543 ( 
.A1(n_514),
.A2(n_93),
.B(n_96),
.Y(n_543)
);

OAI221xp5_ASAP7_75t_L g544 ( 
.A1(n_510),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.C(n_106),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_516),
.A2(n_107),
.B1(n_111),
.B2(n_112),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_521),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_516),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_515),
.A2(n_120),
.B1(n_123),
.B2(n_127),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_508),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_515),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_530),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_540),
.A2(n_514),
.B1(n_517),
.B2(n_506),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_536),
.A2(n_518),
.B1(n_510),
.B2(n_506),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_526),
.A2(n_518),
.B(n_504),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_504),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_539),
.Y(n_558)
);

AOI221xp5_ASAP7_75t_L g559 ( 
.A1(n_544),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.C(n_132),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_538),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

NOR2x1_ASAP7_75t_SL g562 ( 
.A(n_535),
.B(n_137),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_546),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_538),
.A2(n_529),
.B1(n_537),
.B2(n_527),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_532),
.A2(n_545),
.B(n_547),
.C(n_538),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_539),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_530),
.A2(n_548),
.B1(n_541),
.B2(n_550),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_524),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_543),
.A2(n_548),
.B1(n_552),
.B2(n_523),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_549),
.B1(n_533),
.B2(n_534),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_572),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_557),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_561),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_568),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_553),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_570),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_559),
.A2(n_533),
.B1(n_534),
.B2(n_551),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_551),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_571),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_555),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_553),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_566),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_542),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_554),
.B(n_525),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_567),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_577),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_575),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_584),
.B(n_563),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_578),
.Y(n_593)
);

OAI33xp33_ASAP7_75t_L g594 ( 
.A1(n_582),
.A2(n_563),
.A3(n_566),
.B1(n_558),
.B2(n_542),
.B3(n_528),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_575),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_589),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_589),
.B(n_581),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_588),
.B(n_584),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_591),
.B(n_584),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_583),
.Y(n_600)
);

NAND2x1p5_ASAP7_75t_L g601 ( 
.A(n_591),
.B(n_583),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_591),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_582),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_598),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_599),
.A2(n_594),
.B1(n_587),
.B2(n_592),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_602),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_593),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_604),
.B(n_595),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_603),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_607),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_606),
.B(n_600),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_605),
.B(n_565),
.C(n_581),
.Y(n_612)
);

BUFx2_ASAP7_75t_SL g613 ( 
.A(n_609),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_612),
.B(n_590),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_610),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_615),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_614),
.B(n_612),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_L g618 ( 
.A(n_617),
.B(n_613),
.C(n_579),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_619),
.B(n_616),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_620),
.B(n_611),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_SL g622 ( 
.A(n_621),
.B(n_565),
.C(n_560),
.Y(n_622)
);

AND2x2_ASAP7_75t_SL g623 ( 
.A(n_622),
.B(n_608),
.Y(n_623)
);

AND2x4_ASAP7_75t_SL g624 ( 
.A(n_623),
.B(n_564),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_624),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_625),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_626),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_627),
.A2(n_601),
.B1(n_586),
.B2(n_576),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_627),
.B(n_562),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_628),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_630),
.Y(n_631)
);

AOI221xp5_ASAP7_75t_L g632 ( 
.A1(n_631),
.A2(n_573),
.B1(n_586),
.B2(n_556),
.C(n_578),
.Y(n_632)
);

AOI211xp5_ASAP7_75t_L g633 ( 
.A1(n_632),
.A2(n_585),
.B(n_580),
.C(n_528),
.Y(n_633)
);


endmodule