module fake_jpeg_19844_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_38),
.B1(n_41),
.B2(n_16),
.Y(n_89)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_20),
.CON(n_58),
.SN(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_16),
.B(n_21),
.C(n_17),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_65),
.B1(n_69),
.B2(n_30),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_20),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_16),
.B1(n_21),
.B2(n_17),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_42),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_75),
.B(n_80),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_85),
.Y(n_112)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_46),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_82),
.B(n_88),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_46),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_20),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_91),
.Y(n_131)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_20),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_106),
.B(n_19),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_38),
.B1(n_41),
.B2(n_17),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_41),
.B1(n_29),
.B2(n_21),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_107),
.B1(n_19),
.B2(n_23),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_44),
.C(n_39),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.C(n_44),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_26),
.B(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_44),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_108),
.Y(n_114)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_34),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_66),
.B(n_22),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_103),
.C(n_74),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_42),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_113),
.B(n_121),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_44),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_119),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_134),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_79),
.B1(n_106),
.B2(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_42),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_136),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_39),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_76),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_39),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_141),
.A2(n_34),
.B1(n_23),
.B2(n_33),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_101),
.B1(n_96),
.B2(n_83),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_137),
.B1(n_111),
.B2(n_19),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_90),
.B1(n_98),
.B2(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_90),
.B1(n_98),
.B2(n_104),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_140),
.B1(n_114),
.B2(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_119),
.B1(n_120),
.B2(n_118),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_102),
.C(n_106),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_164),
.C(n_33),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_80),
.B(n_110),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_19),
.B(n_23),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_110),
.B1(n_87),
.B2(n_70),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_172),
.B1(n_131),
.B2(n_127),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_100),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_22),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_78),
.B1(n_84),
.B2(n_97),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_139),
.B1(n_84),
.B2(n_111),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_86),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_81),
.B1(n_97),
.B2(n_85),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_34),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_91),
.B1(n_105),
.B2(n_72),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_179),
.B1(n_183),
.B2(n_199),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_203),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_116),
.B1(n_72),
.B2(n_81),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_19),
.A3(n_22),
.B1(n_116),
.B2(n_18),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_188),
.B1(n_197),
.B2(n_172),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_33),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_186),
.A2(n_168),
.B(n_25),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_162),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_19),
.B1(n_25),
.B2(n_18),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_34),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_191),
.A2(n_154),
.B(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_201),
.B1(n_143),
.B2(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_200),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_18),
.C(n_1),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_34),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_25),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_143),
.A2(n_150),
.A3(n_158),
.B1(n_149),
.B2(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_25),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_206),
.A2(n_211),
.B1(n_220),
.B2(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_200),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_217),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_174),
.A2(n_152),
.B1(n_158),
.B2(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_216),
.B(n_12),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_156),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_195),
.B1(n_177),
.B2(n_202),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_191),
.A2(n_166),
.B(n_159),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_185),
.B(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_226),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_166),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_225),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_168),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_168),
.B1(n_165),
.B2(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_176),
.C(n_18),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_198),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_244),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_213),
.Y(n_263)
);

OAI211xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_180),
.B(n_201),
.C(n_194),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_227),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_189),
.B1(n_175),
.B2(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_226),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_188),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_233),
.B1(n_223),
.B2(n_228),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_225),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_208),
.B(n_198),
.C(n_189),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_231),
.C(n_221),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_175),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_256),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_230),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_214),
.B(n_196),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_270),
.B1(n_252),
.B2(n_249),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_218),
.C(n_219),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_218),
.C(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_263),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_237),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_267),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_254),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_R g266 ( 
.A(n_256),
.B(n_210),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_266),
.A2(n_250),
.B1(n_248),
.B2(n_215),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_232),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_271),
.Y(n_288)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_235),
.A2(n_214),
.B1(n_229),
.B2(n_212),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_220),
.B1(n_242),
.B2(n_215),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_238),
.B(n_235),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_280),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_234),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_273),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_253),
.C(n_243),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_283),
.C(n_268),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_236),
.C(n_249),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_284),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_290),
.B1(n_257),
.B2(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_196),
.B1(n_244),
.B2(n_11),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_288),
.B1(n_285),
.B2(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_302),
.C(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_301),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_268),
.B(n_274),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_4),
.B(n_6),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_272),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_274),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_1),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_310),
.C(n_300),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_306),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_282),
.B1(n_5),
.B2(n_6),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_4),
.C(n_5),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_297),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_4),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_302),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_316),
.B(n_292),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_292),
.C(n_299),
.Y(n_316)
);

NAND2x1_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_304),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_7),
.B(n_8),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_305),
.B1(n_308),
.B2(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.C(n_317),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_318),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_319),
.B(n_8),
.C(n_9),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_7),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_9),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_9),
.C(n_10),
.Y(n_329)
);


endmodule