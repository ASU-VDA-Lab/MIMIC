module fake_jpeg_21567_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_26),
.B(n_29),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_26),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_4),
.B(n_5),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_52),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_54),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_24),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_55),
.C(n_61),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_30),
.B1(n_28),
.B2(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_30),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_15),
.B1(n_16),
.B2(n_12),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_60),
.B(n_6),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_12),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_21),
.C(n_13),
.Y(n_61)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_73),
.B1(n_60),
.B2(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_34),
.B(n_35),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_54),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_52),
.C(n_51),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_79),
.C(n_81),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_49),
.B1(n_51),
.B2(n_73),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_63),
.C(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_86),
.B(n_87),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_63),
.C(n_62),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_79),
.B1(n_49),
.B2(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_66),
.A3(n_78),
.B1(n_79),
.B2(n_70),
.C1(n_11),
.C2(n_10),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_71),
.B1(n_68),
.B2(n_33),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_48),
.B1(n_40),
.B2(n_34),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_40),
.B(n_33),
.C(n_50),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_62),
.C(n_50),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_95),
.C(n_21),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_89),
.C(n_91),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_45),
.B(n_57),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.C(n_56),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_100),
.A3(n_56),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_6),
.Y(n_103)
);


endmodule