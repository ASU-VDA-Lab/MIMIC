module fake_jpeg_6359_n_89 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_89);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_89;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_10),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_2),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_32),
.B(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_20),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_12),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_33),
.Y(n_35)
);

AND2x4_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_41),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_16),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_50),
.C(n_38),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_42),
.B(n_52),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_16),
.B(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_15),
.B1(n_11),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_42),
.B1(n_47),
.B2(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_51),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_27),
.B(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_61),
.B(n_51),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B1(n_36),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_45),
.B1(n_37),
.B2(n_50),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_50),
.B(n_45),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_56),
.B(n_64),
.C(n_60),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_35),
.C(n_34),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_39),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_44),
.C(n_40),
.Y(n_72)
);

NOR4xp25_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.C(n_53),
.D(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_63),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_83),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_71),
.B(n_64),
.C(n_66),
.Y(n_84)
);

OAI21x1_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_78),
.B(n_77),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_85),
.B(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_88),
.Y(n_89)
);


endmodule