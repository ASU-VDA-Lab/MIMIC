module real_jpeg_19779_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_1),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_49),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_26),
.B1(n_33),
.B2(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_44),
.B1(n_47),
.B2(n_56),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_3),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_126),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_3),
.A2(n_44),
.B1(n_47),
.B2(n_126),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_126),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_4),
.A2(n_44),
.B1(n_47),
.B2(n_131),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_131),
.Y(n_185)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_5),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_7),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_138),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_7),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_168)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_9),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_124),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_124),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_9),
.A2(n_44),
.B1(n_47),
.B2(n_124),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_10),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_14),
.B(n_62),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_10),
.A2(n_44),
.B1(n_47),
.B2(n_129),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_10),
.A2(n_104),
.B1(n_185),
.B2(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_86),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_10),
.B(n_31),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_10),
.A2(n_31),
.B(n_214),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_12),
.A2(n_36),
.B1(n_44),
.B2(n_47),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_13),
.A2(n_34),
.B1(n_44),
.B2(n_47),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_13),
.A2(n_34),
.B1(n_61),
.B2(n_62),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_14),
.A2(n_44),
.B(n_59),
.C(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_93),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_77),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_77),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_69),
.C(n_72),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_69),
.B2(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_23),
.A2(n_37),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_23),
.A2(n_37),
.B1(n_144),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_23),
.A2(n_264),
.B(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_23),
.A2(n_83),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_24),
.B(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_24),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_24),
.A2(n_29),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_25),
.B(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_26),
.B(n_129),
.CON(n_128),
.SN(n_128)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_28),
.A2(n_30),
.B1(n_128),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_29),
.B(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_30),
.A2(n_44),
.A3(n_46),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_43),
.B(n_45),
.C(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_45),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_32),
.A2(n_37),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_37),
.B(n_129),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_42),
.A2(n_51),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_43),
.A2(n_52),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_43),
.A2(n_52),
.B1(n_123),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_43),
.A2(n_52),
.B1(n_156),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_43),
.A2(n_50),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_43),
.A2(n_52),
.B1(n_75),
.B2(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_45),
.B(n_47),
.Y(n_215)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_47),
.A2(n_63),
.B(n_129),
.C(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_74),
.B(n_76),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_51),
.A2(n_76),
.B(n_87),
.Y(n_266)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_67),
.C(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_57),
.A2(n_66),
.B1(n_73),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_60),
.B(n_64),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_64),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_58),
.A2(n_60),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_58),
.A2(n_60),
.B1(n_181),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_58),
.A2(n_60),
.B1(n_203),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_58),
.A2(n_221),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_58),
.A2(n_60),
.B1(n_111),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_58),
.A2(n_119),
.B(n_256),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_60),
.B(n_129),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_61),
.B(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_65),
.B(n_120),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_69),
.C(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_69),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_72),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_73),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_315),
.A3(n_325),
.B1(n_328),
.B2(n_329),
.C(n_332),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_295),
.B(n_314),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_271),
.B(n_294),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_161),
.B(n_246),
.C(n_270),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_149),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_98),
.B(n_149),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_132),
.B2(n_148),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_101),
.B(n_116),
.C(n_148),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_110),
.B2(n_115),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_102),
.B(n_115),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B(n_107),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_106),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_109),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_104),
.A2(n_171),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_104),
.A2(n_173),
.B(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_104),
.A2(n_105),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_129),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_108),
.A2(n_169),
.B(n_206),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_112),
.B(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_127),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_141),
.C(n_146),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_136),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_150),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_155),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_157),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_245),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_239),
.B(n_244),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_226),
.B(n_238),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_208),
.B(n_225),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_195),
.B(n_207),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_182),
.B(n_194),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_178),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_189),
.B(n_193),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_188),
.Y(n_193)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_197),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_206),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_210),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_216),
.B1(n_223),
.B2(n_224),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_234),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_235),
.C(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_248),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_268),
.B2(n_269),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_258),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_258),
.C(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_267),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_266),
.C(n_267),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_293),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_286),
.B2(n_287),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_287),
.C(n_293),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_281),
.C(n_285),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_279),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_284),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_289),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_305),
.B(n_309),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_291),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_297),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_312),
.B2(n_313),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_304),
.C(n_313),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B(n_303),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_317),
.C(n_322),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_303),
.B(n_317),
.CI(n_322),
.CON(n_327),
.SN(n_327)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_323),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_323),
.Y(n_329)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_327),
.Y(n_331)
);


endmodule