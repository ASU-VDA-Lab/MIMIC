module real_jpeg_33327_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_316, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_316;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_0),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_0),
.Y(n_164)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_142),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_4),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_5),
.A2(n_52),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_5),
.A2(n_52),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_6),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_6),
.Y(n_107)
);

OAI22x1_ASAP7_75t_L g152 ( 
.A1(n_6),
.A2(n_107),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_107),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_7),
.A2(n_139),
.B1(n_142),
.B2(n_146),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_8),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_92),
.B1(n_96),
.B2(n_101),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_9),
.B(n_188),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_9),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_9),
.B(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_10),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_58),
.B1(n_62),
.B2(n_64),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_64),
.B1(n_247),
.B2(n_252),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_216),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_215),
.Y(n_14)
);

INVxp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_165),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_17),
.B(n_165),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_65),
.C(n_113),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_18),
.B(n_66),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_47),
.B1(n_56),
.B2(n_57),
.Y(n_18)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_19),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g297 ( 
.A1(n_19),
.A2(n_47),
.B1(n_233),
.B2(n_298),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_34),
.Y(n_19)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_20),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_24),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_24),
.Y(n_162)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_24),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_24),
.Y(n_271)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_28),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_33),
.Y(n_225)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_33),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_55),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_57),
.A2(n_168),
.B(n_170),
.Y(n_167)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_91),
.B(n_102),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_68),
.B(n_104),
.Y(n_214)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_83),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_80),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_82),
.Y(n_213)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_94),
.Y(n_211)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_98),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_101),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_101),
.B(n_237),
.Y(n_236)
);

OA21x2_ASAP7_75t_R g259 ( 
.A1(n_101),
.A2(n_260),
.B(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_101),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_114),
.A2(n_115),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_136),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_136),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_124),
.B2(n_130),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_129),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2x1_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_151),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_147),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_138),
.A2(n_160),
.B1(n_196),
.B2(n_202),
.Y(n_195)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_139),
.B(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_145),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_151),
.A2(n_223),
.B(n_227),
.Y(n_222)
);

NAND2x1_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_160),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_152),
.B(n_238),
.Y(n_241)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_159),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_160),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_185),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g258 ( 
.A1(n_168),
.A2(n_170),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_171),
.Y(n_298)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_205),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B(n_214),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g301 ( 
.A(n_206),
.Y(n_301)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI321xp33_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_294),
.A3(n_306),
.B1(n_312),
.B2(n_314),
.C(n_316),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_243),
.C(n_257),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_234),
.B(n_242),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_232),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_240),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_240),
.A2(n_241),
.B(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_268),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_279),
.B1(n_280),
.B2(n_285),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.C(n_302),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_300),
.Y(n_311)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);


endmodule