module real_aes_5420_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_958, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_958;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_954;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_922;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g273 ( .A(n_0), .Y(n_273) );
INVx1_ASAP7_75t_L g669 ( .A(n_1), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_2), .A2(n_17), .B1(n_138), .B2(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g643 ( .A(n_3), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_4), .B(n_123), .Y(n_249) );
INVx1_ASAP7_75t_SL g593 ( .A(n_5), .Y(n_593) );
BUFx2_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g920 ( .A(n_6), .Y(n_920) );
INVxp67_ASAP7_75t_L g931 ( .A(n_6), .Y(n_931) );
NAND3xp33_ASAP7_75t_SL g950 ( .A(n_6), .B(n_951), .C(n_952), .Y(n_950) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_7), .B(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_8), .A2(n_39), .B1(n_122), .B2(n_235), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_9), .A2(n_45), .B1(n_157), .B2(n_184), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_10), .A2(n_66), .B1(n_192), .B2(n_295), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_11), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g267 ( .A(n_12), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_13), .B(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_14), .A2(n_54), .B1(n_193), .B2(n_251), .Y(n_621) );
INVx1_ASAP7_75t_L g271 ( .A(n_15), .Y(n_271) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_16), .A2(n_70), .B(n_148), .Y(n_147) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_16), .A2(n_70), .B(n_148), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_18), .A2(n_68), .B1(n_192), .B2(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_19), .B(n_159), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_20), .A2(n_82), .B1(n_236), .B2(n_246), .Y(n_640) );
INVx2_ASAP7_75t_L g585 ( .A(n_21), .Y(n_585) );
INVx1_ASAP7_75t_L g264 ( .A(n_22), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_23), .A2(n_26), .B1(n_216), .B2(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g923 ( .A(n_24), .Y(n_923) );
BUFx8_ASAP7_75t_SL g925 ( .A(n_24), .Y(n_925) );
O2A1O1Ixp5_ASAP7_75t_L g581 ( .A1(n_25), .A2(n_129), .B(n_184), .C(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_27), .A2(n_63), .B1(n_185), .B2(n_555), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_28), .Y(n_613) );
AO22x1_ASAP7_75t_L g244 ( .A1(n_29), .A2(n_80), .B1(n_140), .B2(n_245), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_30), .Y(n_127) );
AND2x2_ASAP7_75t_L g156 ( .A(n_31), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_32), .B(n_140), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_33), .A2(n_83), .B1(n_628), .B2(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g903 ( .A(n_34), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_34), .B(n_905), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_34), .A2(n_87), .B1(n_903), .B2(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g915 ( .A(n_35), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_35), .B(n_81), .Y(n_949) );
INVx1_ASAP7_75t_L g576 ( .A(n_36), .Y(n_576) );
AOI22x1_ASAP7_75t_L g190 ( .A1(n_37), .A2(n_99), .B1(n_191), .B2(n_192), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_38), .B(n_195), .Y(n_237) );
AND2x2_ASAP7_75t_L g952 ( .A(n_40), .B(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_41), .B(n_573), .Y(n_664) );
INVx2_ASAP7_75t_L g583 ( .A(n_42), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_43), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_44), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g556 ( .A(n_46), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_47), .B(n_219), .Y(n_662) );
INVx1_ASAP7_75t_SL g596 ( .A(n_48), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_49), .B(n_216), .Y(n_215) );
AOI22x1_ASAP7_75t_L g105 ( .A1(n_50), .A2(n_106), .B1(n_906), .B2(n_916), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_51), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g609 ( .A(n_52), .Y(n_609) );
INVx1_ASAP7_75t_L g148 ( .A(n_53), .Y(n_148) );
AND2x4_ASAP7_75t_L g144 ( .A(n_55), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g579 ( .A(n_55), .B(n_145), .Y(n_579) );
INVx1_ASAP7_75t_L g599 ( .A(n_56), .Y(n_599) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
INVx2_ASAP7_75t_L g297 ( .A(n_58), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_59), .A2(n_103), .B1(n_944), .B2(n_954), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_60), .A2(n_75), .B1(n_122), .B2(n_191), .Y(n_231) );
CKINVDCx14_ASAP7_75t_R g253 ( .A(n_61), .Y(n_253) );
AND2x2_ASAP7_75t_L g165 ( .A(n_62), .B(n_140), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_64), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_65), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_67), .B(n_208), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_69), .B(n_152), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_71), .A2(n_86), .B1(n_909), .B2(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_71), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_72), .B(n_942), .Y(n_941) );
CKINVDCx14_ASAP7_75t_R g199 ( .A(n_73), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_74), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_76), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_77), .B(n_123), .Y(n_213) );
OR2x6_ASAP7_75t_L g912 ( .A(n_78), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g951 ( .A(n_78), .Y(n_951) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_79), .B(n_217), .Y(n_597) );
INVx1_ASAP7_75t_L g914 ( .A(n_81), .Y(n_914) );
INVx1_ASAP7_75t_L g953 ( .A(n_84), .Y(n_953) );
BUFx5_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx1_ASAP7_75t_L g187 ( .A(n_85), .Y(n_187) );
INVx1_ASAP7_75t_L g910 ( .A(n_86), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_87), .Y(n_939) );
INVx2_ASAP7_75t_L g275 ( .A(n_88), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_89), .B(n_562), .Y(n_594) );
INVx2_ASAP7_75t_L g559 ( .A(n_90), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_91), .Y(n_937) );
NAND2xp33_ASAP7_75t_L g161 ( .A(n_92), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g565 ( .A(n_93), .Y(n_565) );
INVx2_ASAP7_75t_L g616 ( .A(n_94), .Y(n_616) );
INVx2_ASAP7_75t_SL g145 ( .A(n_95), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_96), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_97), .B(n_168), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_98), .B(n_208), .Y(n_657) );
AO32x2_ASAP7_75t_L g539 ( .A1(n_100), .A2(n_143), .A3(n_540), .B1(n_546), .B2(n_547), .Y(n_539) );
AO22x2_ASAP7_75t_L g746 ( .A1(n_100), .A2(n_540), .B1(n_747), .B2(n_749), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_101), .B(n_150), .Y(n_149) );
AO21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_923), .B(n_924), .Y(n_103) );
NAND2x1p5_ASAP7_75t_SL g104 ( .A(n_105), .B(n_921), .Y(n_104) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g921 ( .A(n_107), .B(n_922), .Y(n_921) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_531), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx8_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AOI31xp33_ASAP7_75t_L g532 ( .A1(n_111), .A2(n_533), .A3(n_800), .B(n_903), .Y(n_532) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_426), .Y(n_112) );
NAND4xp25_ASAP7_75t_SL g113 ( .A(n_114), .B(n_317), .C(n_363), .D(n_395), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_255), .B(n_276), .Y(n_114) );
OAI21xp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_201), .B(n_222), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_116), .A2(n_375), .B1(n_379), .B2(n_381), .Y(n_374) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_178), .Y(n_117) );
INVx2_ASAP7_75t_L g307 ( .A(n_118), .Y(n_307) );
AND2x2_ASAP7_75t_L g424 ( .A(n_118), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_154), .Y(n_118) );
AND2x2_ASAP7_75t_L g341 ( .A(n_119), .B(n_226), .Y(n_341) );
AND2x2_ASAP7_75t_L g391 ( .A(n_119), .B(n_361), .Y(n_391) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_119), .B(n_180), .Y(n_418) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_146), .B(n_149), .Y(n_119) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_120), .A2(n_146), .B(n_149), .Y(n_286) );
OAI21x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_135), .B(n_143), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_129), .B2(n_131), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g140 ( .A(n_124), .Y(n_140) );
INVx2_ASAP7_75t_L g193 ( .A(n_124), .Y(n_193) );
INVx2_ASAP7_75t_L g219 ( .A(n_124), .Y(n_219) );
INVx2_ASAP7_75t_L g544 ( .A(n_124), .Y(n_544) );
INVx1_ASAP7_75t_L g666 ( .A(n_124), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_L g182 ( .A1(n_128), .A2(n_183), .B1(n_188), .B2(n_190), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_128), .B(n_578), .Y(n_611) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_129), .A2(n_212), .B(n_213), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_129), .B(n_229), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_129), .A2(n_541), .B1(n_543), .B2(n_545), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_129), .A2(n_660), .B(n_662), .Y(n_659) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_130), .Y(n_142) );
INVxp67_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
INVx1_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_130), .B(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_130), .B(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g270 ( .A(n_130), .Y(n_270) );
INVx3_ASAP7_75t_L g301 ( .A(n_130), .Y(n_301) );
INVx1_ASAP7_75t_L g607 ( .A(n_132), .Y(n_607) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g629 ( .A(n_133), .Y(n_629) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g138 ( .A(n_134), .Y(n_138) );
INVx6_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
INVx3_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B(n_141), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_137), .B(n_266), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_137), .A2(n_140), .B1(n_269), .B2(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g577 ( .A(n_137), .Y(n_577) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_138), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_140), .A2(n_301), .B(n_596), .C(n_597), .Y(n_595) );
INVxp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_SL g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g220 ( .A(n_142), .Y(n_220) );
INVx1_ASAP7_75t_L g243 ( .A(n_142), .Y(n_243) );
INVx1_ASAP7_75t_L g545 ( .A(n_142), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_142), .A2(n_559), .B(n_560), .C(n_561), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_142), .A2(n_592), .B(n_593), .C(n_594), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_142), .B(n_623), .Y(n_622) );
AO31x2_ASAP7_75t_L g181 ( .A1(n_143), .A2(n_182), .A3(n_194), .B(n_198), .Y(n_181) );
AO31x2_ASAP7_75t_L g288 ( .A1(n_143), .A2(n_182), .A3(n_194), .B(n_198), .Y(n_288) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx3_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
INVx1_ASAP7_75t_L g241 ( .A(n_144), .Y(n_241) );
AND2x2_ASAP7_75t_L g638 ( .A(n_144), .B(n_173), .Y(n_638) );
AND2x2_ASAP7_75t_L g747 ( .A(n_144), .B(n_748), .Y(n_747) );
INVx3_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx2_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
OR2x2_ASAP7_75t_L g240 ( .A(n_150), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x2_ASAP7_75t_L g296 ( .A(n_151), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
OR2x2_ASAP7_75t_L g343 ( .A(n_154), .B(n_288), .Y(n_343) );
AND2x2_ASAP7_75t_L g366 ( .A(n_154), .B(n_288), .Y(n_366) );
AND2x4_ASAP7_75t_L g412 ( .A(n_154), .B(n_285), .Y(n_412) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_164), .B(n_172), .Y(n_154) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_155), .A2(n_164), .B(n_172), .Y(n_282) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B(n_163), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_157), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_158), .A2(n_544), .B1(n_613), .B2(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_158), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
INVx1_ASAP7_75t_L g168 ( .A(n_159), .Y(n_168) );
INVx2_ASAP7_75t_SL g542 ( .A(n_159), .Y(n_542) );
INVx1_ASAP7_75t_L g555 ( .A(n_159), .Y(n_555) );
INVx2_ASAP7_75t_L g571 ( .A(n_159), .Y(n_571) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
OAI21x1_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_170), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_169), .B(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g177 ( .A(n_169), .Y(n_177) );
AOI21x1_ASAP7_75t_L g248 ( .A1(n_171), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp33_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_175), .B(n_177), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_174), .B(n_230), .Y(n_590) );
NAND3xp33_ASAP7_75t_SL g293 ( .A(n_175), .B(n_260), .C(n_270), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_175), .B(n_260), .C(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2x1_ASAP7_75t_L g221 ( .A(n_176), .B(n_208), .Y(n_221) );
INVx1_ASAP7_75t_L g305 ( .A(n_178), .Y(n_305) );
AND2x2_ASAP7_75t_L g486 ( .A(n_178), .B(n_412), .Y(n_486) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g254 ( .A(n_179), .Y(n_254) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g413 ( .A(n_180), .B(n_402), .Y(n_413) );
INVx1_ASAP7_75t_L g481 ( .A(n_180), .Y(n_481) );
AND2x2_ASAP7_75t_L g528 ( .A(n_180), .B(n_282), .Y(n_528) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g467 ( .A(n_181), .B(n_334), .Y(n_467) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g562 ( .A(n_186), .Y(n_562) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g247 ( .A(n_187), .Y(n_247) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_189), .B(n_229), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_189), .B(n_623), .Y(n_631) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_196), .B(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_SL g598 ( .A(n_196), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_197), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g260 ( .A(n_197), .Y(n_260) );
INVx1_ASAP7_75t_L g548 ( .A(n_197), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_197), .B(n_230), .Y(n_563) );
NOR2xp67_ASAP7_75t_L g623 ( .A(n_197), .B(n_230), .Y(n_623) );
BUFx3_ASAP7_75t_L g625 ( .A(n_197), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_197), .B(n_230), .Y(n_670) );
INVx1_ASAP7_75t_L g748 ( .A(n_197), .Y(n_748) );
NOR2xp67_ASAP7_75t_SL g198 ( .A(n_199), .B(n_200), .Y(n_198) );
OR2x2_ASAP7_75t_L g252 ( .A(n_200), .B(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g650 ( .A1(n_200), .A2(n_602), .B(n_615), .Y(n_650) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g437 ( .A(n_204), .B(n_325), .Y(n_437) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g355 ( .A(n_205), .B(n_239), .Y(n_355) );
AND2x2_ASAP7_75t_L g387 ( .A(n_205), .B(n_291), .Y(n_387) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g238 ( .A(n_206), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g315 ( .A(n_206), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g370 ( .A(n_206), .Y(n_370) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_210), .Y(n_206) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_209), .B(n_275), .Y(n_274) );
BUFx3_ASAP7_75t_L g546 ( .A(n_209), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_209), .B(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_209), .B(n_643), .Y(n_642) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_221), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_218), .B(n_220), .Y(n_214) );
INVx1_ASAP7_75t_L g592 ( .A(n_216), .Y(n_592) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g236 ( .A(n_217), .Y(n_236) );
INVx1_ASAP7_75t_L g251 ( .A(n_217), .Y(n_251) );
INVx1_ASAP7_75t_L g661 ( .A(n_217), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_254), .Y(n_222) );
INVx1_ASAP7_75t_L g484 ( .A(n_223), .Y(n_484) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_238), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g365 ( .A(n_225), .Y(n_365) );
INVx1_ASAP7_75t_L g408 ( .A(n_225), .Y(n_408) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g309 ( .A(n_226), .Y(n_309) );
AND2x2_ASAP7_75t_L g333 ( .A(n_226), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_226), .B(n_281), .Y(n_380) );
INVx2_ASAP7_75t_L g402 ( .A(n_226), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_227), .B(n_232), .Y(n_226) );
AND2x2_ASAP7_75t_L g361 ( .A(n_227), .B(n_232), .Y(n_361) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_231), .Y(n_227) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_237), .Y(n_232) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g295 ( .A(n_236), .Y(n_295) );
AND2x2_ASAP7_75t_L g289 ( .A(n_238), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g327 ( .A(n_238), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_238), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_SL g316 ( .A(n_239), .Y(n_316) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_242), .B(n_252), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_240), .A2(n_242), .B(n_252), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_241), .B(n_259), .Y(n_258) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_248), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_243), .A2(n_300), .B1(n_640), .B2(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g560 ( .A(n_247), .Y(n_560) );
OR2x2_ASAP7_75t_L g331 ( .A(n_254), .B(n_332), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_255), .B(n_526), .C(n_529), .Y(n_525) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g471 ( .A(n_256), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g475 ( .A(n_256), .B(n_376), .Y(n_475) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g290 ( .A(n_257), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g313 ( .A(n_257), .Y(n_313) );
OR2x2_ASAP7_75t_L g347 ( .A(n_257), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g354 ( .A(n_257), .Y(n_354) );
AND2x2_ASAP7_75t_L g386 ( .A(n_257), .B(n_316), .Y(n_386) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B(n_274), .Y(n_257) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND3xp33_ASAP7_75t_SL g261 ( .A(n_262), .B(n_265), .C(n_268), .Y(n_261) );
NOR2xp33_ASAP7_75t_SL g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_270), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g573 ( .A(n_270), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_270), .B(n_669), .Y(n_668) );
AOI31xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_303), .A3(n_308), .B(n_310), .Y(n_276) );
INVx1_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_283), .B(n_289), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g512 ( .A(n_280), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVxp67_ASAP7_75t_L g362 ( .A(n_282), .Y(n_362) );
INVx2_ASAP7_75t_L g394 ( .A(n_282), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_283), .B(n_308), .Y(n_320) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_283), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_285), .Y(n_400) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g334 ( .A(n_286), .Y(n_334) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g393 ( .A(n_288), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g323 ( .A(n_290), .B(n_324), .Y(n_323) );
NAND2x1_ASAP7_75t_SL g388 ( .A(n_290), .B(n_315), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_290), .B(n_376), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_290), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g516 ( .A(n_290), .Y(n_516) );
INVx2_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
AND2x2_ASAP7_75t_L g329 ( .A(n_291), .B(n_313), .Y(n_329) );
INVx1_ASAP7_75t_L g339 ( .A(n_291), .Y(n_339) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_291), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_291), .Y(n_357) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_291), .Y(n_373) );
INVx1_ASAP7_75t_L g436 ( .A(n_291), .Y(n_436) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_298), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_296), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_300), .B(n_578), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_300), .B(n_578), .C(n_609), .Y(n_608) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_301), .A2(n_554), .B(n_556), .C(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g518 ( .A(n_307), .B(n_425), .Y(n_518) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_310), .A2(n_399), .B1(n_401), .B2(n_403), .Y(n_398) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
AND2x2_ASAP7_75t_L g404 ( .A(n_312), .B(n_376), .Y(n_404) );
AND2x2_ASAP7_75t_L g502 ( .A(n_312), .B(n_355), .Y(n_502) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g356 ( .A(n_315), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g325 ( .A(n_316), .Y(n_325) );
INVx1_ASAP7_75t_L g472 ( .A(n_316), .Y(n_472) );
AOI221x1_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_330), .C(n_335), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_323), .A2(n_337), .B1(n_415), .B2(n_416), .Y(n_414) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
OR2x2_ASAP7_75t_L g422 ( .A(n_327), .B(n_338), .Y(n_422) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g421 ( .A(n_329), .B(n_355), .Y(n_421) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g444 ( .A(n_333), .Y(n_444) );
INVx1_ASAP7_75t_L g350 ( .A(n_334), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_334), .B(n_402), .Y(n_513) );
OAI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B1(n_344), .B2(n_349), .C(n_351), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_SL g381 ( .A(n_338), .B(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_338), .Y(n_483) );
OR2x2_ASAP7_75t_L g521 ( .A(n_338), .B(n_437), .Y(n_521) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g345 ( .A(n_339), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_341), .B(n_392), .Y(n_458) );
AND2x2_ASAP7_75t_L g480 ( .A(n_341), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_341), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g407 ( .A(n_342), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_342), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g349 ( .A(n_343), .B(n_350), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_343), .A2(n_384), .B1(n_388), .B2(n_389), .Y(n_383) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_345), .A2(n_450), .B(n_455), .Y(n_449) );
AND2x2_ASAP7_75t_L g410 ( .A(n_346), .B(n_373), .Y(n_410) );
INVx1_ASAP7_75t_L g509 ( .A(n_346), .Y(n_509) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g369 ( .A(n_347), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g454 ( .A(n_348), .Y(n_454) );
AND3x2_ASAP7_75t_L g358 ( .A(n_350), .B(n_359), .C(n_362), .Y(n_358) );
OR2x2_ASAP7_75t_L g379 ( .A(n_350), .B(n_380), .Y(n_379) );
OAI21xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_356), .B(n_358), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx2_ASAP7_75t_L g378 ( .A(n_353), .Y(n_378) );
INVx2_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
INVx1_ASAP7_75t_L g440 ( .A(n_355), .Y(n_440) );
AND2x2_ASAP7_75t_L g488 ( .A(n_357), .B(n_370), .Y(n_488) );
AND2x2_ASAP7_75t_L g430 ( .A(n_359), .B(n_393), .Y(n_430) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g417 ( .A(n_360), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g425 ( .A(n_360), .Y(n_425) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B(n_374), .C(n_383), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g405 ( .A1(n_369), .A2(n_406), .B1(n_409), .B2(n_411), .C(n_414), .Y(n_405) );
INVxp67_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
INVx2_ASAP7_75t_L g376 ( .A(n_370), .Y(n_376) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_370), .Y(n_470) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_371), .Y(n_496) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
OR2x2_ASAP7_75t_L g520 ( .A(n_376), .B(n_378), .Y(n_520) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g501 ( .A(n_380), .Y(n_501) );
OR2x2_ASAP7_75t_L g515 ( .A(n_382), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_386), .B(n_436), .Y(n_460) );
BUFx3_ASAP7_75t_L g489 ( .A(n_386), .Y(n_489) );
INVx2_ASAP7_75t_L g508 ( .A(n_387), .Y(n_508) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp67_ASAP7_75t_SL g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AND2x4_ASAP7_75t_L g455 ( .A(n_391), .B(n_393), .Y(n_455) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g478 ( .A(n_393), .Y(n_478) );
INVx1_ASAP7_75t_L g466 ( .A(n_394), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_405), .C(n_419), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g415 ( .A(n_402), .B(n_412), .Y(n_415) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_408), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g494 ( .A(n_408), .Y(n_494) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
BUFx3_ASAP7_75t_L g448 ( .A(n_412), .Y(n_448) );
AND2x4_ASAP7_75t_SL g495 ( .A(n_412), .B(n_481), .Y(n_495) );
INVx2_ASAP7_75t_L g433 ( .A(n_413), .Y(n_433) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_418), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_423), .Y(n_419) );
OAI222xp33_ASAP7_75t_L g461 ( .A1(n_420), .A2(n_462), .B1(n_468), .B2(n_473), .C1(n_477), .C2(n_479), .Y(n_461) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_490), .Y(n_426) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_428), .B(n_445), .C(n_461), .D(n_482), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_429), .B(n_438), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_432), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g476 ( .A(n_436), .B(n_454), .Y(n_476) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .C(n_456), .Y(n_445) );
INVx2_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_463), .B(n_494), .Y(n_524) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI32xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .A3(n_485), .B1(n_487), .B2(n_958), .Y(n_482) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_487), .A2(n_507), .B1(n_523), .B2(n_524), .C(n_525), .Y(n_522) );
NAND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AOI211x1_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_497), .B(n_499), .C(n_522), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp67_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .C(n_510), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_514), .B1(n_517), .B2(n_519), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_904), .Y(n_531) );
INVxp33_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g905 ( .A(n_534), .B(n_801), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_731), .Y(n_534) );
NOR3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_681), .C(n_709), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_586), .B1(n_632), .B2(n_644), .C(n_651), .Y(n_536) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_537), .A2(n_682), .B(n_684), .C(n_695), .Y(n_681) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_549), .Y(n_537) );
AND2x2_ASAP7_75t_L g680 ( .A(n_538), .B(n_673), .Y(n_680) );
AND2x2_ASAP7_75t_L g711 ( .A(n_538), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g739 ( .A(n_538), .Y(n_739) );
AND2x4_ASAP7_75t_L g805 ( .A(n_538), .B(n_752), .Y(n_805) );
INVx1_ASAP7_75t_L g828 ( .A(n_538), .Y(n_828) );
AND2x2_ASAP7_75t_SL g833 ( .A(n_538), .B(n_550), .Y(n_833) );
AND2x2_ASAP7_75t_L g886 ( .A(n_538), .B(n_794), .Y(n_886) );
BUFx8_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g703 ( .A(n_539), .Y(n_703) );
AND2x2_ASAP7_75t_L g773 ( .A(n_539), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_542), .B(n_583), .Y(n_582) );
AO31x2_ASAP7_75t_L g567 ( .A1(n_546), .A2(n_568), .A3(n_580), .B(n_584), .Y(n_567) );
INVx2_ASAP7_75t_L g749 ( .A(n_546), .Y(n_749) );
INVxp67_ASAP7_75t_L g601 ( .A(n_547), .Y(n_601) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_548), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g633 ( .A(n_550), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g694 ( .A(n_550), .B(n_635), .Y(n_694) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_566), .Y(n_550) );
INVx2_ASAP7_75t_L g674 ( .A(n_551), .Y(n_674) );
BUFx3_ASAP7_75t_L g699 ( .A(n_551), .Y(n_699) );
INVx1_ASAP7_75t_L g755 ( .A(n_551), .Y(n_755) );
AND2x2_ASAP7_75t_L g794 ( .A(n_551), .B(n_567), .Y(n_794) );
AND2x4_ASAP7_75t_L g891 ( .A(n_551), .B(n_703), .Y(n_891) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_558), .A3(n_563), .B(n_564), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_560), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g673 ( .A(n_567), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g705 ( .A(n_567), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_567), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g810 ( .A(n_567), .B(n_714), .Y(n_810) );
AOI221x1_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B1(n_575), .B2(n_577), .C(n_578), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g575 ( .A(n_573), .B(n_576), .Y(n_575) );
INVx4_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_617), .Y(n_587) );
AND2x2_ASAP7_75t_L g799 ( .A(n_588), .B(n_721), .Y(n_799) );
AND2x2_ASAP7_75t_L g806 ( .A(n_588), .B(n_717), .Y(n_806) );
INVx1_ASAP7_75t_L g869 ( .A(n_588), .Y(n_869) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_600), .Y(n_588) );
INVx2_ASAP7_75t_L g649 ( .A(n_589), .Y(n_649) );
INVx1_ASAP7_75t_L g671 ( .A(n_589), .Y(n_671) );
INVx2_ASAP7_75t_L g688 ( .A(n_589), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_589), .Y(n_693) );
OR2x2_ASAP7_75t_L g814 ( .A(n_589), .B(n_650), .Y(n_814) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_589), .Y(n_855) );
AO31x2_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .A3(n_595), .B(n_598), .Y(n_589) );
AND2x2_ASAP7_75t_L g707 ( .A(n_600), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g736 ( .A(n_600), .B(n_722), .Y(n_736) );
AND2x2_ASAP7_75t_L g743 ( .A(n_600), .B(n_618), .Y(n_743) );
AND2x2_ASAP7_75t_L g879 ( .A(n_600), .B(n_678), .Y(n_879) );
AO21x2_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_615), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_610), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_607), .B2(n_608), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g646 ( .A(n_617), .Y(n_646) );
AND2x2_ASAP7_75t_L g685 ( .A(n_617), .B(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_618), .Y(n_728) );
AND2x2_ASAP7_75t_L g784 ( .A(n_618), .B(n_679), .Y(n_784) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g717 ( .A(n_619), .B(n_656), .Y(n_717) );
AND2x2_ASAP7_75t_L g721 ( .A(n_619), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g764 ( .A(n_619), .Y(n_764) );
INVx1_ASAP7_75t_L g823 ( .A(n_619), .Y(n_823) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_620), .B(n_626), .Y(n_619) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_620), .B(n_626), .Y(n_654) );
OA21x2_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_624), .Y(n_620) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI21xp33_ASAP7_75t_SL g804 ( .A1(n_633), .A2(n_805), .B(n_806), .Y(n_804) );
NAND2x1p5_ASAP7_75t_L g816 ( .A(n_634), .B(n_794), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_634), .B(n_745), .Y(n_870) );
INVx4_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g672 ( .A(n_635), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g697 ( .A(n_635), .Y(n_697) );
HB1xp67_ASAP7_75t_SL g831 ( .A(n_635), .Y(n_831) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g774 ( .A(n_636), .Y(n_774) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g714 ( .A(n_637), .Y(n_714) );
INVx1_ASAP7_75t_L g753 ( .A(n_637), .Y(n_753) );
AOI21x1_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_642), .Y(n_637) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
NOR2x1p5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g716 ( .A(n_648), .B(n_717), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g758 ( .A(n_648), .B(n_759), .Y(n_758) );
AND2x4_ASAP7_75t_L g819 ( .A(n_648), .B(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_649), .Y(n_676) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_649), .Y(n_841) );
INVx2_ASAP7_75t_L g679 ( .A(n_650), .Y(n_679) );
BUFx2_ASAP7_75t_L g720 ( .A(n_650), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_672), .B1(n_675), .B2(n_680), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_671), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_653), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g708 ( .A(n_654), .Y(n_708) );
INVx1_ASAP7_75t_L g759 ( .A(n_654), .Y(n_759) );
AND2x2_ASAP7_75t_L g771 ( .A(n_654), .B(n_655), .Y(n_771) );
INVx1_ASAP7_75t_L g826 ( .A(n_655), .Y(n_826) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g678 ( .A(n_656), .Y(n_678) );
INVx2_ASAP7_75t_L g722 ( .A(n_656), .Y(n_722) );
AND2x2_ASAP7_75t_L g742 ( .A(n_656), .B(n_688), .Y(n_742) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_656), .Y(n_783) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_663), .B(n_670), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g683 ( .A(n_671), .B(n_678), .Y(n_683) );
AND2x2_ASAP7_75t_L g738 ( .A(n_673), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g772 ( .A(n_673), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g797 ( .A(n_673), .B(n_761), .Y(n_797) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_673), .Y(n_835) );
AND2x4_ASAP7_75t_L g745 ( .A(n_674), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g787 ( .A(n_674), .B(n_753), .Y(n_787) );
NOR2xp67_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g730 ( .A(n_678), .Y(n_730) );
AND2x4_ASAP7_75t_L g686 ( .A(n_679), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g706 ( .A(n_683), .B(n_707), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B(n_694), .Y(n_684) );
AND2x4_ASAP7_75t_L g729 ( .A(n_686), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g768 ( .A(n_686), .B(n_721), .Y(n_768) );
AND2x2_ASAP7_75t_L g770 ( .A(n_686), .B(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_686), .B(n_759), .Y(n_871) );
INVx1_ASAP7_75t_L g883 ( .A(n_686), .Y(n_883) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g789 ( .A(n_692), .B(n_783), .Y(n_789) );
AND2x2_ASAP7_75t_L g878 ( .A(n_692), .B(n_823), .Y(n_878) );
INVxp67_ASAP7_75t_L g894 ( .A(n_692), .Y(n_894) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_700), .B(n_706), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
AND2x2_ASAP7_75t_L g760 ( .A(n_698), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g856 ( .A(n_698), .Y(n_856) );
AND2x2_ASAP7_75t_L g881 ( .A(n_698), .B(n_809), .Y(n_881) );
INVx2_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_L g865 ( .A(n_699), .B(n_746), .Y(n_865) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_701), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_703), .B(n_705), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_703), .B(n_774), .Y(n_847) );
INVx2_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g752 ( .A(n_705), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g857 ( .A(n_705), .Y(n_857) );
OAI22xp33_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_715), .B1(n_723), .B2(n_726), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g868 ( .A(n_713), .Y(n_868) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_714), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_718), .A2(n_770), .B1(n_772), .B2(n_775), .Y(n_769) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
NAND5xp2_ASAP7_75t_L g853 ( .A(n_719), .B(n_826), .C(n_854), .D(n_856), .E(n_857), .Y(n_853) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_720), .B(n_721), .Y(n_899) );
NAND2xp67_ASAP7_75t_L g812 ( .A(n_721), .B(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g893 ( .A(n_721), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g776 ( .A(n_725), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g734 ( .A(n_728), .B(n_735), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_765), .C(n_790), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_737), .B1(n_740), .B2(n_744), .C(n_750), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_733), .A2(n_899), .B(n_900), .Y(n_898) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
OR2x6_ASAP7_75t_L g840 ( .A(n_736), .B(n_841), .Y(n_840) );
INVxp67_ASAP7_75t_L g851 ( .A(n_736), .Y(n_851) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
AND2x2_ASAP7_75t_L g763 ( .A(n_742), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g837 ( .A(n_742), .B(n_784), .Y(n_837) );
AND2x4_ASAP7_75t_L g788 ( .A(n_743), .B(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_744), .B(n_809), .Y(n_808) );
INVx4_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_745), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g901 ( .A(n_745), .B(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g756 ( .A(n_746), .Y(n_756) );
INVx1_ASAP7_75t_L g795 ( .A(n_746), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_757), .B1(n_760), .B2(n_762), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_752), .Y(n_780) );
AND2x2_ASAP7_75t_L g890 ( .A(n_752), .B(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g761 ( .A(n_753), .Y(n_761) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_753), .Y(n_820) );
INVx1_ASAP7_75t_L g766 ( .A(n_754), .Y(n_766) );
AND2x2_ASAP7_75t_L g843 ( .A(n_754), .B(n_844), .Y(n_843) );
AND2x4_ASAP7_75t_SL g754 ( .A(n_755), .B(n_756), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_757), .A2(n_808), .B1(n_811), .B2(n_815), .Y(n_807) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g844 ( .A(n_761), .Y(n_844) );
BUFx3_ASAP7_75t_L g885 ( .A(n_761), .Y(n_885) );
BUFx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g850 ( .A(n_764), .Y(n_850) );
OAI211xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B(n_769), .C(n_778), .Y(n_765) );
OAI322xp33_ASAP7_75t_L g866 ( .A1(n_766), .A2(n_840), .A3(n_867), .B1(n_869), .B2(n_870), .C1(n_871), .C2(n_872), .Y(n_866) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g791 ( .A(n_770), .Y(n_791) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_777), .B(n_865), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_781), .B1(n_785), .B2(n_788), .Y(n_778) );
AND2x4_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B1(n_796), .B2(n_798), .Y(n_790) );
OAI32xp33_ASAP7_75t_L g817 ( .A1(n_792), .A2(n_818), .A3(n_821), .B1(n_824), .B2(n_827), .Y(n_817) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx2_ASAP7_75t_L g846 ( .A(n_794), .Y(n_846) );
INVx2_ASAP7_75t_L g897 ( .A(n_794), .Y(n_897) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVxp33_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND4xp25_ASAP7_75t_L g801 ( .A(n_802), .B(n_829), .C(n_858), .D(n_882), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_817), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_807), .Y(n_803) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g902 ( .A(n_810), .Y(n_902) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OR2x2_ASAP7_75t_L g875 ( .A(n_814), .B(n_850), .Y(n_875) );
INVx3_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_819), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g896 ( .A(n_820), .Y(n_896) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AOI311xp33_ASAP7_75t_L g882 ( .A1(n_822), .A2(n_883), .A3(n_884), .B(n_887), .C(n_898), .Y(n_882) );
BUFx3_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_838), .C(n_852), .Y(n_829) );
AOI31xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .A3(n_834), .B(n_836), .Y(n_830) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_842), .B1(n_845), .B2(n_848), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g862 ( .A(n_840), .Y(n_862) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OR2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g873 ( .A(n_847), .Y(n_873) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
AND2x4_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
AND2x2_ASAP7_75t_L g854 ( .A(n_850), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g861 ( .A(n_850), .Y(n_861) );
INVxp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
AOI211xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_863), .B(n_866), .C(n_874), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_860), .B(n_862), .Y(n_859) );
INVxp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
AOI21xp33_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B(n_880), .Y(n_874) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
AND2x4_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
INVx1_ASAP7_75t_L g888 ( .A(n_879), .Y(n_888) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_892), .B2(n_895), .Y(n_887) );
INVx2_ASAP7_75t_SL g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
OR2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_905), .A2(n_933), .B1(n_934), .B2(n_935), .Y(n_932) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_905), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_911), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_908), .B(n_911), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_911), .B(n_931), .Y(n_930) );
INVx8_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
OR2x6_ASAP7_75t_L g919 ( .A(n_912), .B(n_920), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
INVx2_ASAP7_75t_R g916 ( .A(n_917), .Y(n_916) );
BUFx3_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B(n_941), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_932), .Y(n_926) );
BUFx4f_ASAP7_75t_SL g927 ( .A(n_928), .Y(n_927) );
BUFx12f_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
BUFx8_ASAP7_75t_SL g943 ( .A(n_929), .Y(n_943) );
BUFx6f_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_940), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g940 ( .A(n_938), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
BUFx3_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
BUFx4_ASAP7_75t_SL g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g956 ( .A(n_948), .Y(n_956) );
OR2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_955), .Y(n_954) );
BUFx4_ASAP7_75t_SL g955 ( .A(n_956), .Y(n_955) );
endmodule