module fake_aes_7674_n_722 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_722);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_722;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_65), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_35), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_16), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_52), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_76), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_63), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_19), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_68), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_79), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_32), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_60), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_62), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_29), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_21), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_0), .Y(n_98) );
NOR2xp33_ASAP7_75t_L g99 ( .A(n_50), .B(n_22), .Y(n_99) );
NOR2xp33_ASAP7_75t_L g100 ( .A(n_64), .B(n_33), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_55), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_5), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_49), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_45), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_15), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_34), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_56), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_37), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_7), .B(n_36), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_1), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_10), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_4), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_24), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_17), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_18), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_15), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_6), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_51), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_9), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_109), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_129), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_119), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_82), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_90), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_126), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_102), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_121), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_111), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_113), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_80), .B(n_38), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_123), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_103), .B(n_2), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_80), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_114), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_105), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_105), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_108), .B(n_4), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_84), .B(n_5), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_108), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_87), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_88), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_88), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_89), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_89), .B(n_6), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_116), .B(n_7), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_128), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_81), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_116), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_120), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_92), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_131), .B(n_91), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_130), .B(n_107), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_157), .B(n_127), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_165), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_165), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_146), .B(n_101), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_157), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_130), .B(n_85), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_155), .B(n_97), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_170), .B(n_104), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_155), .B(n_104), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_156), .B(n_110), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_165), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_171), .B(n_127), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_140), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_158), .A2(n_110), .B1(n_93), .B2(n_96), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_171), .B(n_124), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_158), .B(n_120), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_166), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_137), .B(n_92), .Y(n_210) );
AND2x6_ASAP7_75t_L g211 ( .A(n_158), .B(n_115), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_143), .B(n_93), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_149), .B(n_124), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_147), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_148), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
NOR2xp33_ASAP7_75t_SL g218 ( .A(n_147), .B(n_115), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_147), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_148), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_134), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_134), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
INVxp67_ASAP7_75t_L g226 ( .A(n_145), .Y(n_226) );
INVx6_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_147), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_139), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_147), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_138), .B(n_118), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_147), .Y(n_232) );
OAI221xp5_ASAP7_75t_L g233 ( .A1(n_152), .A2(n_122), .B1(n_125), .B2(n_98), .C(n_94), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_168), .B(n_122), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_168), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_142), .B(n_112), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_142), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_162), .B(n_118), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_174), .B(n_173), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_236), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_179), .B(n_172), .Y(n_244) );
NOR2xp33_ASAP7_75t_R g245 ( .A(n_218), .B(n_132), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_228), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_239), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_226), .B(n_133), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_217), .Y(n_250) );
O2A1O1Ixp5_ASAP7_75t_L g251 ( .A1(n_195), .A2(n_167), .B(n_159), .C(n_163), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_239), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_236), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_194), .B(n_173), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_195), .B(n_152), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_203), .B(n_142), .Y(n_256) );
AND2x6_ASAP7_75t_L g257 ( .A(n_228), .B(n_112), .Y(n_257) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_186), .A2(n_163), .B(n_153), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_236), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_195), .B(n_153), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_233), .B(n_169), .C(n_154), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_181), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_239), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_236), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_223), .Y(n_267) );
NOR3xp33_ASAP7_75t_SL g268 ( .A(n_182), .B(n_169), .C(n_154), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_194), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_180), .B(n_150), .Y(n_271) );
BUFx4f_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_209), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_194), .B(n_164), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_223), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_228), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_194), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_187), .B(n_164), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_185), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_215), .B(n_96), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_237), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_224), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_176), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_211), .A2(n_161), .B1(n_160), .B2(n_151), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_235), .B(n_161), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_189), .B(n_160), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_211), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g290 ( .A1(n_200), .A2(n_145), .B1(n_135), .B2(n_151), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_215), .B(n_141), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_176), .B(n_141), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_238), .Y(n_293) );
AND3x1_ASAP7_75t_SL g294 ( .A(n_201), .B(n_8), .C(n_10), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_237), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_200), .B(n_99), .Y(n_297) );
NOR2xp33_ASAP7_75t_R g298 ( .A(n_211), .B(n_215), .Y(n_298) );
BUFx4_ASAP7_75t_SL g299 ( .A(n_183), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_219), .A2(n_95), .B(n_100), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_237), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_228), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_230), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_213), .B(n_8), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_177), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_201), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_177), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_175), .B(n_11), .C(n_12), .Y(n_309) );
AND3x1_ASAP7_75t_SL g310 ( .A(n_200), .B(n_11), .C(n_13), .Y(n_310) );
AND3x1_ASAP7_75t_SL g311 ( .A(n_200), .B(n_14), .C(n_17), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_SL g312 ( .A1(n_178), .A2(n_44), .B(n_77), .C(n_75), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_254), .B(n_211), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_262), .B(n_234), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_277), .A2(n_211), .B1(n_227), .B2(n_235), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
AOI21x1_ASAP7_75t_L g317 ( .A1(n_275), .A2(n_191), .B(n_192), .Y(n_317) );
NAND2xp33_ASAP7_75t_L g318 ( .A(n_298), .B(n_230), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_270), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_271), .A2(n_227), .B1(n_234), .B2(n_206), .Y(n_320) );
BUFx4f_ASAP7_75t_L g321 ( .A(n_257), .Y(n_321) );
NOR2x1p5_ASAP7_75t_SL g322 ( .A(n_243), .B(n_188), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_246), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_271), .B(n_238), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_262), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_253), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_291), .A2(n_232), .B(n_219), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_281), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_227), .B1(n_234), .B2(n_206), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_284), .B(n_214), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_273), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_272), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_272), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_247), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_273), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_253), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_259), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_259), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_297), .B(n_227), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_263), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_264), .B(n_206), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_250), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_307), .B(n_214), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_247), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_298), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_291), .A2(n_232), .B(n_219), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_247), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_241), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_297), .A2(n_235), .B1(n_234), .B2(n_206), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_263), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_255), .A2(n_232), .B(n_230), .Y(n_356) );
INVx5_ASAP7_75t_SL g357 ( .A(n_247), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_269), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_274), .B(n_238), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_289), .Y(n_360) );
INVxp33_ASAP7_75t_L g361 ( .A(n_244), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_285), .A2(n_196), .B1(n_202), .B2(n_240), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_289), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_266), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_255), .A2(n_230), .B(n_231), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_285), .A2(n_196), .B1(n_202), .B2(n_230), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_299), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_316), .A2(n_251), .B(n_286), .C(n_309), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_367), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_314), .B(n_241), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_331), .A2(n_290), .B1(n_279), .B2(n_249), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_361), .B(n_242), .Y(n_373) );
OAI21xp33_ASAP7_75t_SL g374 ( .A1(n_341), .A2(n_331), .B(n_354), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_337), .A2(n_249), .B1(n_292), .B2(n_288), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_346), .B(n_278), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_323), .B(n_249), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_341), .A2(n_245), .B1(n_258), .B2(n_305), .Y(n_381) );
OA21x2_ASAP7_75t_L g382 ( .A1(n_317), .A2(n_301), .B(n_220), .Y(n_382) );
INVx4_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_324), .B(n_256), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_314), .B(n_248), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_316), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_337), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_324), .B(n_261), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_341), .A2(n_245), .B1(n_258), .B2(n_286), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_367), .Y(n_390) );
BUFx4f_ASAP7_75t_L g391 ( .A(n_341), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_345), .A2(n_252), .B1(n_265), .B2(n_280), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_330), .A2(n_268), .B1(n_210), .B2(n_229), .C(n_225), .Y(n_393) );
AND2x6_ASAP7_75t_L g394 ( .A(n_314), .B(n_269), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_314), .B(n_260), .Y(n_395) );
NAND2x1_ASAP7_75t_L g396 ( .A(n_352), .B(n_257), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_320), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_326), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_320), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_327), .A2(n_343), .B1(n_321), .B2(n_360), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_343), .Y(n_401) );
INVxp33_ASAP7_75t_L g402 ( .A(n_370), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_SL g403 ( .A1(n_384), .A2(n_352), .B(n_204), .C(n_197), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_399), .A2(n_344), .B1(n_330), .B2(n_359), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_378), .B(n_344), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_399), .A2(n_359), .B1(n_343), .B2(n_313), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_391), .A2(n_313), .B1(n_343), .B2(n_321), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_401), .B(n_350), .Y(n_409) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_376), .A2(n_353), .B1(n_350), .B2(n_315), .C1(n_294), .C2(n_319), .Y(n_410) );
OAI22xp5_ASAP7_75t_SL g411 ( .A1(n_372), .A2(n_311), .B1(n_310), .B2(n_353), .Y(n_411) );
INVx2_ASAP7_75t_SL g412 ( .A(n_391), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g414 ( .A1(n_377), .A2(n_363), .B1(n_360), .B2(n_321), .C1(n_362), .C2(n_327), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_397), .A2(n_321), .B1(n_363), .B2(n_348), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_379), .B(n_225), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_368), .A2(n_318), .B(n_356), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g419 ( .A1(n_373), .A2(n_280), .B1(n_366), .B2(n_334), .C1(n_229), .C2(n_257), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_374), .B(n_352), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_387), .A2(n_348), .B1(n_334), .B2(n_325), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_394), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_375), .A2(n_352), .B1(n_257), .B2(n_325), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_368), .A2(n_356), .B(n_365), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_373), .B(n_326), .Y(n_425) );
OAI21x1_ASAP7_75t_L g426 ( .A1(n_382), .A2(n_317), .B(n_365), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_257), .B1(n_334), .B2(n_335), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_394), .Y(n_428) );
BUFx8_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_404), .A2(n_383), .B1(n_384), .B2(n_380), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_417), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_425), .Y(n_433) );
BUFx12f_ASAP7_75t_L g434 ( .A(n_429), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_420), .B(n_383), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_383), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_406), .B(n_381), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_430), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_429), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_425), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_410), .B(n_393), .C(n_389), .D(n_392), .Y(n_441) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_410), .A2(n_390), .B(n_369), .C(n_400), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_411), .A2(n_395), .B1(n_385), .B2(n_371), .Y(n_444) );
NOR4xp25_ASAP7_75t_SL g445 ( .A(n_405), .B(n_312), .C(n_390), .D(n_396), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_411), .A2(n_395), .B1(n_385), .B2(n_371), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_426), .A2(n_220), .B(n_193), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_404), .A2(n_385), .B1(n_395), .B2(n_312), .C(n_212), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_402), .B(n_335), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_405), .A2(n_207), .B1(n_212), .B2(n_205), .C(n_199), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_423), .A2(n_382), .B(n_205), .C(n_207), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_420), .B(n_382), .Y(n_452) );
NAND2xp33_ASAP7_75t_SL g453 ( .A(n_412), .B(n_334), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_409), .B(n_394), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_416), .B(n_394), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_407), .A2(n_302), .B1(n_266), .B2(n_282), .Y(n_456) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_424), .A2(n_193), .B(n_222), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_413), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_419), .B(n_208), .C(n_199), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_413), .B(n_322), .Y(n_461) );
AOI33xp33_ASAP7_75t_L g462 ( .A1(n_416), .A2(n_198), .A3(n_178), .B1(n_190), .B2(n_191), .B3(n_192), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_418), .A2(n_216), .B(n_204), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_409), .B(n_339), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_414), .B(n_322), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g467 ( .A1(n_414), .A2(n_364), .B(n_355), .Y(n_467) );
AOI211xp5_ASAP7_75t_L g468 ( .A1(n_442), .A2(n_415), .B(n_421), .C(n_408), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_443), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_435), .B(n_422), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_433), .B(n_422), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_458), .B(n_428), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_440), .B(n_412), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_458), .B(n_428), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_459), .B(n_14), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_465), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_437), .B(n_408), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_437), .B(n_18), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_434), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_434), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_438), .B(n_427), .C(n_429), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_431), .B(n_429), .C(n_419), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_452), .B(n_19), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_436), .B(n_403), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_459), .B(n_20), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_436), .B(n_20), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_449), .B(n_208), .C(n_198), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_441), .B(n_208), .C(n_190), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_465), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_439), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_444), .B(n_364), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_364), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_435), .B(n_326), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_441), .A2(n_300), .A3(n_287), .B(n_302), .Y(n_498) );
OAI31xp33_ASAP7_75t_L g499 ( .A1(n_446), .A2(n_300), .A3(n_287), .B(n_282), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_435), .B(n_328), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_439), .B(n_328), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_461), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_454), .B(n_328), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_448), .B(n_208), .C(n_184), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_461), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_452), .B(n_338), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_461), .B(n_338), .Y(n_508) );
OR2x6_ASAP7_75t_SL g509 ( .A(n_466), .B(n_338), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
OR2x6_ASAP7_75t_L g511 ( .A(n_466), .B(n_358), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_455), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
NOR2xp33_ASAP7_75t_SL g516 ( .A(n_467), .B(n_358), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_467), .B(n_355), .Y(n_517) );
OAI31xp33_ASAP7_75t_L g518 ( .A1(n_453), .A2(n_295), .A3(n_260), .B(n_355), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_462), .B(n_208), .C(n_222), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_456), .B(n_342), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_469), .B(n_457), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_503), .B(n_457), .Y(n_522) );
NOR4xp25_ASAP7_75t_SL g523 ( .A(n_474), .B(n_445), .C(n_450), .D(n_460), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_479), .B(n_457), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_492), .B(n_457), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_503), .B(n_464), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_506), .B(n_464), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_513), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_480), .B(n_464), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_483), .B(n_25), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_485), .B(n_460), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_506), .B(n_464), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_483), .B(n_26), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_471), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_475), .B(n_451), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_486), .Y(n_536) );
INVx3_ASAP7_75t_SL g537 ( .A(n_474), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_486), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_510), .B(n_447), .Y(n_539) );
AND4x1_ASAP7_75t_L g540 ( .A(n_468), .B(n_445), .C(n_28), .D(n_30), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_502), .B(n_447), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_482), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_478), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_510), .B(n_447), .Y(n_544) );
OR2x6_ASAP7_75t_L g545 ( .A(n_511), .B(n_447), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_514), .B(n_339), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_507), .B(n_197), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_507), .B(n_188), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_516), .B(n_357), .Y(n_549) );
OAI21xp33_ASAP7_75t_L g550 ( .A1(n_487), .A2(n_216), .B(n_221), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_481), .B(n_342), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_508), .B(n_184), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_508), .B(n_221), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_480), .B(n_342), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_493), .B(n_27), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_488), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_511), .B(n_39), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_476), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_472), .B(n_339), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_511), .B(n_40), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_472), .Y(n_561) );
NAND2xp33_ASAP7_75t_SL g562 ( .A(n_509), .B(n_340), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_473), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_481), .B(n_340), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_494), .B(n_340), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_473), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_511), .B(n_41), .Y(n_567) );
AOI33xp33_ASAP7_75t_L g568 ( .A1(n_477), .A2(n_295), .A3(n_306), .B1(n_308), .B2(n_48), .B3(n_54), .Y(n_568) );
BUFx2_ASAP7_75t_SL g569 ( .A(n_482), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_512), .B(n_357), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_509), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_501), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_477), .B(n_42), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_496), .B(n_358), .Y(n_575) );
INVx4_ASAP7_75t_L g576 ( .A(n_470), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_497), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_489), .B(n_357), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_512), .B(n_357), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_534), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_574), .B(n_497), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_571), .A2(n_484), .B1(n_470), .B2(n_500), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_569), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_536), .A2(n_491), .B1(n_495), .B2(n_504), .C(n_505), .Y(n_584) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_531), .A2(n_498), .B(n_490), .Y(n_585) );
AND2x4_ASAP7_75t_SL g586 ( .A(n_576), .B(n_500), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_577), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_558), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_531), .A2(n_515), .B(n_520), .Y(n_589) );
INVx3_ASAP7_75t_L g590 ( .A(n_576), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g591 ( .A1(n_538), .A2(n_470), .B1(n_515), .B2(n_517), .C1(n_513), .C2(n_519), .Y(n_591) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_537), .A2(n_499), .B(n_518), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_572), .B(n_43), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_521), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_521), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_576), .A2(n_336), .B1(n_351), .B2(n_347), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_537), .A2(n_329), .B(n_349), .C(n_336), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_563), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_529), .B(n_47), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_529), .B(n_59), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_542), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_559), .Y(n_603) );
OAI32xp33_ASAP7_75t_L g604 ( .A1(n_562), .A2(n_347), .A3(n_351), .B1(n_67), .B2(n_69), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_562), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_568), .A2(n_329), .B(n_349), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_566), .B(n_61), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_557), .A2(n_357), .B1(n_351), .B2(n_347), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_556), .B(n_66), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_524), .B(n_70), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_557), .A2(n_308), .B1(n_306), .B2(n_78), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_530), .B(n_72), .C(n_73), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_543), .B(n_269), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_535), .A2(n_269), .B1(n_276), .B2(n_303), .C(n_304), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_528), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
OA21x2_ASAP7_75t_L g617 ( .A1(n_525), .A2(n_276), .B(n_303), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_533), .B(n_276), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_541), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_528), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_578), .B(n_276), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_539), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_565), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_546), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_522), .Y(n_625) );
XNOR2x2_ASAP7_75t_L g626 ( .A(n_560), .B(n_303), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_522), .B(n_303), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_526), .B(n_527), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_526), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_568), .B(n_304), .C(n_540), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_527), .B(n_304), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_620), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_602), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_588), .A2(n_551), .B1(n_564), .B2(n_532), .C(n_573), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_580), .Y(n_635) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_583), .B(n_590), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_604), .A2(n_549), .B(n_545), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_581), .B(n_545), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_582), .A2(n_567), .B1(n_545), .B2(n_553), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_586), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_603), .B(n_575), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_619), .B(n_539), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_595), .B(n_544), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_628), .B(n_545), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_596), .B(n_544), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_599), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_593), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_587), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_628), .B(n_579), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_623), .B(n_547), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_616), .B(n_579), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_622), .B(n_553), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_594), .B(n_570), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_624), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_625), .B(n_552), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_629), .B(n_547), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_608), .B(n_575), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_585), .A2(n_549), .B(n_605), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_592), .B(n_570), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_591), .B(n_548), .Y(n_660) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_626), .B(n_555), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_590), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_607), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_615), .B(n_552), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_600), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_600), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_640), .B(n_589), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_659), .A2(n_585), .B1(n_612), .B2(n_584), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_640), .B(n_611), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_659), .A2(n_601), .B1(n_609), .B2(n_610), .C1(n_630), .C2(n_606), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_639), .A2(n_601), .B1(n_610), .B2(n_631), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_636), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_637), .A2(n_597), .B(n_618), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_633), .Y(n_675) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_664), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_664), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_661), .B(n_614), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_664), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_660), .A2(n_621), .B1(n_548), .B2(n_627), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_635), .Y(n_681) );
O2A1O1Ixp5_ASAP7_75t_SL g682 ( .A1(n_647), .A2(n_613), .B(n_523), .C(n_598), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_646), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_648), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_654), .A2(n_555), .B1(n_550), .B2(n_617), .C(n_304), .Y(n_685) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_658), .A2(n_617), .B(n_657), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_644), .B(n_638), .Y(n_687) );
INVxp33_ASAP7_75t_L g688 ( .A(n_661), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_688), .A2(n_663), .B1(n_662), .B2(n_641), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_675), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_686), .A2(n_634), .B(n_666), .C(n_665), .Y(n_691) );
BUFx2_ASAP7_75t_L g692 ( .A(n_676), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_681), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_680), .B(n_655), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_683), .Y(n_695) );
AOI21xp33_ASAP7_75t_SL g696 ( .A1(n_688), .A2(n_653), .B(n_651), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_684), .B(n_678), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_679), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_677), .B(n_651), .Y(n_699) );
NAND4xp25_ASAP7_75t_SL g700 ( .A(n_668), .B(n_649), .C(n_642), .D(n_650), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_674), .A2(n_653), .B(n_656), .C(n_645), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_667), .A2(n_652), .B1(n_643), .B2(n_632), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_673), .A2(n_669), .B1(n_687), .B2(n_671), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_673), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_672), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_682), .B(n_670), .C(n_669), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_685), .B(n_672), .C(n_687), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_682), .A2(n_688), .B(n_686), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_690), .Y(n_709) );
INVx1_ASAP7_75t_SL g710 ( .A(n_692), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_689), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_703), .Y(n_712) );
AOI21x1_ASAP7_75t_L g713 ( .A1(n_704), .A2(n_706), .B(n_697), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_710), .B(n_708), .C(n_691), .D(n_696), .Y(n_714) );
AOI221xp5_ASAP7_75t_SL g715 ( .A1(n_712), .A2(n_694), .B1(n_699), .B2(n_705), .C(n_691), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_711), .A2(n_700), .B1(n_707), .B2(n_698), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_714), .A2(n_709), .B(n_701), .Y(n_717) );
BUFx8_ASAP7_75t_L g718 ( .A(n_715), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_717), .B(n_716), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
AOI22xp5_ASAP7_75t_SL g721 ( .A1(n_720), .A2(n_709), .B1(n_713), .B2(n_693), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_719), .B1(n_702), .B2(n_695), .C(n_705), .Y(n_722) );
endmodule