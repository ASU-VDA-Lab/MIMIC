module fake_jpeg_621_n_62 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_62);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_25),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_21),
.C(n_20),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_2),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_4),
.B(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_56),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_51),
.B1(n_57),
.B2(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_50),
.Y(n_62)
);


endmodule