module fake_jpeg_14592_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_3),
.B(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_38),
.B(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_32),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_48),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_10),
.B(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_63),
.B1(n_7),
.B2(n_8),
.Y(n_97)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_24),
.B1(n_21),
.B2(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_37),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_20),
.B(n_13),
.Y(n_121)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_82),
.Y(n_106)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_25),
.B1(n_33),
.B2(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_63),
.B1(n_20),
.B2(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_35),
.B1(n_33),
.B2(n_29),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_90),
.B1(n_92),
.B2(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_102),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_42),
.A2(n_22),
.B1(n_27),
.B2(n_35),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_27),
.B1(n_26),
.B2(n_31),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_26),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_100),
.B(n_65),
.C(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_41),
.B(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_44),
.B(n_31),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_117),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_129),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_10),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_114),
.B1(n_129),
.B2(n_127),
.Y(n_143)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_125),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_30),
.B1(n_20),
.B2(n_28),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_121),
.B(n_87),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_20),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_123),
.C(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_124),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_30),
.B(n_28),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_12),
.B1(n_14),
.B2(n_81),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_126),
.A2(n_76),
.B1(n_87),
.B2(n_77),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_130),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_70),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_64),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_134),
.B1(n_124),
.B2(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_138),
.B(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_109),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_156),
.B(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_151),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_71),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_148),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_79),
.B1(n_72),
.B2(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_160),
.B1(n_137),
.B2(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_98),
.B(n_77),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_69),
.C(n_71),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_135),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_69),
.B(n_106),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_174),
.C(n_180),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_179),
.B(n_183),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_161),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_103),
.B1(n_111),
.B2(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_111),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_183),
.B(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_177),
.B1(n_136),
.B2(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_145),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_146),
.B1(n_143),
.B2(n_148),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_162),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_153),
.B(n_151),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_184),
.Y(n_187)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_185),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_159),
.C(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_171),
.C(n_173),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_177),
.B1(n_166),
.B2(n_165),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_199),
.B1(n_170),
.B2(n_184),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_175),
.B1(n_179),
.B2(n_178),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_205),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_182),
.C(n_164),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_214),
.B(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_195),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_213),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_189),
.B(n_200),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_218),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_204),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_221),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_216),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_205),
.C(n_203),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_194),
.C(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_209),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_234),
.B(n_225),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_229),
.B1(n_226),
.B2(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_194),
.C(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_237),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_232),
.C(n_207),
.Y(n_238)
);

AOI211xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_239),
.B(n_207),
.C(n_201),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_198),
.Y(n_241)
);


endmodule