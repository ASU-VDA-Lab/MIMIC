module fake_jpeg_20582_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_55),
.B1(n_75),
.B2(n_74),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_54),
.B1(n_72),
.B2(n_76),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_76),
.B1(n_73),
.B2(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_85),
.Y(n_99)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_78),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_73),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_60),
.B1(n_77),
.B2(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_96),
.B1(n_93),
.B2(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_118),
.B1(n_59),
.B2(n_65),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_70),
.B1(n_77),
.B2(n_68),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_69),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_0),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_108),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_139),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_117),
.B1(n_118),
.B2(n_3),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_58),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_136),
.B(n_21),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_19),
.B(n_49),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_144),
.B1(n_4),
.B2(n_6),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_27),
.C(n_48),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_12),
.C(n_14),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_1),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_148),
.B(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_155),
.B1(n_140),
.B2(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_152),
.B(n_151),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_160),
.B1(n_153),
.B2(n_158),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_142),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_156),
.C(n_29),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_16),
.B(n_32),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_37),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_167),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_39),
.B(n_40),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_46),
.CI(n_47),
.CON(n_171),
.SN(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_50),
.Y(n_172)
);


endmodule