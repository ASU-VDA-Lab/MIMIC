module fake_jpeg_5562_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_39),
.B1(n_29),
.B2(n_37),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_50),
.B1(n_54),
.B2(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_27),
.B1(n_30),
.B2(n_23),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_30),
.B1(n_15),
.B2(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_22),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_21),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_74),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_35),
.B(n_17),
.C(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

CKINVDCx11_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_51),
.B1(n_48),
.B2(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_44),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_53),
.C(n_56),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_91),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_57),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_66),
.B(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_43),
.C(n_44),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_81),
.B1(n_77),
.B2(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_63),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_68),
.B1(n_71),
.B2(n_64),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_97),
.B(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_118),
.C(n_86),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_64),
.B(n_74),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_100),
.B(n_92),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_116),
.B(n_28),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_119),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_68),
.B(n_76),
.C(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_120),
.B1(n_111),
.B2(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_100),
.B(n_93),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_65),
.B1(n_67),
.B2(n_52),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_31),
.B1(n_37),
.B2(n_32),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_98),
.B1(n_90),
.B2(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_124),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_65),
.B1(n_32),
.B2(n_37),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_135),
.B1(n_139),
.B2(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_132),
.C(n_133),
.Y(n_157)
);

NOR4xp25_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_85),
.C(n_92),
.D(n_87),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_130),
.B(n_1),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_101),
.A3(n_86),
.B1(n_44),
.B2(n_104),
.C1(n_13),
.C2(n_14),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_138),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_38),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_117),
.C(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_124),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_32),
.B(n_31),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_88),
.B1(n_31),
.B2(n_28),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_0),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_38),
.B(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_134),
.A2(n_119),
.B1(n_122),
.B2(n_110),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_150),
.B(n_126),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_117),
.B1(n_112),
.B2(n_105),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_151),
.B1(n_155),
.B2(n_2),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_88),
.B1(n_80),
.B2(n_38),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_154),
.Y(n_159)
);

OA21x2_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_3),
.B(n_4),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_80),
.B1(n_14),
.B2(n_13),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_133),
.C(n_132),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_144),
.C(n_145),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_130),
.B1(n_141),
.B2(n_140),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_167),
.B1(n_5),
.B2(n_6),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_130),
.B(n_142),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_164),
.B(n_169),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_3),
.B(n_4),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_175),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_178),
.B(n_170),
.Y(n_184)
);

AOI31xp67_ASAP7_75t_L g175 ( 
.A1(n_164),
.A2(n_150),
.A3(n_148),
.B(n_154),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_151),
.C(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_5),
.C(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_167),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_185),
.B1(n_174),
.B2(n_7),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_7),
.B(n_9),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_165),
.B(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_159),
.B1(n_161),
.B2(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_177),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_190),
.C(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_188),
.B(n_6),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_7),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_189),
.C(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

OAI31xp33_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_198),
.A3(n_195),
.B(n_10),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_202),
.Y(n_204)
);


endmodule