module fake_netlist_5_1852_n_2880 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_520, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2880);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_520;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2880;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_549;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_1462;
wire n_1799;
wire n_854;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_2538;
wire n_2105;
wire n_877;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_556;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_976;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_553;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_1880;
wire n_888;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_571;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_586;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_931;
wire n_1711;
wire n_599;
wire n_1891;
wire n_1662;
wire n_870;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_1798;
wire n_2022;
wire n_776;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_1539;
wire n_946;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_2029;
wire n_742;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_2565;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2111;
wire n_1724;
wire n_2521;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_701;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_1954;
wire n_802;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1735;
wire n_1697;
wire n_1575;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_555;
wire n_1848;
wire n_1928;
wire n_783;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_693;
wire n_1506;
wire n_2653;
wire n_990;
wire n_836;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_2259;
wire n_1702;
wire n_2794;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_1499;
wire n_711;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1929;
wire n_1597;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2201;
wire n_1737;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1584;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1944;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_2695;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_927;
wire n_2044;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g543 ( 
.A(n_387),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_192),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_347),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_409),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_354),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_215),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

BUFx2_ASAP7_75t_SL g550 ( 
.A(n_355),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_382),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_393),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_135),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_536),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_248),
.Y(n_555)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_399),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_242),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_222),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_335),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_209),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_356),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_414),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_425),
.Y(n_565)
);

BUFx2_ASAP7_75t_SL g566 ( 
.A(n_172),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_231),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_496),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_348),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_442),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_483),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_405),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_348),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_498),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_527),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_115),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_80),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_495),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_280),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_80),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_10),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

BUFx8_ASAP7_75t_SL g583 ( 
.A(n_388),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_219),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_532),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_39),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_47),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_166),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_424),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_469),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_406),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_8),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_342),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_266),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_195),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_113),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_141),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_473),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_518),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_380),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_205),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_169),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_481),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_266),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_365),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_354),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_366),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_476),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_415),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_283),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_511),
.Y(n_612)
);

BUFx5_ASAP7_75t_L g613 ( 
.A(n_140),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_450),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_18),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_91),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_308),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_402),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_360),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_195),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_48),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_500),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_513),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_504),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_419),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_421),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_82),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_398),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_262),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_519),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_332),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_203),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_412),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_535),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_1),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_13),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_458),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_358),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_123),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_127),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_292),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_378),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_221),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_124),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_86),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_368),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_140),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_411),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_106),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_515),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_60),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_149),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_147),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_155),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_205),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_115),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_29),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_523),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_391),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_457),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_462),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_238),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_355),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_350),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_141),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_522),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_497),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_256),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_171),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_232),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_209),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_318),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_1),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_100),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_88),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_338),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_153),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_418),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_318),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_390),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_430),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_252),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_403),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_329),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_220),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_365),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_485),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_489),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_539),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_445),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_246),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_427),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_507),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_294),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_3),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_240),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_53),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_372),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_130),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_128),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_509),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_410),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_103),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_317),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_358),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_506),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_186),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_499),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_392),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_344),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_400),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_337),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_512),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_38),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_433),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_49),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_431),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_219),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_192),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_323),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_101),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_163),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_437),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_203),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_438),
.Y(n_725)
);

BUFx2_ASAP7_75t_SL g726 ( 
.A(n_171),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_143),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_467),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_475),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_276),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_413),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_163),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_542),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_103),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_31),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_196),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_304),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_102),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_460),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_517),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_516),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_137),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_81),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_213),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_164),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_164),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_494),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_230),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_363),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_102),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_108),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_490),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_301),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_101),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_119),
.Y(n_755)
);

BUFx5_ASAP7_75t_L g756 ( 
.A(n_484),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_172),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_453),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_72),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_528),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_155),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_23),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_277),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_471),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_357),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_379),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_477),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_43),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_255),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_389),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_131),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_263),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_465),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_320),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_149),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_144),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_370),
.Y(n_777)
);

BUFx10_ASAP7_75t_L g778 ( 
.A(n_56),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_311),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_315),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_385),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_530),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_531),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_503),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_441),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_466),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_429),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_346),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_456),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_76),
.Y(n_790)
);

INVxp33_ASAP7_75t_R g791 ( 
.A(n_492),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_451),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_367),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_446),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_435),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_284),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_534),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_158),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_327),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_486),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_181),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_18),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_243),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_329),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_146),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_51),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_151),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_182),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_533),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_62),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_459),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_36),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_375),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_92),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_353),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_224),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_468),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_255),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_260),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_434),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_397),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_525),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_463),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_488),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_323),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_386),
.Y(n_826)
);

CKINVDCx14_ASAP7_75t_R g827 ( 
.A(n_452),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_383),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_50),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_298),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_420),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_330),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_35),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_207),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_364),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_444),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_464),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_461),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_284),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_123),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_396),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_24),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_432),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_5),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_253),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_394),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_491),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_278),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_114),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_24),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_166),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_361),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_374),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_296),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_423),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_27),
.Y(n_856)
);

BUFx10_ASAP7_75t_L g857 ( 
.A(n_67),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_98),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_493),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_119),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_455),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_331),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_362),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_142),
.Y(n_864)
);

BUFx8_ASAP7_75t_SL g865 ( 
.A(n_39),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_114),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_336),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_9),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_188),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_36),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_56),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_44),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_147),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_520),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_356),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_487),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_474),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_367),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_440),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_373),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_334),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_302),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_259),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_121),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_90),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_479),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_154),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_529),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_514),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_66),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_23),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_447),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_401),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_28),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_395),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_537),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_324),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_65),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_48),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_480),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_117),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_185),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_94),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_254),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_252),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_349),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_482),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_120),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_230),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_87),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_408),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_297),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_454),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_281),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_508),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_505),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_247),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_524),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_42),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_250),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_422),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_381),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_448),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_241),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_502),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_352),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_59),
.Y(n_927)
);

BUFx8_ASAP7_75t_SL g928 ( 
.A(n_137),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_521),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_211),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_384),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_38),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_229),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_72),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_204),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_262),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_526),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_470),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_282),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_105),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_212),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_112),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_215),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_334),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_478),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_144),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_404),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_416),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_52),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_303),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_449),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_472),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_201),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_407),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_63),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_359),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_217),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_207),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_237),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_351),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_436),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_201),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_60),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_540),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_538),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_541),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_353),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_132),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_319),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_35),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_337),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_210),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_417),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_234),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_288),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_70),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_510),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_100),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_73),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_235),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_613),
.Y(n_981)
);

CKINVDCx16_ASAP7_75t_R g982 ( 
.A(n_647),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_613),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_613),
.Y(n_984)
);

INVxp33_ASAP7_75t_L g985 ( 
.A(n_757),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_641),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_939),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_865),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_716),
.Y(n_989)
);

INVxp33_ASAP7_75t_L g990 ( 
.A(n_738),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_582),
.Y(n_991)
);

INVxp33_ASAP7_75t_SL g992 ( 
.A(n_544),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_928),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_613),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_613),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_613),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_758),
.B(n_0),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_953),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_613),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_613),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_602),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_581),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_602),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_705),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_705),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_615),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_812),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_812),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_SL g1009 ( 
.A(n_708),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_801),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_829),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_581),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_829),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_926),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_926),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_619),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_830),
.Y(n_1017)
);

INVxp67_ASAP7_75t_SL g1018 ( 
.A(n_688),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_941),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_941),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_581),
.Y(n_1021)
);

INVxp33_ASAP7_75t_SL g1022 ( 
.A(n_544),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_636),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_581),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_597),
.Y(n_1025)
);

INVxp33_ASAP7_75t_SL g1026 ( 
.A(n_545),
.Y(n_1026)
);

CKINVDCx16_ASAP7_75t_R g1027 ( 
.A(n_599),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_581),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_670),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_616),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_670),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_794),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_640),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_652),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_670),
.Y(n_1035)
);

INVxp33_ASAP7_75t_SL g1036 ( 
.A(n_545),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_703),
.Y(n_1037)
);

INVxp67_ASAP7_75t_SL g1038 ( 
.A(n_795),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_670),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_925),
.Y(n_1040)
);

CKINVDCx16_ASAP7_75t_R g1041 ( 
.A(n_827),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_620),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_759),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_759),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_759),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_759),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_759),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_890),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_727),
.Y(n_1049)
);

INVxp67_ASAP7_75t_SL g1050 ( 
.A(n_582),
.Y(n_1050)
);

INVxp67_ASAP7_75t_SL g1051 ( 
.A(n_660),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_890),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_890),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1053),
.Y(n_1054)
);

BUFx12f_ASAP7_75t_L g1055 ( 
.A(n_993),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_991),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_995),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1053),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_998),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_986),
.B(n_636),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_996),
.A2(n_585),
.B(n_571),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1032),
.B(n_556),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1002),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_996),
.A2(n_585),
.B(n_571),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1050),
.B(n_761),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1002),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1012),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1012),
.Y(n_1068)
);

OA21x2_ASAP7_75t_L g1069 ( 
.A1(n_981),
.A2(n_678),
.B(n_650),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_995),
.A2(n_678),
.B(n_650),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_983),
.A2(n_698),
.B(n_692),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1045),
.Y(n_1072)
);

XNOR2x2_ASAP7_75t_L g1073 ( 
.A(n_989),
.B(n_704),
.Y(n_1073)
);

CKINVDCx6p67_ASAP7_75t_R g1074 ( 
.A(n_1027),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1051),
.B(n_890),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1045),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_1025),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1025),
.A2(n_762),
.B1(n_806),
.B2(n_743),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_991),
.B(n_761),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1047),
.Y(n_1080)
);

OA22x2_ASAP7_75t_L g1081 ( 
.A1(n_1001),
.A2(n_819),
.B1(n_772),
.B2(n_654),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1021),
.B(n_846),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1047),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_984),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1003),
.B(n_772),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_1038),
.B(n_556),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1024),
.B(n_846),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_994),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_999),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1000),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1028),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1004),
.B(n_819),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1029),
.A2(n_698),
.B(n_692),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1031),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1035),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1039),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_1043),
.A2(n_859),
.B(n_549),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_997),
.A2(n_878),
.B1(n_899),
.B2(n_835),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1048),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_993),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1005),
.B(n_971),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_1041),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1052),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1007),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1008),
.B(n_660),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1011),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1013),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1014),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1015),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1019),
.Y(n_1111)
);

CKINVDCx6p67_ASAP7_75t_R g1112 ( 
.A(n_1040),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_998),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_1077),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1091),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1101),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_1074),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1055),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1055),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1055),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1091),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1108),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1091),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1074),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_1074),
.B(n_1006),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1112),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1108),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1062),
.B(n_992),
.Y(n_1128)
);

AOI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1075),
.A2(n_554),
.B(n_543),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1108),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1095),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1057),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1112),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1112),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1105),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1056),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1056),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1056),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1059),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1113),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1103),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1073),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1086),
.B(n_992),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_1103),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1089),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1103),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1103),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1106),
.B(n_709),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1103),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1057),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1103),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1103),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1065),
.B(n_1018),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1078),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1078),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_R g1156 ( 
.A(n_1065),
.B(n_1006),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1105),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1079),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1099),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_1088),
.B(n_1016),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1099),
.Y(n_1161)
);

XNOR2xp5_ASAP7_75t_L g1162 ( 
.A(n_1073),
.B(n_1030),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1107),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1079),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_1075),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1106),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1095),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1095),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1106),
.B(n_987),
.Y(n_1169)
);

BUFx10_ASAP7_75t_L g1170 ( 
.A(n_1106),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1057),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1128),
.B(n_1143),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1170),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1158),
.B(n_990),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1156),
.B(n_1088),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1135),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1145),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1157),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1122),
.B(n_1088),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1170),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1165),
.B(n_1022),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1170),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1169),
.B(n_1016),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1142),
.B(n_1081),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1145),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1115),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1163),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1127),
.B(n_1088),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1130),
.B(n_1090),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1148),
.B(n_1109),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1153),
.B(n_1090),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1145),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1114),
.Y(n_1194)
);

XOR2xp5_ASAP7_75t_L g1195 ( 
.A(n_1114),
.B(n_1030),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1162),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1139),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1148),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1148),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1132),
.Y(n_1200)
);

OAI22x1_ASAP7_75t_L g1201 ( 
.A1(n_1159),
.A2(n_1023),
.B1(n_1010),
.B2(n_1017),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1115),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1166),
.B(n_1109),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1165),
.B(n_1022),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1121),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1136),
.B(n_1109),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1132),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_R g1208 ( 
.A(n_1124),
.B(n_988),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1121),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1132),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1125),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1145),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1150),
.B(n_1090),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1150),
.B(n_1090),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1150),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1164),
.B(n_1042),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_1171),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1161),
.B(n_982),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1164),
.B(n_1026),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1116),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1171),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1138),
.B(n_1026),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1171),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1123),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1123),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1140),
.B(n_1042),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1131),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1160),
.B(n_1089),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1154),
.B(n_985),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1126),
.B(n_1060),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_1131),
.B(n_859),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1167),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1167),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1133),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1144),
.B(n_1089),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1168),
.Y(n_1236)
);

NOR2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1118),
.B(n_1119),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1120),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1168),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1141),
.A2(n_600),
.B1(n_604),
.B2(n_575),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1134),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1129),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1146),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1117),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1147),
.B(n_1036),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1149),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1117),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1155),
.B(n_1060),
.Y(n_1248)
);

AND2x6_ASAP7_75t_L g1249 ( 
.A(n_1151),
.B(n_709),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1186),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1186),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1174),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1202),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1202),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1205),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1173),
.B(n_1180),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1172),
.A2(n_1081),
.B1(n_931),
.B2(n_911),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1205),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1203),
.B(n_1206),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1191),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1172),
.B(n_1152),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1191),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1183),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1173),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1209),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1240),
.B(n_1033),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1216),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1203),
.B(n_1107),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1219),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1248),
.A2(n_1155),
.B1(n_1033),
.B2(n_1037),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1209),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1191),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1222),
.B(n_1034),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1176),
.Y(n_1274)
);

OAI221xp5_ASAP7_75t_L g1275 ( 
.A1(n_1184),
.A2(n_1178),
.B1(n_1187),
.B2(n_1190),
.C(n_1198),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1199),
.A2(n_626),
.B1(n_782),
.B2(n_741),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1210),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_SL g1278 ( 
.A(n_1220),
.B(n_988),
.Y(n_1278)
);

BUFx2_ASAP7_75t_SL g1279 ( 
.A(n_1247),
.Y(n_1279)
);

AO22x2_ASAP7_75t_L g1280 ( 
.A1(n_1196),
.A2(n_550),
.B1(n_726),
.B2(n_566),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1217),
.B(n_1036),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1208),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1206),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1203),
.B(n_1110),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1192),
.A2(n_1081),
.B1(n_931),
.B2(n_911),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1217),
.B(n_1084),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1206),
.B(n_789),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1223),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1208),
.Y(n_1289)
);

AO22x2_ASAP7_75t_L g1290 ( 
.A1(n_1194),
.A2(n_871),
.B1(n_872),
.B2(n_714),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1224),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1222),
.B(n_1034),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1224),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1192),
.B(n_1084),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1232),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1231),
.B(n_1084),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1184),
.A2(n_1231),
.B1(n_1235),
.B2(n_1236),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1232),
.Y(n_1299)
);

AO22x2_ASAP7_75t_L g1300 ( 
.A1(n_1195),
.A2(n_884),
.B1(n_654),
.B2(n_682),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1233),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1219),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1173),
.B(n_1110),
.Y(n_1303)
);

AO22x2_ASAP7_75t_L g1304 ( 
.A1(n_1229),
.A2(n_682),
.B1(n_788),
.B2(n_605),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1233),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1173),
.B(n_1111),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1180),
.B(n_1182),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1175),
.B(n_791),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1239),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1239),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1175),
.B(n_1089),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1200),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1247),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1181),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1200),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1225),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1211),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1207),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1207),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1180),
.B(n_1111),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1180),
.B(n_1102),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1225),
.Y(n_1322)
);

AO22x2_ASAP7_75t_L g1323 ( 
.A1(n_1218),
.A2(n_788),
.B1(n_818),
.B2(n_605),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1227),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1215),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1215),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1211),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1204),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1182),
.B(n_1102),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1221),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1204),
.B(n_1085),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1182),
.B(n_1085),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1226),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1197),
.B(n_1092),
.Y(n_1334)
);

OAI221xp5_ASAP7_75t_L g1335 ( 
.A1(n_1184),
.A2(n_897),
.B1(n_548),
.B2(n_573),
.C(n_557),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1221),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1182),
.B(n_800),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1235),
.A2(n_832),
.B1(n_844),
.B2(n_818),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1245),
.B(n_847),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1245),
.B(n_1037),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1227),
.Y(n_1341)
);

AOI211xp5_ASAP7_75t_L g1342 ( 
.A1(n_1234),
.A2(n_1020),
.B(n_1092),
.C(n_576),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1179),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1201),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1188),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1244),
.Y(n_1346)
);

AO22x2_ASAP7_75t_L g1347 ( 
.A1(n_1243),
.A2(n_844),
.B1(n_971),
.B2(n_832),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1246),
.A2(n_951),
.B1(n_977),
.B2(n_622),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1189),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1228),
.B(n_1089),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1228),
.A2(n_1049),
.B1(n_817),
.B2(n_614),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1237),
.B(n_773),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1261),
.A2(n_1242),
.B(n_1214),
.C(n_1213),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1286),
.A2(n_1212),
.B(n_1185),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1281),
.B(n_1249),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1350),
.A2(n_1212),
.B(n_1185),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1294),
.A2(n_1070),
.B(n_1242),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1275),
.A2(n_563),
.B(n_574),
.C(n_564),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1263),
.A2(n_618),
.B(n_625),
.C(n_587),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1250),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1331),
.B(n_1249),
.Y(n_1361)
);

AOI21xp33_ASAP7_75t_L g1362 ( 
.A1(n_1266),
.A2(n_1238),
.B(n_1049),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1314),
.B(n_1241),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1250),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1311),
.A2(n_1212),
.B(n_1193),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1297),
.A2(n_1070),
.B(n_1064),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1259),
.B(n_1212),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1296),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1283),
.B(n_1249),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1251),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1259),
.B(n_1343),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1343),
.A2(n_1193),
.B(n_1177),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1269),
.A2(n_630),
.B(n_646),
.C(n_628),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1345),
.A2(n_1177),
.B(n_1064),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1328),
.B(n_1009),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1345),
.A2(n_1064),
.B(n_1061),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1251),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1308),
.A2(n_1249),
.B1(n_612),
.B2(n_624),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1332),
.B(n_546),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1302),
.A2(n_702),
.B(n_706),
.C(n_658),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1349),
.A2(n_1064),
.B(n_1061),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1335),
.A2(n_731),
.B(n_739),
.C(n_723),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1264),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1349),
.A2(n_1329),
.B(n_1262),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1254),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_L g1386 ( 
.A(n_1339),
.B(n_843),
.C(n_590),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1340),
.A2(n_1267),
.B1(n_1292),
.B2(n_1273),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1329),
.A2(n_1061),
.B(n_1069),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1254),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1260),
.A2(n_1061),
.B(n_1069),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1272),
.A2(n_1069),
.B(n_1070),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1332),
.A2(n_1069),
.B(n_1057),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1252),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1306),
.A2(n_1071),
.B(n_1093),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1351),
.A2(n_764),
.B(n_767),
.C(n_752),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1274),
.B(n_1249),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1306),
.A2(n_1071),
.B(n_1093),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1334),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1268),
.B(n_546),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1298),
.B(n_1268),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1255),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1264),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1336),
.A2(n_1071),
.B(n_1093),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1255),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1336),
.A2(n_1097),
.B(n_1089),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1293),
.A2(n_1058),
.B(n_1054),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1276),
.A2(n_958),
.B1(n_960),
.B2(n_935),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1348),
.A2(n_777),
.B(n_811),
.C(n_809),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1321),
.A2(n_1097),
.B(n_1098),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1279),
.Y(n_1410)
);

AND2x2_ASAP7_75t_SL g1411 ( 
.A(n_1278),
.B(n_551),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1284),
.B(n_1257),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1299),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1284),
.A2(n_821),
.B(n_823),
.C(n_822),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1287),
.B(n_636),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1301),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1253),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1309),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1310),
.A2(n_1058),
.B(n_1054),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1270),
.B(n_631),
.C(n_629),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1277),
.A2(n_831),
.B(n_853),
.C(n_837),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1313),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1264),
.B(n_1352),
.Y(n_1423)
);

AOI21xp33_ASAP7_75t_L g1424 ( 
.A1(n_1333),
.A2(n_969),
.B(n_962),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1338),
.B(n_1094),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1282),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1312),
.A2(n_1097),
.B(n_1098),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1258),
.A2(n_1097),
.B(n_1087),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1315),
.A2(n_728),
.B(n_551),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1304),
.B(n_778),
.Y(n_1430)
);

O2A1O1Ixp5_ASAP7_75t_L g1431 ( 
.A1(n_1337),
.A2(n_1087),
.B(n_1082),
.C(n_895),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1342),
.B(n_552),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1318),
.A2(n_728),
.B(n_551),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1338),
.B(n_1288),
.Y(n_1434)
);

AOI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1319),
.A2(n_1066),
.B(n_1063),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1325),
.A2(n_1066),
.B(n_1063),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1326),
.A2(n_728),
.B(n_551),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1317),
.B(n_1009),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1330),
.A2(n_728),
.B(n_551),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1285),
.B(n_1094),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1256),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1307),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1303),
.A2(n_770),
.B(n_728),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1265),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1271),
.A2(n_896),
.B(n_880),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1346),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1320),
.A2(n_921),
.B(n_770),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1327),
.B(n_1009),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1291),
.A2(n_921),
.B(n_770),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1347),
.B(n_1096),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1383),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1387),
.B(n_1289),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1413),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

O2A1O1Ixp5_ASAP7_75t_L g1455 ( 
.A1(n_1395),
.A2(n_1352),
.B(n_1295),
.C(n_1305),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1383),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1446),
.B(n_1344),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1374),
.A2(n_1322),
.B(n_1316),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1368),
.B(n_1347),
.Y(n_1459)
);

NOR3xp33_ASAP7_75t_SL g1460 ( 
.A(n_1420),
.B(n_555),
.C(n_547),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1368),
.B(n_1304),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1362),
.B(n_1324),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1386),
.A2(n_1341),
.B(n_907),
.C(n_948),
.Y(n_1463)
);

NOR2xp67_ASAP7_75t_L g1464 ( 
.A(n_1371),
.B(n_369),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1385),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_R g1466 ( 
.A(n_1426),
.B(n_552),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1411),
.A2(n_1400),
.B1(n_1398),
.B2(n_1412),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1415),
.B(n_1323),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1407),
.A2(n_1290),
.B1(n_1300),
.B2(n_1280),
.C(n_1323),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1353),
.A2(n_921),
.B(n_770),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1422),
.B(n_980),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1401),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1355),
.A2(n_921),
.B(n_770),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1361),
.A2(n_965),
.B(n_921),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1408),
.A2(n_553),
.B(n_580),
.C(n_579),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1378),
.B(n_371),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1434),
.A2(n_1280),
.B1(n_1290),
.B2(n_1300),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1360),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1384),
.A2(n_565),
.B1(n_568),
.B2(n_562),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1422),
.B(n_562),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1372),
.A2(n_965),
.B(n_1082),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1373),
.A2(n_594),
.B(n_603),
.C(n_588),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1363),
.A2(n_568),
.B1(n_570),
.B2(n_565),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1418),
.A2(n_572),
.B1(n_578),
.B2(n_570),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1393),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1364),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1403),
.A2(n_952),
.B(n_923),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1357),
.A2(n_965),
.B(n_954),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1423),
.B(n_778),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1423),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1370),
.B(n_1377),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1424),
.B(n_572),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1380),
.A2(n_608),
.B(n_617),
.C(n_607),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1389),
.B(n_1404),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1410),
.B(n_1375),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1438),
.B(n_708),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1402),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1399),
.B(n_1379),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1402),
.B(n_773),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1444),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1430),
.B(n_778),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1396),
.A2(n_591),
.B1(n_592),
.B2(n_578),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1442),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1417),
.B(n_591),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1432),
.B(n_592),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1357),
.A2(n_965),
.B(n_1076),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1359),
.A2(n_627),
.B(n_635),
.C(n_621),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1441),
.B(n_1096),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1450),
.B(n_601),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1369),
.A2(n_609),
.B1(n_610),
.B2(n_601),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1441),
.B(n_609),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1354),
.A2(n_965),
.B(n_1076),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1425),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1365),
.A2(n_1080),
.B(n_1076),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1406),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1392),
.A2(n_1083),
.B(n_1080),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1367),
.A2(n_747),
.B1(n_893),
.B2(n_610),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1448),
.B(n_1442),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1356),
.A2(n_1083),
.B(n_1080),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1442),
.B(n_644),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1358),
.A2(n_1440),
.B1(n_1414),
.B2(n_1445),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1431),
.B(n_857),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1421),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1382),
.B(n_747),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1443),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1428),
.B(n_1376),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1419),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1388),
.A2(n_900),
.B1(n_913),
.B2(n_893),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1435),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_SL g1530 ( 
.A1(n_1429),
.A2(n_651),
.B(n_656),
.C(n_645),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1428),
.B(n_900),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1436),
.B(n_663),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1381),
.A2(n_1083),
.B(n_633),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1447),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_SL g1535 ( 
.A1(n_1433),
.A2(n_1104),
.B(n_1100),
.C(n_664),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1409),
.A2(n_634),
.B(n_623),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1366),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1427),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1394),
.A2(n_637),
.B1(n_648),
.B2(n_642),
.Y(n_1539)
);

NOR2xp67_ASAP7_75t_SL g1540 ( 
.A(n_1397),
.B(n_547),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1390),
.A2(n_661),
.B(n_659),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1391),
.B(n_555),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1405),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1437),
.B(n_913),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1439),
.Y(n_1545)
);

O2A1O1Ixp5_ASAP7_75t_L g1546 ( 
.A1(n_1449),
.A2(n_672),
.B(n_673),
.C(n_669),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1413),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1422),
.B(n_1067),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1387),
.B(n_915),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1413),
.Y(n_1550)
);

INVx5_ASAP7_75t_L g1551 ( 
.A(n_1383),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1442),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1485),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1552),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1549),
.A2(n_667),
.B1(n_680),
.B2(n_666),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1548),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1461),
.B(n_708),
.Y(n_1557)
);

INVx5_ASAP7_75t_L g1558 ( 
.A(n_1552),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1552),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1480),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1467),
.B(n_558),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1457),
.B(n_674),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1457),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1453),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1497),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1454),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

NAND2x1_ASAP7_75t_L g1568 ( 
.A(n_1478),
.B(n_1067),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1486),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1489),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1551),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1551),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

INVx5_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1490),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1465),
.Y(n_1576)
);

BUFx2_ASAP7_75t_R g1577 ( 
.A(n_1471),
.Y(n_1577)
);

BUFx12f_ASAP7_75t_L g1578 ( 
.A(n_1520),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1527),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1503),
.Y(n_1580)
);

INVx3_ASAP7_75t_SL g1581 ( 
.A(n_1520),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_SL g1582 ( 
.A(n_1503),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1462),
.B(n_1452),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1490),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1495),
.Y(n_1585)
);

BUFx4f_ASAP7_75t_SL g1586 ( 
.A(n_1518),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1451),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1459),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1451),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1513),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1511),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1456),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1491),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1508),
.B(n_376),
.Y(n_1594)
);

BUFx5_ASAP7_75t_L g1595 ( 
.A(n_1538),
.Y(n_1595)
);

BUFx2_ASAP7_75t_SL g1596 ( 
.A(n_1456),
.Y(n_1596)
);

INVx5_ASAP7_75t_SL g1597 ( 
.A(n_1508),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1494),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1492),
.B(n_558),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1472),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1550),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1515),
.Y(n_1602)
);

NAND2x1p5_ASAP7_75t_L g1603 ( 
.A(n_1500),
.B(n_1464),
.Y(n_1603)
);

INVx5_ASAP7_75t_L g1604 ( 
.A(n_1523),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1532),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1498),
.A2(n_560),
.B1(n_567),
.B2(n_561),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1499),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1529),
.Y(n_1608)
);

BUFx8_ASAP7_75t_L g1609 ( 
.A(n_1501),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1532),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1455),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1469),
.A2(n_711),
.B1(n_857),
.B2(n_756),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1526),
.Y(n_1613)
);

BUFx2_ASAP7_75t_R g1614 ( 
.A(n_1468),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1464),
.B(n_1068),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1542),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1543),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1509),
.B(n_1477),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1475),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1458),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1460),
.B(n_377),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1525),
.Y(n_1622)
);

BUFx2_ASAP7_75t_SL g1623 ( 
.A(n_1476),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1487),
.Y(n_1624)
);

INVx6_ASAP7_75t_SL g1625 ( 
.A(n_1466),
.Y(n_1625)
);

BUFx2_ASAP7_75t_SL g1626 ( 
.A(n_1476),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1504),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1505),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1534),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1483),
.B(n_559),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1522),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1496),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1544),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1521),
.A2(n_683),
.B1(n_687),
.B2(n_681),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1524),
.A2(n_711),
.B1(n_857),
.B2(n_756),
.Y(n_1635)
);

AOI222xp33_ASAP7_75t_L g1636 ( 
.A1(n_1583),
.A2(n_696),
.B1(n_685),
.B2(n_710),
.C1(n_686),
.C2(n_677),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1563),
.Y(n_1637)
);

INVx6_ASAP7_75t_L g1638 ( 
.A(n_1574),
.Y(n_1638)
);

AO31x2_ASAP7_75t_L g1639 ( 
.A1(n_1624),
.A2(n_1470),
.A3(n_1488),
.B(n_1506),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1589),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1624),
.A2(n_1512),
.B(n_1473),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1620),
.A2(n_1474),
.B(n_1514),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1620),
.A2(n_1519),
.B(n_1516),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1611),
.A2(n_1481),
.B(n_1545),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1573),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1604),
.A2(n_1531),
.B(n_1533),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1623),
.B(n_1536),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1573),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1632),
.A2(n_1463),
.B1(n_1484),
.B2(n_1517),
.Y(n_1649)
);

O2A1O1Ixp33_ASAP7_75t_SL g1650 ( 
.A1(n_1618),
.A2(n_1507),
.B(n_1535),
.C(n_1528),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1569),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1579),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1634),
.A2(n_1541),
.B(n_1539),
.Y(n_1653)
);

AOI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1579),
.A2(n_1540),
.B(n_1502),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1613),
.A2(n_1546),
.B(n_1493),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1613),
.B(n_1510),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1608),
.Y(n_1657)
);

INVx5_ASAP7_75t_L g1658 ( 
.A(n_1604),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1626),
.B(n_1631),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1625),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1576),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1616),
.A2(n_1479),
.B1(n_638),
.B2(n_639),
.Y(n_1662)
);

INVx3_ASAP7_75t_SL g1663 ( 
.A(n_1581),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1608),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1564),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1617),
.A2(n_1482),
.B(n_1072),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1566),
.Y(n_1667)
);

AO31x2_ASAP7_75t_L g1668 ( 
.A1(n_1602),
.A2(n_712),
.A3(n_720),
.B(n_719),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1617),
.A2(n_1072),
.B(n_1068),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1590),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1590),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1567),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1602),
.A2(n_1530),
.B(n_732),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1603),
.A2(n_1104),
.B(n_1100),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1588),
.B(n_1631),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1629),
.A2(n_1104),
.B(n_1100),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1629),
.A2(n_1605),
.B(n_1610),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1589),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1605),
.A2(n_1104),
.B(n_1100),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1622),
.A2(n_1593),
.B(n_1594),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1619),
.A2(n_735),
.B(n_721),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1599),
.A2(n_749),
.B1(n_750),
.B2(n_748),
.Y(n_1682)
);

AND2x4_ASAP7_75t_SL g1683 ( 
.A(n_1571),
.B(n_711),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1553),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1565),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1595),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1600),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1568),
.A2(n_753),
.B(n_751),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1606),
.A2(n_905),
.B1(n_940),
.B2(n_589),
.C(n_560),
.Y(n_1689)
);

AO31x2_ASAP7_75t_L g1690 ( 
.A1(n_1598),
.A2(n_763),
.A3(n_793),
.B(n_780),
.Y(n_1690)
);

OAI211xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1630),
.A2(n_816),
.B(n_842),
.C(n_807),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1600),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1586),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1598),
.A2(n_850),
.B(n_848),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1645),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_1631),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1648),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1686),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1652),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1641),
.A2(n_1635),
.B(n_1612),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1671),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1677),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1657),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1664),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1672),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1675),
.B(n_1633),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1665),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1691),
.A2(n_1591),
.B1(n_1561),
.B2(n_1627),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1660),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1667),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1668),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1668),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1658),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1691),
.A2(n_1628),
.B1(n_1621),
.B2(n_1560),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1644),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1684),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1668),
.Y(n_1718)
);

OR2x6_ASAP7_75t_L g1719 ( 
.A(n_1680),
.B(n_1633),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1668),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1690),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1658),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1690),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1690),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1643),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1658),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1642),
.A2(n_1646),
.B(n_1676),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1651),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1658),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1661),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1639),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1669),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1685),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1694),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1639),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1659),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1659),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1639),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1694),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1639),
.B(n_1595),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1646),
.A2(n_1615),
.B(n_1595),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1735),
.B(n_1637),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1717),
.Y(n_1745)
);

INVx5_ASAP7_75t_SL g1746 ( 
.A(n_1719),
.Y(n_1746)
);

AO31x2_ASAP7_75t_L g1747 ( 
.A1(n_1713),
.A2(n_1656),
.A3(n_1572),
.B(n_1687),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1719),
.B(n_1659),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1735),
.B(n_1637),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1706),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1717),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1698),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1706),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1696),
.B(n_1692),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1709),
.A2(n_1682),
.B1(n_1604),
.B2(n_1649),
.Y(n_1755)
);

NAND2xp33_ASAP7_75t_R g1756 ( 
.A(n_1710),
.B(n_1585),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1723),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_R g1758 ( 
.A(n_1738),
.B(n_1660),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1707),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1696),
.B(n_1663),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1715),
.B(n_1636),
.C(n_1681),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1711),
.Y(n_1762)
);

BUFx4f_ASAP7_75t_SL g1763 ( 
.A(n_1707),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1696),
.Y(n_1764)
);

CKINVDCx16_ASAP7_75t_R g1765 ( 
.A(n_1739),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1719),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_L g1767 ( 
.A1(n_1715),
.A2(n_1636),
.B(n_1682),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1696),
.B(n_1663),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1719),
.A2(n_1621),
.B1(n_1578),
.B2(n_1633),
.Y(n_1769)
);

NOR3xp33_ASAP7_75t_SL g1770 ( 
.A(n_1736),
.B(n_1681),
.C(n_1689),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1719),
.B(n_1638),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1719),
.A2(n_1653),
.B1(n_1689),
.B2(n_1609),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1696),
.B(n_1693),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1723),
.B(n_1640),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1698),
.B(n_1570),
.Y(n_1775)
);

NOR2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1640),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1711),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1706),
.B(n_1595),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1739),
.Y(n_1779)
);

NAND2xp33_ASAP7_75t_R g1780 ( 
.A(n_1738),
.B(n_1562),
.Y(n_1780)
);

OR2x6_ASAP7_75t_L g1781 ( 
.A(n_1743),
.B(n_1638),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1709),
.B(n_1607),
.Y(n_1782)
);

BUFx4f_ASAP7_75t_SL g1783 ( 
.A(n_1738),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1711),
.B(n_1678),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1697),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1708),
.B(n_1595),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1738),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1695),
.B(n_1678),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1697),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1708),
.B(n_1614),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_SL g1791 ( 
.A(n_1736),
.B(n_1555),
.C(n_1662),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1730),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1704),
.B(n_1557),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1743),
.B(n_1638),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1730),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1704),
.B(n_1705),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1759),
.B(n_1703),
.Y(n_1797)
);

INVx2_ASAP7_75t_SL g1798 ( 
.A(n_1776),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1750),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1753),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1785),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1761),
.A2(n_1653),
.B(n_1743),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1789),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1792),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1770),
.B(n_1726),
.C(n_1741),
.Y(n_1806)
);

AND2x4_ASAP7_75t_SL g1807 ( 
.A(n_1748),
.B(n_1728),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1762),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1777),
.Y(n_1809)
);

AND2x4_ASAP7_75t_SL g1810 ( 
.A(n_1748),
.B(n_1728),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1795),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1752),
.B(n_1703),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1744),
.B(n_1749),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1796),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1771),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1787),
.B(n_1703),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1771),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1747),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1783),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1781),
.B(n_1794),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1765),
.B(n_1745),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1751),
.B(n_1703),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1757),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1781),
.B(n_1794),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1786),
.Y(n_1826)
);

CKINVDCx12_ASAP7_75t_R g1827 ( 
.A(n_1775),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1748),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1801),
.Y(n_1829)
);

INVx4_ASAP7_75t_R g1830 ( 
.A(n_1820),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1822),
.B(n_1774),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1824),
.B(n_1779),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1801),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1801),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1760),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1798),
.B(n_1828),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1822),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1814),
.B(n_1768),
.Y(n_1838)
);

AOI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1812),
.A2(n_1782),
.B(n_1755),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1802),
.A2(n_1761),
.B(n_1755),
.C(n_1767),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1802),
.A2(n_1767),
.B1(n_1772),
.B2(n_1770),
.C(n_1769),
.Y(n_1841)
);

INVx4_ASAP7_75t_SL g1842 ( 
.A(n_1820),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1803),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1803),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1814),
.B(n_1773),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1824),
.B(n_1793),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1806),
.A2(n_1791),
.B(n_1771),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1803),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1800),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1821),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1823),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1800),
.Y(n_1852)
);

AOI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1806),
.A2(n_1791),
.B(n_1793),
.C(n_881),
.Y(n_1853)
);

OAI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1828),
.A2(n_561),
.B(n_559),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1798),
.A2(n_1650),
.B(n_1647),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1828),
.Y(n_1856)
);

OAI21x1_ASAP7_75t_L g1857 ( 
.A1(n_1813),
.A2(n_1725),
.B(n_1716),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1798),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1799),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1848),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1851),
.B(n_1826),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1837),
.B(n_1840),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1829),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1849),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1836),
.B(n_1821),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1842),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1836),
.B(n_1821),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1852),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1833),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1850),
.B(n_1821),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_SL g1871 ( 
.A(n_1841),
.B(n_1766),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1846),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1858),
.Y(n_1873)
);

INVx4_ASAP7_75t_L g1874 ( 
.A(n_1842),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1856),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1834),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1850),
.B(n_1825),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1853),
.A2(n_1746),
.B1(n_1818),
.B2(n_1816),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1856),
.B(n_1826),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1843),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1844),
.B(n_1805),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1859),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1832),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1856),
.B(n_1825),
.Y(n_1884)
);

INVxp67_ASAP7_75t_SL g1885 ( 
.A(n_1839),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1831),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1857),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1830),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1830),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1847),
.B(n_1838),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1845),
.Y(n_1891)
);

INVx5_ASAP7_75t_SL g1892 ( 
.A(n_1854),
.Y(n_1892)
);

NOR3xp33_ASAP7_75t_L g1893 ( 
.A(n_1862),
.B(n_1854),
.C(n_1466),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1865),
.B(n_1825),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1866),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1865),
.B(n_1825),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1864),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1873),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1867),
.B(n_1835),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1864),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1888),
.B(n_1823),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1874),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1867),
.B(n_1816),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1874),
.B(n_1807),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1863),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1888),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1868),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1874),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1884),
.B(n_1818),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1884),
.B(n_1810),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1871),
.B(n_1758),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1868),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1875),
.B(n_1810),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1869),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1872),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1889),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1875),
.B(n_1810),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1861),
.B(n_1805),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1869),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1863),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1861),
.B(n_1804),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1876),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1889),
.B(n_1812),
.Y(n_1923)
);

NAND2x1_ASAP7_75t_L g1924 ( 
.A(n_1904),
.B(n_1874),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1908),
.Y(n_1925)
);

NAND2x1p5_ASAP7_75t_L g1926 ( 
.A(n_1904),
.B(n_1875),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1898),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1915),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1897),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1895),
.B(n_1883),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1902),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1902),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1897),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1906),
.B(n_1890),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1908),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1916),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1899),
.B(n_1891),
.Y(n_1937)
);

NAND2x1p5_ASAP7_75t_L g1938 ( 
.A(n_1904),
.B(n_1574),
.Y(n_1938)
);

NOR2xp67_ASAP7_75t_L g1939 ( 
.A(n_1908),
.B(n_1877),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1899),
.B(n_1891),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1900),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1910),
.B(n_1909),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1893),
.B(n_1871),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1911),
.B(n_1878),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1900),
.B(n_1886),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1907),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1907),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1910),
.B(n_1883),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1913),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1923),
.B(n_1886),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1912),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1909),
.B(n_1870),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1912),
.Y(n_1953)
);

NAND2x1p5_ASAP7_75t_L g1954 ( 
.A(n_1913),
.B(n_1574),
.Y(n_1954)
);

O2A1O1Ixp33_ASAP7_75t_L g1955 ( 
.A1(n_1914),
.A2(n_1885),
.B(n_1892),
.C(n_1879),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1901),
.B(n_1881),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1903),
.B(n_1892),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1903),
.B(n_1870),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1914),
.B(n_1860),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1919),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1919),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1920),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1905),
.B(n_1860),
.Y(n_1963)
);

INVxp67_ASAP7_75t_L g1964 ( 
.A(n_1917),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1917),
.Y(n_1965)
);

AND2x2_ASAP7_75t_SL g1966 ( 
.A(n_1894),
.B(n_1683),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1918),
.B(n_1881),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1927),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1926),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1930),
.B(n_1918),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1924),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1942),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1934),
.A2(n_1892),
.B1(n_1780),
.B2(n_1855),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1931),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1936),
.B(n_1892),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1931),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1936),
.B(n_1894),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1949),
.B(n_1896),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1932),
.Y(n_1979)
);

CKINVDCx16_ASAP7_75t_R g1980 ( 
.A(n_1944),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1964),
.B(n_1896),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1932),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1965),
.B(n_1905),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1929),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1939),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1928),
.B(n_1625),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1925),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1937),
.B(n_1922),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1952),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1933),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1941),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1940),
.B(n_1922),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1946),
.Y(n_1993)
);

INVx1_ASAP7_75t_SL g1994 ( 
.A(n_1935),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1948),
.B(n_1877),
.Y(n_1995)
);

INVx4_ASAP7_75t_L g1996 ( 
.A(n_1966),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1947),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1957),
.B(n_1877),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1958),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1944),
.B(n_1877),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1951),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1938),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1943),
.B(n_1920),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1953),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_L g2005 ( 
.A(n_1939),
.B(n_1921),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1944),
.A2(n_1921),
.B1(n_1790),
.B2(n_1813),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1960),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1956),
.B(n_1876),
.Y(n_2008)
);

OR2x6_ASAP7_75t_L g2009 ( 
.A(n_1955),
.B(n_1562),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1961),
.Y(n_2010)
);

OAI33xp33_ASAP7_75t_L g2011 ( 
.A1(n_1945),
.A2(n_584),
.A3(n_569),
.B1(n_586),
.B2(n_577),
.B3(n_567),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1962),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1954),
.B(n_1880),
.Y(n_2013)
);

OR2x6_ASAP7_75t_L g2014 ( 
.A(n_1967),
.B(n_1607),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1950),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1959),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1945),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1963),
.B(n_1880),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1963),
.B(n_1882),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1959),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1936),
.B(n_1882),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1927),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1942),
.B(n_1797),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1927),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_1936),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1966),
.B(n_1763),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1927),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1927),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1944),
.A2(n_1746),
.B1(n_1887),
.B2(n_1807),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1927),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1927),
.B(n_1887),
.Y(n_2031)
);

OAI31xp33_ASAP7_75t_L g2032 ( 
.A1(n_2006),
.A2(n_2025),
.A3(n_1979),
.B(n_2028),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_2025),
.B(n_1971),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2030),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1969),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2005),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2000),
.B(n_1807),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1978),
.B(n_1797),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1980),
.B(n_1815),
.Y(n_2039)
);

NOR3xp33_ASAP7_75t_SL g2040 ( 
.A(n_1975),
.B(n_1756),
.C(n_577),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1977),
.B(n_1815),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1985),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1979),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1972),
.B(n_1974),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1995),
.B(n_1813),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1970),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1976),
.B(n_1804),
.Y(n_2047)
);

AND3x2_ASAP7_75t_L g2048 ( 
.A(n_1982),
.B(n_1556),
.C(n_1609),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1968),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2022),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1987),
.B(n_1813),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1987),
.B(n_1817),
.Y(n_2052)
);

NOR2xp67_ASAP7_75t_SL g2053 ( 
.A(n_1996),
.B(n_1571),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1996),
.B(n_1827),
.Y(n_2054)
);

INVx4_ASAP7_75t_L g2055 ( 
.A(n_2024),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1994),
.B(n_1817),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1994),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2027),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2021),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1988),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1992),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1981),
.B(n_1811),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_2026),
.A2(n_2006),
.B(n_2009),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1989),
.B(n_854),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1999),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1998),
.A2(n_1746),
.B1(n_1794),
.B2(n_1781),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2015),
.B(n_2020),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2003),
.B(n_883),
.Y(n_2068)
);

AOI22x1_ASAP7_75t_L g2069 ( 
.A1(n_2002),
.A2(n_2013),
.B1(n_2016),
.B2(n_2017),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1986),
.B(n_1808),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2009),
.B(n_1808),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2009),
.B(n_1808),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2023),
.B(n_1809),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1983),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_2014),
.Y(n_2075)
);

CKINVDCx16_ASAP7_75t_R g2076 ( 
.A(n_1973),
.Y(n_2076)
);

BUFx2_ASAP7_75t_L g2077 ( 
.A(n_2014),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1984),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1990),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2018),
.B(n_901),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2012),
.B(n_902),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_2014),
.Y(n_2082)
);

NAND2xp33_ASAP7_75t_L g2083 ( 
.A(n_1973),
.B(n_569),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1991),
.B(n_1993),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2029),
.B(n_1809),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2019),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1997),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2001),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2004),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2007),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2008),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2010),
.Y(n_2092)
);

OAI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_2031),
.A2(n_1683),
.B(n_1577),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2031),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2011),
.Y(n_2095)
);

NAND3xp33_ASAP7_75t_SL g2096 ( 
.A(n_2025),
.B(n_589),
.C(n_586),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_2028),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2025),
.B(n_903),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_SL g2099 ( 
.A(n_1980),
.B(n_1582),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2005),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2025),
.B(n_1811),
.Y(n_2101)
);

NAND2x1p5_ASAP7_75t_L g2102 ( 
.A(n_2025),
.B(n_1558),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2025),
.B(n_908),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2025),
.B(n_1809),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2028),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2028),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2000),
.B(n_1799),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2028),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2028),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2000),
.B(n_1799),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2005),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_2025),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2028),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2005),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2028),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2025),
.B(n_910),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2000),
.B(n_1754),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2025),
.B(n_914),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2033),
.B(n_919),
.Y(n_2119)
);

OAI322xp33_ASAP7_75t_L g2120 ( 
.A1(n_2112),
.A2(n_2097),
.A3(n_2043),
.B1(n_2076),
.B2(n_2113),
.C1(n_2115),
.C2(n_2034),
.Y(n_2120)
);

O2A1O1Ixp33_ASAP7_75t_SL g2121 ( 
.A1(n_2057),
.A2(n_927),
.B(n_930),
.C(n_920),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2033),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_2032),
.A2(n_593),
.B(n_584),
.Y(n_2123)
);

NOR3xp33_ASAP7_75t_L g2124 ( 
.A(n_2083),
.B(n_934),
.C(n_933),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2034),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2035),
.Y(n_2126)
);

AOI21xp33_ASAP7_75t_L g2127 ( 
.A1(n_2054),
.A2(n_595),
.B(n_593),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2105),
.A2(n_957),
.B1(n_950),
.B2(n_942),
.C(n_598),
.Y(n_2128)
);

NOR3xp33_ASAP7_75t_L g2129 ( 
.A(n_2044),
.B(n_596),
.C(n_595),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2113),
.Y(n_2130)
);

OA21x2_ASAP7_75t_L g2131 ( 
.A1(n_2036),
.A2(n_598),
.B(n_596),
.Y(n_2131)
);

OAI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2063),
.A2(n_611),
.B(n_606),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2035),
.B(n_2046),
.Y(n_2133)
);

AOI222xp33_ASAP7_75t_L g2134 ( 
.A1(n_2100),
.A2(n_775),
.B1(n_611),
.B2(n_894),
.C1(n_774),
.C2(n_606),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2042),
.B(n_2106),
.Y(n_2135)
);

NOR3xp33_ASAP7_75t_L g2136 ( 
.A(n_2055),
.B(n_775),
.C(n_774),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2115),
.B(n_894),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_2108),
.B(n_0),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2055),
.B(n_898),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2037),
.B(n_1754),
.Y(n_2140)
);

OAI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2111),
.A2(n_904),
.B(n_898),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2109),
.Y(n_2142)
);

OAI32xp33_ASAP7_75t_L g2143 ( 
.A1(n_2114),
.A2(n_1819),
.A3(n_906),
.B1(n_909),
.B2(n_905),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2091),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2048),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2096),
.A2(n_906),
.B(n_904),
.Y(n_2146)
);

NAND3xp33_ASAP7_75t_L g2147 ( 
.A(n_2069),
.B(n_912),
.C(n_909),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_2099),
.B(n_1827),
.Y(n_2148)
);

OAI221xp5_ASAP7_75t_L g2149 ( 
.A1(n_2093),
.A2(n_924),
.B1(n_932),
.B2(n_917),
.C(n_912),
.Y(n_2149)
);

AOI221xp5_ASAP7_75t_L g2150 ( 
.A1(n_2049),
.A2(n_932),
.B1(n_936),
.B2(n_924),
.C(n_917),
.Y(n_2150)
);

AO22x1_ASAP7_75t_L g2151 ( 
.A1(n_2051),
.A2(n_1558),
.B1(n_940),
.B2(n_943),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2065),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2045),
.A2(n_943),
.B1(n_944),
.B2(n_936),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2040),
.B(n_2038),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2067),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_2117),
.A2(n_2095),
.B1(n_2061),
.B2(n_2060),
.Y(n_2156)
);

NOR2x1_ASAP7_75t_L g2157 ( 
.A(n_2116),
.B(n_1594),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2118),
.Y(n_2158)
);

OAI21xp5_ASAP7_75t_SL g2159 ( 
.A1(n_2039),
.A2(n_1607),
.B(n_1722),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2075),
.B(n_944),
.Y(n_2160)
);

NAND2xp33_ASAP7_75t_SL g2161 ( 
.A(n_2053),
.B(n_1582),
.Y(n_2161)
);

OAI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_2050),
.A2(n_2058),
.B(n_2059),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2086),
.Y(n_2163)
);

AOI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_2094),
.A2(n_975),
.B1(n_976),
.B2(n_949),
.C(n_946),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2074),
.B(n_1764),
.Y(n_2165)
);

OAI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_2102),
.A2(n_1819),
.B1(n_1714),
.B2(n_1731),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2089),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2077),
.B(n_946),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2089),
.Y(n_2169)
);

AO22x1_ASAP7_75t_L g2170 ( 
.A1(n_2051),
.A2(n_1558),
.B1(n_975),
.B2(n_976),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2090),
.Y(n_2171)
);

OAI33xp33_ASAP7_75t_L g2172 ( 
.A1(n_2084),
.A2(n_978),
.A3(n_979),
.B1(n_949),
.B2(n_653),
.B3(n_643),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2090),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2082),
.Y(n_2174)
);

OR4x1_ASAP7_75t_L g2175 ( 
.A(n_2078),
.B(n_1559),
.C(n_1554),
.D(n_1741),
.Y(n_2175)
);

INVx1_ASAP7_75t_SL g2176 ( 
.A(n_2104),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2092),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_2101),
.Y(n_2178)
);

INVxp67_ASAP7_75t_L g2179 ( 
.A(n_2082),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2070),
.B(n_2107),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2092),
.Y(n_2181)
);

OAI31xp33_ASAP7_75t_L g2182 ( 
.A1(n_2085),
.A2(n_1714),
.A3(n_1650),
.B(n_1722),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2068),
.B(n_978),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2066),
.A2(n_1819),
.B1(n_979),
.B2(n_1705),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2098),
.B(n_632),
.Y(n_2185)
);

INVx1_ASAP7_75t_SL g2186 ( 
.A(n_2052),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2110),
.Y(n_2187)
);

OAI21xp5_ASAP7_75t_SL g2188 ( 
.A1(n_2047),
.A2(n_1731),
.B(n_1722),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2081),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2073),
.Y(n_2190)
);

A2O1A1Ixp33_ASAP7_75t_L g2191 ( 
.A1(n_2103),
.A2(n_655),
.B(n_657),
.C(n_649),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2080),
.B(n_662),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2064),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2079),
.B(n_1784),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_2071),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2087),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2088),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2041),
.Y(n_2198)
);

OAI221xp5_ASAP7_75t_L g2199 ( 
.A1(n_2056),
.A2(n_671),
.B1(n_675),
.B2(n_668),
.C(n_665),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2072),
.B(n_2062),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2033),
.B(n_676),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_2057),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2057),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_2112),
.B(n_679),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_2032),
.A2(n_691),
.B(n_684),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2112),
.B(n_694),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2057),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2057),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2033),
.Y(n_2209)
);

AOI222xp33_ASAP7_75t_L g2210 ( 
.A1(n_2083),
.A2(n_695),
.B1(n_699),
.B2(n_707),
.C1(n_700),
.C2(n_697),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_2032),
.A2(n_1724),
.B1(n_1721),
.B2(n_1712),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2112),
.B(n_1788),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2033),
.Y(n_2213)
);

AOI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2032),
.A2(n_722),
.B(n_718),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2112),
.B(n_1788),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2112),
.B(n_1597),
.Y(n_2216)
);

OAI221xp5_ASAP7_75t_SL g2217 ( 
.A1(n_2032),
.A2(n_1647),
.B1(n_1714),
.B2(n_1731),
.C(n_1722),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2033),
.B(n_724),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2057),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2032),
.A2(n_734),
.B(n_730),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2057),
.Y(n_2221)
);

OA22x2_ASAP7_75t_L g2222 ( 
.A1(n_2048),
.A2(n_737),
.B1(n_742),
.B2(n_736),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2076),
.A2(n_808),
.B1(n_860),
.B2(n_796),
.Y(n_2223)
);

AOI221xp5_ASAP7_75t_L g2224 ( 
.A1(n_2032),
.A2(n_746),
.B1(n_754),
.B2(n_745),
.C(n_744),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2033),
.B(n_755),
.Y(n_2225)
);

OAI322xp33_ASAP7_75t_SL g2226 ( 
.A1(n_2043),
.A2(n_771),
.A3(n_768),
.B1(n_776),
.B2(n_779),
.C1(n_769),
.C2(n_765),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_2053),
.B(n_1571),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_2033),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2033),
.B(n_790),
.Y(n_2229)
);

OAI211xp5_ASAP7_75t_L g2230 ( 
.A1(n_2032),
.A2(n_799),
.B(n_802),
.C(n_798),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2099),
.A2(n_803),
.B1(n_805),
.B2(n_804),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2033),
.B(n_810),
.Y(n_2232)
);

NOR2x2_ASAP7_75t_L g2233 ( 
.A(n_2091),
.B(n_1647),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2057),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2112),
.B(n_814),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2099),
.A2(n_815),
.B1(n_833),
.B2(n_825),
.Y(n_2236)
);

AOI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_2032),
.A2(n_839),
.B(n_834),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2112),
.B(n_1597),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2033),
.B(n_840),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2033),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_2112),
.B(n_1721),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2057),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2112),
.B(n_1575),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2033),
.Y(n_2244)
);

NAND2x1_ASAP7_75t_L g2245 ( 
.A(n_2033),
.B(n_1580),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2033),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_2032),
.A2(n_849),
.B(n_845),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2057),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2057),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_2032),
.A2(n_1724),
.B1(n_1718),
.B2(n_1720),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2076),
.A2(n_1786),
.B1(n_1718),
.B2(n_1720),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2033),
.B(n_851),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2112),
.B(n_1584),
.Y(n_2253)
);

NOR3xp33_ASAP7_75t_L g2254 ( 
.A(n_2076),
.B(n_856),
.C(n_852),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_2033),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2057),
.Y(n_2256)
);

OAI31xp33_ASAP7_75t_L g2257 ( 
.A1(n_2032),
.A2(n_1731),
.A3(n_1712),
.B(n_1725),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2057),
.Y(n_2258)
);

INVxp67_ASAP7_75t_SL g2259 ( 
.A(n_2057),
.Y(n_2259)
);

AOI322xp5_ASAP7_75t_L g2260 ( 
.A1(n_2112),
.A2(n_864),
.A3(n_862),
.B1(n_866),
.B2(n_867),
.C1(n_863),
.C2(n_858),
.Y(n_2260)
);

INVx2_ASAP7_75t_SL g2261 ( 
.A(n_2033),
.Y(n_2261)
);

OAI21xp33_ASAP7_75t_L g2262 ( 
.A1(n_2099),
.A2(n_869),
.B(n_868),
.Y(n_2262)
);

XOR2x2_ASAP7_75t_L g2263 ( 
.A(n_2054),
.B(n_2),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2076),
.A2(n_956),
.B1(n_970),
.B2(n_873),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2112),
.B(n_870),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2057),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2033),
.B(n_875),
.Y(n_2267)
);

AOI21xp33_ASAP7_75t_SL g2268 ( 
.A1(n_2032),
.A2(n_885),
.B(n_882),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2255),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2255),
.B(n_2228),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2261),
.B(n_887),
.Y(n_2271)
);

INVxp67_ASAP7_75t_SL g2272 ( 
.A(n_2209),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2259),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2122),
.B(n_891),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2133),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2213),
.B(n_955),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2240),
.Y(n_2277)
);

NAND2x1p5_ASAP7_75t_L g2278 ( 
.A(n_2243),
.B(n_1580),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2244),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2179),
.B(n_959),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2246),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_2148),
.Y(n_2282)
);

NAND2x1p5_ASAP7_75t_L g2283 ( 
.A(n_2253),
.B(n_1589),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2126),
.B(n_963),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2154),
.B(n_967),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2268),
.B(n_1725),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2135),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2174),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_2202),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2145),
.B(n_968),
.Y(n_2290)
);

NOR2x1_ASAP7_75t_L g2291 ( 
.A(n_2120),
.B(n_2),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2203),
.B(n_3),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2207),
.Y(n_2293)
);

INVxp67_ASAP7_75t_L g2294 ( 
.A(n_2208),
.Y(n_2294)
);

AOI21xp33_ASAP7_75t_SL g2295 ( 
.A1(n_2230),
.A2(n_974),
.B(n_972),
.Y(n_2295)
);

NAND2x1_ASAP7_75t_L g2296 ( 
.A(n_2195),
.B(n_1587),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2268),
.B(n_4),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_2219),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2221),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_SL g2300 ( 
.A(n_2234),
.B(n_1587),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_2245),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2242),
.B(n_4),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_2248),
.B(n_2249),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2195),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2256),
.B(n_5),
.Y(n_2305)
);

INVxp67_ASAP7_75t_L g2306 ( 
.A(n_2258),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2266),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2138),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2224),
.B(n_1713),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2176),
.B(n_6),
.Y(n_2310)
);

HB1xp67_ASAP7_75t_L g2311 ( 
.A(n_2131),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2178),
.B(n_2158),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2125),
.Y(n_2313)
);

NAND2xp33_ASAP7_75t_L g2314 ( 
.A(n_2254),
.B(n_1592),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2186),
.B(n_6),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2216),
.B(n_7),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2227),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2144),
.B(n_7),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2265),
.B(n_8),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2163),
.B(n_9),
.Y(n_2320)
);

OR2x2_ASAP7_75t_L g2321 ( 
.A(n_2187),
.B(n_10),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2257),
.B(n_1730),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2140),
.A2(n_756),
.B1(n_1742),
.B2(n_1716),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2142),
.B(n_2198),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2151),
.B(n_11),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2170),
.B(n_2130),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2119),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2167),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2169),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_2238),
.Y(n_2330)
);

NAND3xp33_ASAP7_75t_L g2331 ( 
.A(n_2156),
.B(n_916),
.C(n_915),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2171),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2180),
.B(n_11),
.Y(n_2333)
);

NOR2x1_ASAP7_75t_L g2334 ( 
.A(n_2147),
.B(n_12),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2173),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2177),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2181),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2165),
.B(n_12),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2212),
.B(n_13),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2190),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2152),
.B(n_14),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2200),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2215),
.B(n_2222),
.Y(n_2343)
);

NAND2xp33_ASAP7_75t_L g2344 ( 
.A(n_2157),
.B(n_1592),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2263),
.B(n_14),
.Y(n_2345)
);

OR2x2_ASAP7_75t_L g2346 ( 
.A(n_2155),
.B(n_15),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2192),
.B(n_15),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2223),
.B(n_16),
.Y(n_2348)
);

AOI22x1_ASAP7_75t_SL g2349 ( 
.A1(n_2193),
.A2(n_918),
.B1(n_922),
.B2(n_916),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2223),
.B(n_16),
.Y(n_2350)
);

OR2x2_ASAP7_75t_L g2351 ( 
.A(n_2162),
.B(n_17),
.Y(n_2351)
);

NOR2x1_ASAP7_75t_L g2352 ( 
.A(n_2205),
.B(n_17),
.Y(n_2352)
);

OR2x2_ASAP7_75t_L g2353 ( 
.A(n_2201),
.B(n_19),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2132),
.B(n_19),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2149),
.B(n_20),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2194),
.B(n_20),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2160),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2121),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_L g2359 ( 
.A(n_2157),
.B(n_1592),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2233),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2189),
.B(n_21),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2196),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2262),
.B(n_21),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2197),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2218),
.B(n_22),
.Y(n_2365)
);

INVxp67_ASAP7_75t_L g2366 ( 
.A(n_2204),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2264),
.B(n_22),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2168),
.Y(n_2368)
);

OAI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2123),
.A2(n_2220),
.B(n_2214),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2225),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2136),
.B(n_25),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2264),
.B(n_1732),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2217),
.A2(n_1701),
.B1(n_1702),
.B2(n_1699),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2231),
.B(n_25),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2229),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2206),
.B(n_26),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2166),
.B(n_1732),
.Y(n_2377)
);

NOR2xp67_ASAP7_75t_L g2378 ( 
.A(n_2236),
.B(n_26),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2235),
.B(n_27),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2153),
.B(n_28),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2134),
.B(n_2210),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2129),
.B(n_29),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2232),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2239),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2172),
.B(n_30),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2131),
.B(n_30),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2183),
.B(n_31),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2269),
.B(n_2260),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2291),
.B(n_2161),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2272),
.B(n_2141),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2311),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2275),
.B(n_2191),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2270),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2291),
.B(n_2185),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2273),
.B(n_2237),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2303),
.B(n_2247),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_2289),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2303),
.B(n_2252),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2279),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_2386),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_2294),
.B(n_2298),
.Y(n_2401)
);

INVx1_ASAP7_75t_SL g2402 ( 
.A(n_2345),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2277),
.Y(n_2403)
);

INVx1_ASAP7_75t_SL g2404 ( 
.A(n_2349),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2281),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2304),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2306),
.B(n_2267),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2338),
.B(n_2139),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2288),
.B(n_2124),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2287),
.A2(n_2184),
.B1(n_2159),
.B2(n_2188),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2343),
.B(n_2137),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2342),
.B(n_2128),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2301),
.B(n_2182),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2333),
.B(n_2199),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2285),
.B(n_2146),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2292),
.Y(n_2416)
);

NOR2x1_ASAP7_75t_L g2417 ( 
.A(n_2334),
.B(n_2241),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2330),
.B(n_2127),
.Y(n_2418)
);

INVxp67_ASAP7_75t_L g2419 ( 
.A(n_2297),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2339),
.B(n_2356),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2360),
.A2(n_2250),
.B1(n_2211),
.B2(n_2150),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2321),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2310),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2316),
.B(n_2164),
.Y(n_2424)
);

NOR2x1_ASAP7_75t_L g2425 ( 
.A(n_2334),
.B(n_2326),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2307),
.B(n_2143),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2320),
.Y(n_2427)
);

NAND2xp33_ASAP7_75t_SL g2428 ( 
.A(n_2296),
.B(n_2251),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2341),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2315),
.Y(n_2430)
);

INVxp67_ASAP7_75t_L g2431 ( 
.A(n_2324),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2293),
.B(n_2226),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2302),
.Y(n_2433)
);

INVx3_ASAP7_75t_L g2434 ( 
.A(n_2278),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2346),
.Y(n_2435)
);

NOR2x1_ASAP7_75t_L g2436 ( 
.A(n_2352),
.B(n_2325),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2305),
.Y(n_2437)
);

NOR2x1_ASAP7_75t_L g2438 ( 
.A(n_2352),
.B(n_2175),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2299),
.B(n_32),
.Y(n_2439)
);

INVxp67_ASAP7_75t_L g2440 ( 
.A(n_2300),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2312),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2308),
.B(n_32),
.Y(n_2442)
);

OR2x2_ASAP7_75t_L g2443 ( 
.A(n_2351),
.B(n_33),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2319),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_2361),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2290),
.B(n_33),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2353),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2365),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2378),
.B(n_34),
.Y(n_2449)
);

AOI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2385),
.A2(n_756),
.B1(n_922),
.B2(n_918),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2318),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2340),
.Y(n_2452)
);

NAND4xp25_ASAP7_75t_L g2453 ( 
.A(n_2282),
.B(n_40),
.C(n_34),
.D(n_37),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2313),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2284),
.Y(n_2455)
);

INVx1_ASAP7_75t_SL g2456 ( 
.A(n_2358),
.Y(n_2456)
);

NOR2x1_ASAP7_75t_L g2457 ( 
.A(n_2331),
.B(n_37),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2371),
.B(n_40),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2317),
.B(n_41),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2347),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2368),
.B(n_41),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2271),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2366),
.B(n_42),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2376),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2379),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2354),
.B(n_43),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2357),
.B(n_44),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2283),
.Y(n_2468)
);

NAND3xp33_ASAP7_75t_L g2469 ( 
.A(n_2328),
.B(n_937),
.C(n_929),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2329),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2327),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_L g2472 ( 
.A(n_2370),
.B(n_45),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2332),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2335),
.Y(n_2474)
);

INVx2_ASAP7_75t_SL g2475 ( 
.A(n_2362),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2387),
.B(n_45),
.Y(n_2476)
);

INVxp67_ASAP7_75t_L g2477 ( 
.A(n_2355),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2369),
.B(n_756),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2280),
.B(n_46),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2295),
.B(n_46),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2295),
.B(n_47),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2375),
.B(n_49),
.Y(n_2482)
);

NOR2x1_ASAP7_75t_L g2483 ( 
.A(n_2274),
.B(n_50),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2336),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2383),
.B(n_51),
.Y(n_2485)
);

NAND2x1p5_ASAP7_75t_L g2486 ( 
.A(n_2364),
.B(n_1688),
.Y(n_2486)
);

CKINVDCx16_ASAP7_75t_R g2487 ( 
.A(n_2374),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_2384),
.B(n_52),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2337),
.Y(n_2489)
);

OAI221xp5_ASAP7_75t_SL g2490 ( 
.A1(n_2381),
.A2(n_1742),
.B1(n_1778),
.B2(n_1732),
.C(n_55),
.Y(n_2490)
);

OAI21xp5_ASAP7_75t_SL g2491 ( 
.A1(n_2348),
.A2(n_1655),
.B(n_53),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2363),
.B(n_54),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2276),
.B(n_54),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2350),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2367),
.B(n_55),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2380),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2382),
.B(n_57),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2314),
.B(n_57),
.Y(n_2498)
);

INVxp33_ASAP7_75t_L g2499 ( 
.A(n_2309),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2286),
.B(n_58),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2372),
.B(n_58),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_L g2502 ( 
.A(n_2344),
.B(n_59),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_2359),
.B(n_61),
.Y(n_2503)
);

INVx1_ASAP7_75t_SL g2504 ( 
.A(n_2377),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2323),
.B(n_2373),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2322),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2311),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2270),
.B(n_61),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2269),
.Y(n_2509)
);

AOI22xp33_ASAP7_75t_SL g2510 ( 
.A1(n_2272),
.A2(n_1596),
.B1(n_756),
.B2(n_1742),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2272),
.B(n_62),
.Y(n_2511)
);

NOR2x1_ASAP7_75t_L g2512 ( 
.A(n_2291),
.B(n_63),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2269),
.B(n_64),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2269),
.B(n_64),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2270),
.Y(n_2515)
);

INVx1_ASAP7_75t_SL g2516 ( 
.A(n_2270),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2270),
.B(n_65),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2273),
.B(n_66),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2269),
.Y(n_2519)
);

CKINVDCx14_ASAP7_75t_R g2520 ( 
.A(n_2345),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2273),
.B(n_67),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2269),
.B(n_68),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2269),
.B(n_68),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2270),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2270),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2270),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2270),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2270),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2269),
.Y(n_2529)
);

INVx1_ASAP7_75t_SL g2530 ( 
.A(n_2270),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2269),
.B(n_69),
.Y(n_2531)
);

OAI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2291),
.A2(n_1699),
.B1(n_1702),
.B2(n_1701),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2270),
.Y(n_2533)
);

NOR3xp33_ASAP7_75t_SL g2534 ( 
.A(n_2270),
.B(n_937),
.C(n_929),
.Y(n_2534)
);

OAI211xp5_ASAP7_75t_L g2535 ( 
.A1(n_2291),
.A2(n_945),
.B(n_947),
.C(n_938),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2272),
.B(n_69),
.Y(n_2536)
);

NAND4xp25_ASAP7_75t_L g2537 ( 
.A(n_2401),
.B(n_1655),
.C(n_73),
.D(n_70),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2391),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2520),
.B(n_71),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2507),
.Y(n_2540)
);

NAND4xp25_ASAP7_75t_L g2541 ( 
.A(n_2402),
.B(n_75),
.C(n_71),
.D(n_74),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2389),
.A2(n_945),
.B(n_938),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2516),
.B(n_74),
.Y(n_2543)
);

O2A1O1Ixp33_ASAP7_75t_L g2544 ( 
.A1(n_2512),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2544)
);

OAI21xp33_ASAP7_75t_L g2545 ( 
.A1(n_2530),
.A2(n_2456),
.B(n_2499),
.Y(n_2545)
);

NOR2x1_ASAP7_75t_L g2546 ( 
.A(n_2535),
.B(n_77),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2516),
.B(n_2511),
.Y(n_2547)
);

O2A1O1Ixp33_ASAP7_75t_L g2548 ( 
.A1(n_2491),
.A2(n_81),
.B(n_78),
.C(n_79),
.Y(n_2548)
);

NOR3xp33_ASAP7_75t_L g2549 ( 
.A(n_2487),
.B(n_947),
.C(n_690),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2536),
.B(n_78),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_L g2551 ( 
.A(n_2425),
.B(n_693),
.C(n_689),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2397),
.B(n_79),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_2400),
.Y(n_2553)
);

NOR3xp33_ASAP7_75t_L g2554 ( 
.A(n_2398),
.B(n_713),
.C(n_701),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2393),
.A2(n_756),
.B1(n_1737),
.B2(n_1733),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2420),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2508),
.Y(n_2557)
);

AOI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2532),
.A2(n_725),
.B1(n_729),
.B2(n_717),
.C(n_715),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2411),
.B(n_82),
.Y(n_2559)
);

AOI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2394),
.A2(n_740),
.B(n_733),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2417),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2408),
.B(n_83),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2404),
.B(n_2445),
.Y(n_2563)
);

NOR3xp33_ASAP7_75t_L g2564 ( 
.A(n_2431),
.B(n_766),
.C(n_760),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2517),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2406),
.B(n_83),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2459),
.B(n_84),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2509),
.B(n_84),
.Y(n_2568)
);

NOR2xp67_ASAP7_75t_L g2569 ( 
.A(n_2434),
.B(n_85),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2515),
.B(n_85),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2519),
.B(n_86),
.Y(n_2571)
);

NAND2x1p5_ASAP7_75t_L g2572 ( 
.A(n_2436),
.B(n_1666),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2529),
.B(n_87),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2470),
.Y(n_2574)
);

INVx2_ASAP7_75t_SL g2575 ( 
.A(n_2483),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2524),
.A2(n_756),
.B1(n_1737),
.B2(n_1733),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2482),
.B(n_2485),
.Y(n_2577)
);

INVx1_ASAP7_75t_SL g2578 ( 
.A(n_2443),
.Y(n_2578)
);

INVxp33_ASAP7_75t_L g2579 ( 
.A(n_2407),
.Y(n_2579)
);

NAND3xp33_ASAP7_75t_L g2580 ( 
.A(n_2413),
.B(n_783),
.C(n_781),
.Y(n_2580)
);

AOI211xp5_ASAP7_75t_SL g2581 ( 
.A1(n_2419),
.A2(n_2440),
.B(n_2396),
.C(n_2399),
.Y(n_2581)
);

AOI211xp5_ASAP7_75t_L g2582 ( 
.A1(n_2491),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_2582)
);

NAND3xp33_ASAP7_75t_L g2583 ( 
.A(n_2525),
.B(n_785),
.C(n_784),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_SL g2584 ( 
.A(n_2453),
.B(n_583),
.Y(n_2584)
);

NAND3xp33_ASAP7_75t_L g2585 ( 
.A(n_2526),
.B(n_787),
.C(n_786),
.Y(n_2585)
);

AOI221xp5_ASAP7_75t_L g2586 ( 
.A1(n_2421),
.A2(n_813),
.B1(n_820),
.B2(n_797),
.C(n_792),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2461),
.B(n_89),
.Y(n_2587)
);

AOI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2478),
.A2(n_826),
.B(n_824),
.Y(n_2588)
);

NOR3xp33_ASAP7_75t_L g2589 ( 
.A(n_2527),
.B(n_836),
.C(n_828),
.Y(n_2589)
);

AOI211xp5_ASAP7_75t_L g2590 ( 
.A1(n_2453),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2467),
.B(n_93),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_2534),
.Y(n_2592)
);

OAI21xp33_ASAP7_75t_L g2593 ( 
.A1(n_2418),
.A2(n_1737),
.B(n_1733),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2528),
.B(n_94),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2533),
.B(n_95),
.Y(n_2595)
);

NOR3xp33_ASAP7_75t_L g2596 ( 
.A(n_2395),
.B(n_841),
.C(n_838),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2438),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2449),
.Y(n_2598)
);

NAND4xp25_ASAP7_75t_L g2599 ( 
.A(n_2388),
.B(n_97),
.C(n_95),
.D(n_96),
.Y(n_2599)
);

NOR2x1_ASAP7_75t_L g2600 ( 
.A(n_2469),
.B(n_96),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2463),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2427),
.B(n_97),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2518),
.B(n_98),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2521),
.B(n_99),
.Y(n_2604)
);

AO21x1_ASAP7_75t_L g2605 ( 
.A1(n_2428),
.A2(n_99),
.B(n_104),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2416),
.B(n_104),
.Y(n_2606)
);

NAND2xp33_ASAP7_75t_L g2607 ( 
.A(n_2435),
.B(n_855),
.Y(n_2607)
);

AOI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2441),
.A2(n_1740),
.B1(n_1700),
.B2(n_1716),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2429),
.B(n_105),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2493),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2434),
.B(n_2475),
.Y(n_2611)
);

OAI211xp5_ASAP7_75t_L g2612 ( 
.A1(n_2403),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2612)
);

BUFx12f_ASAP7_75t_L g2613 ( 
.A(n_2390),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2422),
.B(n_107),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2412),
.B(n_109),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2500),
.Y(n_2616)
);

NAND4xp25_ASAP7_75t_L g2617 ( 
.A(n_2432),
.B(n_111),
.C(n_109),
.D(n_110),
.Y(n_2617)
);

AOI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2415),
.A2(n_874),
.B(n_861),
.Y(n_2618)
);

OAI21xp33_ASAP7_75t_L g2619 ( 
.A1(n_2477),
.A2(n_1740),
.B(n_1695),
.Y(n_2619)
);

OAI21xp33_ASAP7_75t_SL g2620 ( 
.A1(n_2506),
.A2(n_1695),
.B(n_1729),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2426),
.B(n_110),
.Y(n_2621)
);

NOR2x1_ASAP7_75t_L g2622 ( 
.A(n_2469),
.B(n_111),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2513),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2405),
.B(n_112),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2569),
.Y(n_2625)
);

OAI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2611),
.A2(n_2410),
.B(n_2504),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_SL g2627 ( 
.A(n_2545),
.B(n_2392),
.C(n_2424),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2563),
.A2(n_2553),
.B1(n_2613),
.B2(n_2539),
.Y(n_2628)
);

AOI211x1_ASAP7_75t_L g2629 ( 
.A1(n_2605),
.A2(n_2452),
.B(n_2473),
.C(n_2454),
.Y(n_2629)
);

A2O1A1Ixp33_ASAP7_75t_L g2630 ( 
.A1(n_2544),
.A2(n_2502),
.B(n_2503),
.C(n_2501),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2575),
.B(n_2514),
.Y(n_2631)
);

AOI211xp5_ASAP7_75t_SL g2632 ( 
.A1(n_2597),
.A2(n_2409),
.B(n_2494),
.C(n_2423),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2584),
.A2(n_2447),
.B1(n_2448),
.B2(n_2430),
.Y(n_2633)
);

XNOR2xp5_ASAP7_75t_L g2634 ( 
.A(n_2592),
.B(n_2444),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2556),
.A2(n_2496),
.B1(n_2464),
.B2(n_2465),
.Y(n_2635)
);

AOI222xp33_ASAP7_75t_L g2636 ( 
.A1(n_2561),
.A2(n_2474),
.B1(n_2489),
.B2(n_2484),
.C1(n_2433),
.C2(n_2437),
.Y(n_2636)
);

OAI211xp5_ASAP7_75t_L g2637 ( 
.A1(n_2582),
.A2(n_2510),
.B(n_2523),
.C(n_2522),
.Y(n_2637)
);

AOI221x1_ASAP7_75t_L g2638 ( 
.A1(n_2538),
.A2(n_2531),
.B1(n_2439),
.B2(n_2442),
.C(n_2451),
.Y(n_2638)
);

A2O1A1Ixp33_ASAP7_75t_L g2639 ( 
.A1(n_2548),
.A2(n_2488),
.B(n_2472),
.C(n_2490),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2559),
.B(n_2460),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2543),
.B(n_2446),
.Y(n_2641)
);

AOI221xp5_ASAP7_75t_L g2642 ( 
.A1(n_2540),
.A2(n_2468),
.B1(n_2462),
.B2(n_2455),
.C(n_2505),
.Y(n_2642)
);

AOI222xp33_ASAP7_75t_L g2643 ( 
.A1(n_2574),
.A2(n_2471),
.B1(n_2495),
.B2(n_2457),
.C1(n_2480),
.C2(n_2481),
.Y(n_2643)
);

XNOR2x1_ASAP7_75t_L g2644 ( 
.A(n_2621),
.B(n_2414),
.Y(n_2644)
);

AOI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2547),
.A2(n_2607),
.B(n_2577),
.Y(n_2645)
);

AOI211xp5_ASAP7_75t_L g2646 ( 
.A1(n_2579),
.A2(n_2498),
.B(n_2497),
.C(n_2466),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2590),
.B(n_2458),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2578),
.Y(n_2648)
);

AOI221x1_ASAP7_75t_L g2649 ( 
.A1(n_2599),
.A2(n_2476),
.B1(n_2492),
.B2(n_2479),
.C(n_2450),
.Y(n_2649)
);

AOI322xp5_ASAP7_75t_L g2650 ( 
.A1(n_2601),
.A2(n_2450),
.A3(n_2486),
.B1(n_1740),
.B2(n_118),
.C1(n_120),
.C2(n_121),
.Y(n_2650)
);

O2A1O1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2582),
.A2(n_117),
.B(n_113),
.C(n_116),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_R g2652 ( 
.A(n_2557),
.B(n_116),
.Y(n_2652)
);

A2O1A1Ixp33_ASAP7_75t_L g2653 ( 
.A1(n_2590),
.A2(n_124),
.B(n_118),
.C(n_122),
.Y(n_2653)
);

OAI222xp33_ASAP7_75t_L g2654 ( 
.A1(n_2565),
.A2(n_1654),
.B1(n_126),
.B2(n_128),
.C1(n_122),
.C2(n_125),
.Y(n_2654)
);

NAND4xp25_ASAP7_75t_L g2655 ( 
.A(n_2581),
.B(n_127),
.C(n_125),
.D(n_126),
.Y(n_2655)
);

OAI211xp5_ASAP7_75t_SL g2656 ( 
.A1(n_2586),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2541),
.B(n_129),
.Y(n_2657)
);

AOI221xp5_ASAP7_75t_L g2658 ( 
.A1(n_2552),
.A2(n_879),
.B1(n_886),
.B2(n_877),
.C(n_876),
.Y(n_2658)
);

AOI221xp5_ASAP7_75t_L g2659 ( 
.A1(n_2580),
.A2(n_892),
.B1(n_961),
.B2(n_889),
.C(n_888),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2562),
.Y(n_2660)
);

OAI321xp33_ASAP7_75t_L g2661 ( 
.A1(n_2598),
.A2(n_132),
.A3(n_133),
.B1(n_134),
.B2(n_135),
.C(n_136),
.Y(n_2661)
);

A2O1A1Ixp33_ASAP7_75t_L g2662 ( 
.A1(n_2594),
.A2(n_2595),
.B(n_2606),
.C(n_2612),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2615),
.Y(n_2663)
);

OAI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2614),
.A2(n_1674),
.B(n_1679),
.Y(n_2664)
);

OAI31xp33_ASAP7_75t_L g2665 ( 
.A1(n_2537),
.A2(n_136),
.A3(n_133),
.B(n_134),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2550),
.Y(n_2666)
);

NOR3xp33_ASAP7_75t_SL g2667 ( 
.A(n_2617),
.B(n_2623),
.C(n_2571),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2616),
.A2(n_1700),
.B1(n_1716),
.B2(n_1727),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2566),
.B(n_138),
.Y(n_2669)
);

AOI221x1_ASAP7_75t_L g2670 ( 
.A1(n_2549),
.A2(n_142),
.B1(n_138),
.B2(n_139),
.C(n_143),
.Y(n_2670)
);

AOI221xp5_ASAP7_75t_L g2671 ( 
.A1(n_2589),
.A2(n_2554),
.B1(n_2596),
.B2(n_2564),
.C(n_2610),
.Y(n_2671)
);

OAI21xp5_ASAP7_75t_SL g2672 ( 
.A1(n_2570),
.A2(n_139),
.B(n_145),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2572),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2567),
.A2(n_1727),
.B1(n_1734),
.B2(n_1700),
.Y(n_2674)
);

AOI221xp5_ASAP7_75t_L g2675 ( 
.A1(n_2624),
.A2(n_973),
.B1(n_966),
.B2(n_964),
.C(n_148),
.Y(n_2675)
);

NAND4xp25_ASAP7_75t_L g2676 ( 
.A(n_2546),
.B(n_148),
.C(n_145),
.D(n_146),
.Y(n_2676)
);

OAI221xp5_ASAP7_75t_SL g2677 ( 
.A1(n_2620),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.C(n_153),
.Y(n_2677)
);

AOI221xp5_ASAP7_75t_L g2678 ( 
.A1(n_2568),
.A2(n_154),
.B1(n_150),
.B2(n_152),
.C(n_156),
.Y(n_2678)
);

OAI211xp5_ASAP7_75t_SL g2679 ( 
.A1(n_2558),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_2679)
);

NAND5xp2_ASAP7_75t_L g2680 ( 
.A(n_2555),
.B(n_160),
.C(n_157),
.D(n_159),
.E(n_161),
.Y(n_2680)
);

OAI31xp33_ASAP7_75t_L g2681 ( 
.A1(n_2573),
.A2(n_161),
.A3(n_159),
.B(n_160),
.Y(n_2681)
);

AOI221xp5_ASAP7_75t_L g2682 ( 
.A1(n_2609),
.A2(n_167),
.B1(n_162),
.B2(n_165),
.C(n_168),
.Y(n_2682)
);

AOI211x1_ASAP7_75t_L g2683 ( 
.A1(n_2626),
.A2(n_2551),
.B(n_2585),
.C(n_2583),
.Y(n_2683)
);

OAI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2628),
.A2(n_2591),
.B1(n_2587),
.B2(n_2602),
.Y(n_2684)
);

AOI221xp5_ASAP7_75t_L g2685 ( 
.A1(n_2629),
.A2(n_2603),
.B1(n_2604),
.B2(n_2542),
.C(n_2593),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2655),
.B(n_2600),
.Y(n_2686)
);

NOR3xp33_ASAP7_75t_L g2687 ( 
.A(n_2642),
.B(n_2622),
.C(n_2560),
.Y(n_2687)
);

OAI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2665),
.A2(n_2576),
.B1(n_2619),
.B2(n_2618),
.C(n_2588),
.Y(n_2688)
);

AOI21xp33_ASAP7_75t_SL g2689 ( 
.A1(n_2644),
.A2(n_162),
.B(n_165),
.Y(n_2689)
);

NAND4xp75_ASAP7_75t_L g2690 ( 
.A(n_2638),
.B(n_2608),
.C(n_169),
.D(n_167),
.Y(n_2690)
);

NAND3xp33_ASAP7_75t_L g2691 ( 
.A(n_2636),
.B(n_168),
.C(n_170),
.Y(n_2691)
);

OAI21xp5_ASAP7_75t_SL g2692 ( 
.A1(n_2632),
.A2(n_170),
.B(n_173),
.Y(n_2692)
);

NOR2x1_ASAP7_75t_L g2693 ( 
.A(n_2676),
.B(n_173),
.Y(n_2693)
);

AOI21xp33_ASAP7_75t_SL g2694 ( 
.A1(n_2625),
.A2(n_174),
.B(n_175),
.Y(n_2694)
);

AOI211x1_ASAP7_75t_L g2695 ( 
.A1(n_2637),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_2695)
);

NOR4xp25_ASAP7_75t_L g2696 ( 
.A(n_2662),
.B(n_178),
.C(n_176),
.D(n_177),
.Y(n_2696)
);

AOI211x1_ASAP7_75t_L g2697 ( 
.A1(n_2631),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2697)
);

AOI322xp5_ASAP7_75t_L g2698 ( 
.A1(n_2627),
.A2(n_179),
.A3(n_180),
.B1(n_181),
.B2(n_182),
.C1(n_183),
.C2(n_184),
.Y(n_2698)
);

OA22x2_ASAP7_75t_L g2699 ( 
.A1(n_2633),
.A2(n_184),
.B1(n_180),
.B2(n_183),
.Y(n_2699)
);

OAI21xp33_ASAP7_75t_SL g2700 ( 
.A1(n_2643),
.A2(n_185),
.B(n_186),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2648),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2663),
.B(n_187),
.Y(n_2702)
);

AOI221xp5_ASAP7_75t_L g2703 ( 
.A1(n_2677),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_2703)
);

OAI211xp5_ASAP7_75t_L g2704 ( 
.A1(n_2650),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_2704)
);

OAI21xp33_ASAP7_75t_L g2705 ( 
.A1(n_2634),
.A2(n_1727),
.B(n_1734),
.Y(n_2705)
);

AOI322xp5_ASAP7_75t_L g2706 ( 
.A1(n_2660),
.A2(n_191),
.A3(n_193),
.B1(n_194),
.B2(n_196),
.C1(n_197),
.C2(n_198),
.Y(n_2706)
);

A2O1A1Ixp33_ASAP7_75t_L g2707 ( 
.A1(n_2651),
.A2(n_197),
.B(n_193),
.C(n_194),
.Y(n_2707)
);

NOR4xp25_ASAP7_75t_SL g2708 ( 
.A(n_2672),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_2708)
);

AOI221xp5_ASAP7_75t_SL g2709 ( 
.A1(n_2639),
.A2(n_202),
.B1(n_199),
.B2(n_200),
.C(n_204),
.Y(n_2709)
);

NAND4xp25_ASAP7_75t_L g2710 ( 
.A(n_2649),
.B(n_2646),
.C(n_2635),
.D(n_2630),
.Y(n_2710)
);

NOR2xp33_ASAP7_75t_SL g2711 ( 
.A(n_2681),
.B(n_202),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2669),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2647),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2680),
.B(n_206),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2657),
.A2(n_1673),
.B1(n_1700),
.B2(n_1729),
.Y(n_2715)
);

OAI221xp5_ASAP7_75t_SL g2716 ( 
.A1(n_2645),
.A2(n_206),
.B1(n_208),
.B2(n_210),
.C(n_211),
.Y(n_2716)
);

OAI221xp5_ASAP7_75t_L g2717 ( 
.A1(n_2653),
.A2(n_208),
.B1(n_212),
.B2(n_213),
.C(n_214),
.Y(n_2717)
);

NAND3xp33_ASAP7_75t_L g2718 ( 
.A(n_2667),
.B(n_214),
.C(n_216),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2701),
.B(n_2666),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2693),
.B(n_2640),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2699),
.Y(n_2721)
);

AOI321xp33_ASAP7_75t_L g2722 ( 
.A1(n_2687),
.A2(n_2641),
.A3(n_2673),
.B1(n_2671),
.B2(n_2675),
.C(n_2682),
.Y(n_2722)
);

OAI322xp33_ASAP7_75t_L g2723 ( 
.A1(n_2711),
.A2(n_2674),
.A3(n_2661),
.B1(n_2670),
.B2(n_2656),
.C1(n_2679),
.C2(n_2652),
.Y(n_2723)
);

OAI32xp33_ASAP7_75t_L g2724 ( 
.A1(n_2700),
.A2(n_2654),
.A3(n_2661),
.B1(n_2668),
.B2(n_2678),
.Y(n_2724)
);

OAI22xp5_ASAP7_75t_L g2725 ( 
.A1(n_2718),
.A2(n_2658),
.B1(n_2659),
.B2(n_2664),
.Y(n_2725)
);

AND2x4_ASAP7_75t_L g2726 ( 
.A(n_2702),
.B(n_216),
.Y(n_2726)
);

OAI221xp5_ASAP7_75t_L g2727 ( 
.A1(n_2692),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.C(n_221),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2714),
.Y(n_2728)
);

A2O1A1Ixp33_ASAP7_75t_L g2729 ( 
.A1(n_2698),
.A2(n_223),
.B(n_218),
.C(n_222),
.Y(n_2729)
);

OAI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2710),
.A2(n_1700),
.B1(n_225),
.B2(n_223),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2691),
.Y(n_2731)
);

OAI21xp33_ASAP7_75t_L g2732 ( 
.A1(n_2686),
.A2(n_1729),
.B(n_224),
.Y(n_2732)
);

NOR2x1_ASAP7_75t_L g2733 ( 
.A(n_2690),
.B(n_225),
.Y(n_2733)
);

NOR2x1p5_ASAP7_75t_L g2734 ( 
.A(n_2713),
.B(n_226),
.Y(n_2734)
);

INVxp67_ASAP7_75t_SL g2735 ( 
.A(n_2716),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2689),
.B(n_226),
.Y(n_2736)
);

NAND4xp75_ASAP7_75t_L g2737 ( 
.A(n_2695),
.B(n_229),
.C(n_227),
.D(n_228),
.Y(n_2737)
);

OAI321xp33_ASAP7_75t_L g2738 ( 
.A1(n_2684),
.A2(n_227),
.A3(n_228),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_2738)
);

AOI322xp5_ASAP7_75t_L g2739 ( 
.A1(n_2730),
.A2(n_2685),
.A3(n_2712),
.B1(n_2709),
.B2(n_2703),
.C1(n_2707),
.C2(n_2705),
.Y(n_2739)
);

NAND3xp33_ASAP7_75t_SL g2740 ( 
.A(n_2729),
.B(n_2708),
.C(n_2696),
.Y(n_2740)
);

OR2x2_ASAP7_75t_L g2741 ( 
.A(n_2721),
.B(n_2704),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2720),
.B(n_2694),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2737),
.Y(n_2743)
);

NOR3xp33_ASAP7_75t_L g2744 ( 
.A(n_2728),
.B(n_2717),
.C(n_2688),
.Y(n_2744)
);

CKINVDCx14_ASAP7_75t_R g2745 ( 
.A(n_2719),
.Y(n_2745)
);

OR3x2_ASAP7_75t_L g2746 ( 
.A(n_2731),
.B(n_2683),
.C(n_2697),
.Y(n_2746)
);

AND3x4_ASAP7_75t_L g2747 ( 
.A(n_2733),
.B(n_2726),
.C(n_2723),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2738),
.B(n_2706),
.Y(n_2748)
);

NAND4xp25_ASAP7_75t_L g2749 ( 
.A(n_2722),
.B(n_2715),
.C(n_235),
.D(n_233),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2734),
.Y(n_2750)
);

NAND4xp75_ASAP7_75t_L g2751 ( 
.A(n_2736),
.B(n_2735),
.C(n_2727),
.D(n_2724),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2726),
.B(n_234),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2732),
.B(n_236),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2725),
.Y(n_2754)
);

AND3x4_ASAP7_75t_L g2755 ( 
.A(n_2733),
.B(n_236),
.C(n_237),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2752),
.Y(n_2756)
);

OAI211xp5_ASAP7_75t_SL g2757 ( 
.A1(n_2739),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2755),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2746),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2745),
.B(n_239),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_R g2761 ( 
.A(n_2740),
.B(n_241),
.Y(n_2761)
);

OAI221xp5_ASAP7_75t_SL g2762 ( 
.A1(n_2741),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.C(n_245),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_SL g2763 ( 
.A1(n_2743),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2742),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2750),
.Y(n_2765)
);

CKINVDCx16_ASAP7_75t_R g2766 ( 
.A(n_2754),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2744),
.B(n_247),
.Y(n_2767)
);

INVxp67_ASAP7_75t_SL g2768 ( 
.A(n_2753),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2748),
.B(n_248),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2747),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2751),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_2749),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_2745),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_2745),
.Y(n_2774)
);

NOR2xp67_ASAP7_75t_SL g2775 ( 
.A(n_2774),
.B(n_249),
.Y(n_2775)
);

OR2x2_ASAP7_75t_L g2776 ( 
.A(n_2760),
.B(n_2769),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2773),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2756),
.Y(n_2778)
);

AO21x1_ASAP7_75t_L g2779 ( 
.A1(n_2767),
.A2(n_249),
.B(n_250),
.Y(n_2779)
);

INVx4_ASAP7_75t_L g2780 ( 
.A(n_2766),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2758),
.Y(n_2781)
);

AOI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2770),
.A2(n_1673),
.B1(n_254),
.B2(n_251),
.Y(n_2782)
);

AOI22x1_ASAP7_75t_L g2783 ( 
.A1(n_2771),
.A2(n_256),
.B1(n_251),
.B2(n_253),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2764),
.Y(n_2784)
);

AOI22x1_ASAP7_75t_L g2785 ( 
.A1(n_2759),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2765),
.B(n_257),
.Y(n_2786)
);

XNOR2x1_ASAP7_75t_L g2787 ( 
.A(n_2772),
.B(n_258),
.Y(n_2787)
);

AOI22x1_ASAP7_75t_L g2788 ( 
.A1(n_2768),
.A2(n_2757),
.B1(n_2761),
.B2(n_2762),
.Y(n_2788)
);

OAI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2763),
.A2(n_263),
.B1(n_260),
.B2(n_261),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2774),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2773),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2773),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2773),
.A2(n_265),
.B1(n_261),
.B2(n_264),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2774),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2775),
.B(n_264),
.Y(n_2795)
);

INVx4_ASAP7_75t_L g2796 ( 
.A(n_2780),
.Y(n_2796)
);

OAI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2790),
.A2(n_265),
.B(n_267),
.Y(n_2797)
);

AOI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2794),
.A2(n_267),
.B(n_268),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2778),
.B(n_268),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2789),
.B(n_269),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2775),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2786),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2791),
.B(n_269),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2779),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2787),
.Y(n_2805)
);

AO21x1_ASAP7_75t_L g2806 ( 
.A1(n_2784),
.A2(n_270),
.B(n_271),
.Y(n_2806)
);

XNOR2x1_ASAP7_75t_L g2807 ( 
.A(n_2788),
.B(n_270),
.Y(n_2807)
);

AOI21xp5_ASAP7_75t_SL g2808 ( 
.A1(n_2793),
.A2(n_271),
.B(n_272),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2783),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2806),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2803),
.Y(n_2811)
);

INVx3_ASAP7_75t_L g2812 ( 
.A(n_2799),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2795),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2807),
.Y(n_2814)
);

HB1xp67_ASAP7_75t_L g2815 ( 
.A(n_2804),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2801),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2800),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2796),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2797),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2802),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2809),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2805),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2798),
.Y(n_2823)
);

AOI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2820),
.A2(n_2777),
.B1(n_2792),
.B2(n_2781),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2810),
.B(n_2808),
.Y(n_2825)
);

OAI31xp33_ASAP7_75t_L g2826 ( 
.A1(n_2815),
.A2(n_2776),
.A3(n_2785),
.B(n_2782),
.Y(n_2826)
);

OAI21x1_ASAP7_75t_SL g2827 ( 
.A1(n_2818),
.A2(n_272),
.B(n_273),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2816),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2812),
.Y(n_2829)
);

OAI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2821),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2830)
);

OAI22x1_ASAP7_75t_SL g2831 ( 
.A1(n_2814),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_2831)
);

XOR2xp5_ASAP7_75t_L g2832 ( 
.A(n_2822),
.B(n_279),
.Y(n_2832)
);

AOI22x1_ASAP7_75t_L g2833 ( 
.A1(n_2811),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_2833)
);

AOI22x1_ASAP7_75t_L g2834 ( 
.A1(n_2819),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2812),
.Y(n_2835)
);

HB1xp67_ASAP7_75t_L g2836 ( 
.A(n_2823),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2813),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2817),
.Y(n_2838)
);

OAI22x1_ASAP7_75t_L g2839 ( 
.A1(n_2833),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2832),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2829),
.B(n_287),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2835),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_2842)
);

AOI31xp33_ASAP7_75t_L g2843 ( 
.A1(n_2825),
.A2(n_289),
.A3(n_290),
.B(n_291),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2824),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2827),
.Y(n_2845)
);

INVxp67_ASAP7_75t_L g2846 ( 
.A(n_2831),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2838),
.Y(n_2847)
);

AOI221xp5_ASAP7_75t_L g2848 ( 
.A1(n_2836),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.C(n_296),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2837),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_2849)
);

OAI21x1_ASAP7_75t_SL g2850 ( 
.A1(n_2834),
.A2(n_299),
.B(n_300),
.Y(n_2850)
);

NAND4xp25_ASAP7_75t_SL g2851 ( 
.A(n_2847),
.B(n_2826),
.C(n_2830),
.D(n_2828),
.Y(n_2851)
);

AOI221x1_ASAP7_75t_L g2852 ( 
.A1(n_2845),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.C(n_302),
.Y(n_2852)
);

OAI322xp33_ASAP7_75t_L g2853 ( 
.A1(n_2846),
.A2(n_303),
.A3(n_304),
.B1(n_305),
.B2(n_306),
.C1(n_307),
.C2(n_308),
.Y(n_2853)
);

NOR4xp25_ASAP7_75t_L g2854 ( 
.A(n_2840),
.B(n_305),
.C(n_306),
.D(n_307),
.Y(n_2854)
);

AOI211xp5_ASAP7_75t_SL g2855 ( 
.A1(n_2843),
.A2(n_309),
.B(n_310),
.C(n_311),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2841),
.Y(n_2856)
);

AOI22xp33_ASAP7_75t_L g2857 ( 
.A1(n_2850),
.A2(n_309),
.B1(n_310),
.B2(n_312),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2839),
.Y(n_2858)
);

OAI322xp33_ASAP7_75t_L g2859 ( 
.A1(n_2844),
.A2(n_312),
.A3(n_313),
.B1(n_314),
.B2(n_315),
.C1(n_316),
.C2(n_317),
.Y(n_2859)
);

AOI211xp5_ASAP7_75t_L g2860 ( 
.A1(n_2848),
.A2(n_313),
.B(n_314),
.C(n_316),
.Y(n_2860)
);

O2A1O1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2849),
.A2(n_319),
.B(n_320),
.C(n_321),
.Y(n_2861)
);

INVxp67_ASAP7_75t_L g2862 ( 
.A(n_2842),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2858),
.Y(n_2863)
);

AOI222xp33_ASAP7_75t_L g2864 ( 
.A1(n_2862),
.A2(n_321),
.B1(n_322),
.B2(n_324),
.C1(n_325),
.C2(n_326),
.Y(n_2864)
);

AOI21xp33_ASAP7_75t_SL g2865 ( 
.A1(n_2854),
.A2(n_322),
.B(n_325),
.Y(n_2865)
);

INVxp67_ASAP7_75t_L g2866 ( 
.A(n_2851),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2856),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2857),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_2868)
);

OAI222xp33_ASAP7_75t_L g2869 ( 
.A1(n_2861),
.A2(n_2855),
.B1(n_2860),
.B2(n_2859),
.C1(n_2852),
.C2(n_2853),
.Y(n_2869)
);

OAI21xp5_ASAP7_75t_SL g2870 ( 
.A1(n_2855),
.A2(n_332),
.B(n_333),
.Y(n_2870)
);

AOI22xp5_ASAP7_75t_L g2871 ( 
.A1(n_2851),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2870),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_SL g2873 ( 
.A1(n_2866),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_2873)
);

AOI22xp5_ASAP7_75t_SL g2874 ( 
.A1(n_2863),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_2874)
);

OAI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2868),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2873),
.B(n_2865),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2872),
.A2(n_2871),
.B1(n_2867),
.B2(n_2869),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2875),
.B(n_2864),
.Y(n_2878)
);

NOR3xp33_ASAP7_75t_L g2879 ( 
.A(n_2877),
.B(n_2874),
.C(n_343),
.Y(n_2879)
);

AOI211xp5_ASAP7_75t_L g2880 ( 
.A1(n_2879),
.A2(n_2876),
.B(n_2878),
.C(n_345),
.Y(n_2880)
);


endmodule