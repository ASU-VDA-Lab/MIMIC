module fake_jpeg_16669_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_72),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_66),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_57),
.B(n_64),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_5),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_68),
.Y(n_93)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_14),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_40),
.B1(n_30),
.B2(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_75),
.A2(n_96),
.B1(n_109),
.B2(n_126),
.Y(n_165)
);

CKINVDCx9p33_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_78),
.B(n_97),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_83),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_19),
.B1(n_36),
.B2(n_26),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_39),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_89),
.B(n_101),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_33),
.B(n_24),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_92),
.B(n_96),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_68),
.B1(n_49),
.B2(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_24),
.C(n_21),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_2),
.C(n_3),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_33),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_113),
.B(n_1),
.Y(n_142)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_108),
.B(n_4),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_37),
.B1(n_39),
.B2(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_16),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_113),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_121),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_0),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_16),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g121 ( 
.A(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_18),
.B1(n_26),
.B2(n_19),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_129),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_154),
.B1(n_142),
.B2(n_134),
.Y(n_199)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_135),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_9),
.B1(n_13),
.B2(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_158),
.B1(n_150),
.B2(n_144),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_24),
.Y(n_140)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_35),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_169),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_2),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_150),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_132),
.B1(n_148),
.B2(n_149),
.Y(n_200)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_3),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_157),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_4),
.B1(n_114),
.B2(n_86),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_120),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_4),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_126),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_100),
.B(n_99),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_105),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_114),
.B1(n_80),
.B2(n_86),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_181),
.B1(n_192),
.B2(n_199),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_90),
.B1(n_102),
.B2(n_80),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_180),
.A2(n_185),
.B1(n_193),
.B2(n_152),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_197),
.B(n_159),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_102),
.B1(n_116),
.B2(n_106),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_77),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_189),
.B(n_201),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_133),
.A2(n_125),
.A3(n_107),
.B1(n_124),
.B2(n_123),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_152),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_123),
.B1(n_124),
.B2(n_94),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_91),
.B1(n_94),
.B2(n_139),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_91),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_180),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_147),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_143),
.A2(n_147),
.B1(n_156),
.B2(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_175),
.B1(n_197),
.B2(n_174),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_153),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_128),
.C(n_145),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_212),
.C(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_176),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_136),
.C(n_131),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_135),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_146),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_226),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_235),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_221),
.B(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_148),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_200),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_166),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_205),
.B(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_163),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_223),
.B(n_227),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_196),
.B(n_138),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_231),
.B1(n_186),
.B2(n_187),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_188),
.B(n_184),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_187),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_174),
.C(n_207),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_236),
.C(n_183),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_175),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_206),
.B1(n_181),
.B2(n_175),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_217),
.B(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_194),
.B1(n_195),
.B2(n_190),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_203),
.B1(n_186),
.B2(n_179),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_248),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_251),
.B1(n_243),
.B2(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_173),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_222),
.B(n_216),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_218),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_229),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_234),
.C(n_210),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_260),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_223),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_179),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_277),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_268),
.C(n_272),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_217),
.B(n_224),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_279),
.B(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_212),
.C(n_214),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_226),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_247),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_247),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_221),
.B(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_240),
.B1(n_227),
.B2(n_242),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_219),
.B(n_237),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_242),
.B1(n_262),
.B2(n_261),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_285),
.B1(n_289),
.B2(n_292),
.Y(n_307)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_242),
.B1(n_237),
.B2(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

AOI221xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_250),
.B1(n_253),
.B2(n_240),
.C(n_244),
.Y(n_290)
);

XOR2x2_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_250),
.B(n_258),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_279),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_255),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_272),
.C(n_267),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_245),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_265),
.B1(n_254),
.B2(n_256),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_300),
.B1(n_301),
.B2(n_239),
.Y(n_309)
);

OAI31xp33_ASAP7_75t_L g314 ( 
.A1(n_297),
.A2(n_283),
.A3(n_270),
.B(n_285),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_256),
.B1(n_248),
.B2(n_275),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_275),
.B1(n_239),
.B2(n_273),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_304),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_268),
.C(n_245),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_314),
.B1(n_315),
.B2(n_307),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_270),
.B(n_305),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_263),
.B(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_266),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_313),
.C(n_232),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_293),
.B(n_286),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_273),
.B(n_266),
.C(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_318),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_282),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_319),
.C(n_320),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_303),
.A3(n_302),
.B1(n_299),
.B2(n_304),
.C1(n_228),
.C2(n_232),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_318),
.A2(n_312),
.B(n_308),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_318),
.B1(n_315),
.B2(n_317),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_324),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_202),
.CI(n_322),
.CON(n_325),
.SN(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_325),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_325),
.Y(n_328)
);


endmodule