module fake_jpeg_3176_n_124 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_51),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_37),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_44),
.C(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_71),
.B1(n_72),
.B2(n_62),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_35),
.B1(n_1),
.B2(n_3),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_4),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_32),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_54),
.B1(n_52),
.B2(n_56),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_78),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_59),
.C(n_58),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_6),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_10),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_18),
.C(n_19),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_67),
.B(n_12),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_73),
.Y(n_99)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_11),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_13),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_26),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_107),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_20),
.B(n_21),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_106),
.B(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_85),
.C(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_112),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_92),
.B(n_27),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_104),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_111),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_110),
.B(n_101),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_107),
.C(n_111),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_115),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_100),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_108),
.Y(n_124)
);


endmodule