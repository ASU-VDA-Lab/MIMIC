module fake_jpeg_6893_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_27),
.B1(n_18),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_68),
.B1(n_69),
.B2(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_23),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_32),
.B(n_31),
.C(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_18),
.B1(n_27),
.B2(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_32),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_19),
.B1(n_34),
.B2(n_29),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_82),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_49),
.B1(n_21),
.B2(n_22),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_67),
.B1(n_53),
.B2(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_86),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_42),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_62),
.CI(n_46),
.CON(n_106),
.SN(n_106)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_37),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_36),
.B1(n_31),
.B2(n_21),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_64),
.B1(n_52),
.B2(n_50),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_36),
.B1(n_42),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_89),
.B1(n_49),
.B2(n_50),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_42),
.B1(n_34),
.B2(n_29),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_99),
.B1(n_107),
.B2(n_109),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_114),
.B1(n_87),
.B2(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_66),
.B1(n_51),
.B2(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_101),
.B(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_105),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_83),
.B1(n_85),
.B2(n_79),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_80),
.B(n_87),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_46),
.B1(n_45),
.B2(n_29),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_46),
.B1(n_29),
.B2(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_45),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_118),
.A2(n_137),
.B1(n_101),
.B2(n_106),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_123),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_87),
.B(n_89),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_83),
.B1(n_87),
.B2(n_85),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_42),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_139),
.B(n_97),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_88),
.B(n_28),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_135),
.Y(n_160)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_93),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_88),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_70),
.B1(n_19),
.B2(n_91),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_70),
.B(n_54),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_0),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_91),
.B1(n_54),
.B2(n_28),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_98),
.B1(n_97),
.B2(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_108),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_94),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_116),
.C(n_111),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_168),
.C(n_25),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_135),
.B1(n_117),
.B2(n_126),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_25),
.B(n_26),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_161),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_131),
.B1(n_132),
.B2(n_130),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_106),
.C(n_28),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_25),
.B1(n_26),
.B2(n_3),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_118),
.B1(n_123),
.B2(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_186),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_182),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_177),
.B1(n_183),
.B2(n_156),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_131),
.B(n_127),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_143),
.Y(n_201)
);

OAI22x1_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_131),
.B1(n_126),
.B2(n_122),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_143),
.B1(n_154),
.B2(n_160),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_146),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_194),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_144),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_25),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_168),
.C(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_144),
.B1(n_154),
.B2(n_163),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_189),
.B1(n_26),
.B2(n_4),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_1),
.B(n_2),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_191),
.C(n_180),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_215),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_159),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_145),
.C(n_155),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_25),
.C(n_26),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_26),
.C(n_2),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_185),
.B1(n_187),
.B2(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_175),
.B1(n_188),
.B2(n_172),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_172),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_232),
.B(n_234),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_190),
.B1(n_176),
.B2(n_174),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_174),
.C(n_171),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_195),
.C(n_200),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_5),
.B(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_214),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_204),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_238),
.C(n_246),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_205),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_237),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_201),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_1),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_233),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_1),
.CI(n_4),
.CON(n_244),
.SN(n_244)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_244),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_248),
.B(n_228),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_5),
.C(n_6),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_5),
.C(n_6),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_259),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_230),
.B(n_247),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_253),
.B(n_255),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_258),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_222),
.B1(n_231),
.B2(n_225),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_241),
.B1(n_248),
.B2(n_235),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_227),
.C(n_219),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_227),
.C(n_226),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_9),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_242),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_267),
.B(n_12),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_10),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_7),
.B(n_9),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_10),
.B(n_11),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_251),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_275),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_249),
.C(n_11),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_272),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_10),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_276),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_280),
.B(n_273),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_262),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_265),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_12),
.B(n_13),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.C(n_12),
.Y(n_285)
);

OAI21x1_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_13),
.B(n_14),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_277),
.C(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_15),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_16),
.B(n_279),
.Y(n_290)
);


endmodule