module fake_jpeg_7741_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_20),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_33),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_25),
.B1(n_14),
.B2(n_28),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_34),
.B(n_12),
.C(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_11),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_19),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_14),
.B1(n_12),
.B2(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_30),
.B(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_13),
.C(n_9),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.C(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_35),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_56),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_49),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_55),
.C(n_56),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_61),
.B(n_63),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_27),
.A3(n_14),
.B1(n_35),
.B2(n_26),
.C1(n_8),
.C2(n_13),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_47),
.C(n_27),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_48),
.B(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_57),
.B1(n_35),
.B2(n_52),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_61),
.C(n_62),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_25),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_1),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_26),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_2),
.B(n_4),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_4),
.B(n_5),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.C(n_5),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_6),
.CI(n_7),
.CON(n_77),
.SN(n_77)
);


endmodule