module fake_jpeg_8518_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_24),
.B1(n_32),
.B2(n_29),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_46),
.B1(n_59),
.B2(n_32),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_24),
.B1(n_28),
.B2(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_39),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_24),
.B1(n_28),
.B2(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_27),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_26),
.CON(n_63),
.SN(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_28),
.B(n_16),
.C(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_71),
.Y(n_103)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_88),
.B1(n_32),
.B2(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_31),
.B(n_25),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_39),
.B1(n_40),
.B2(n_37),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_93),
.B1(n_56),
.B2(n_53),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_85),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_47),
.B(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_27),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_19),
.C(n_33),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_23),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_39),
.B1(n_40),
.B2(n_37),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_104),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_116),
.B1(n_117),
.B2(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_35),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_118),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_0),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_68),
.B(n_31),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_53),
.B1(n_45),
.B2(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_40),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_119),
.B(n_17),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_93),
.B1(n_88),
.B2(n_79),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_142),
.B1(n_106),
.B2(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_127),
.A2(n_131),
.B(n_132),
.Y(n_180)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_81),
.B1(n_98),
.B2(n_32),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_92),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_93),
.B(n_112),
.C(n_100),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_136),
.Y(n_158)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_69),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_81),
.B1(n_84),
.B2(n_71),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_146),
.Y(n_179)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_81),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_154),
.B1(n_161),
.B2(n_168),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_114),
.B1(n_95),
.B2(n_111),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_95),
.C(n_106),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_159),
.A2(n_172),
.B(n_173),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_119),
.C(n_102),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_87),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_20),
.C(n_67),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_132),
.B1(n_142),
.B2(n_127),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_126),
.A2(n_98),
.B1(n_99),
.B2(n_17),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_31),
.B(n_33),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_33),
.B(n_19),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_17),
.B(n_19),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_73),
.C(n_82),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_181),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_21),
.B1(n_82),
.B2(n_29),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_122),
.B1(n_131),
.B2(n_21),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_20),
.C(n_30),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_125),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_207),
.C(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_204),
.C(n_205),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_148),
.B1(n_146),
.B2(n_129),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_123),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_144),
.B1(n_130),
.B2(n_143),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_144),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_141),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_128),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_171),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_20),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_169),
.B(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_177),
.B(n_30),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_222),
.C(n_223),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_208),
.B(n_206),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_172),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_167),
.C(n_165),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_167),
.C(n_154),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_159),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_173),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_231),
.C(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_171),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_204),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_157),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_157),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_198),
.B1(n_197),
.B2(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_183),
.A2(n_169),
.B1(n_185),
.B2(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_207),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_213),
.C(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_249),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_SL g248 ( 
.A(n_212),
.B(n_208),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_250),
.B(n_21),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

NOR2x1_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_152),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_205),
.B1(n_191),
.B2(n_188),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_253),
.B1(n_164),
.B2(n_178),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_195),
.B1(n_164),
.B2(n_145),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_217),
.Y(n_255)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_215),
.B1(n_228),
.B2(n_216),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_271),
.B1(n_237),
.B2(n_254),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_223),
.C(n_222),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_6),
.C(n_14),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_15),
.C(n_14),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_225),
.C(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_254),
.C(n_240),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_218),
.C(n_226),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_268),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_242),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_15),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_145),
.B1(n_7),
.B2(n_8),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_274),
.B(n_276),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_259),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_245),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_281),
.B1(n_269),
.B2(n_260),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_236),
.B(n_239),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_239),
.C(n_7),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_285),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_284),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_258),
.B(n_256),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_261),
.B1(n_9),
.B2(n_2),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_12),
.C(n_11),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_295),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_256),
.B(n_265),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_294),
.B(n_1),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_261),
.B(n_11),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_0),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g299 ( 
.A(n_297),
.B(n_285),
.Y(n_299)
);

OAI21x1_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_1),
.B(n_2),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_286),
.B(n_272),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_1),
.B(n_3),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_0),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_305),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_304),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_309),
.B1(n_3),
.B2(n_4),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_312),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_1),
.B(n_3),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_3),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_301),
.B1(n_298),
.B2(n_5),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.C(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_313),
.Y(n_317)
);

AO21x1_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_4),
.B(n_5),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_5),
.Y(n_320)
);


endmodule