module fake_netlist_6_1547_n_359 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_92, n_42, n_96, n_8, n_90, n_24, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_95, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_359);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_95;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_359;

wire n_326;
wire n_256;
wire n_209;
wire n_223;
wire n_278;
wire n_341;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_125;
wire n_168;
wire n_297;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_350;
wire n_142;
wire n_143;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_280;
wire n_287;
wire n_353;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_183;
wire n_338;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_352;
wire n_107;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_293;
wire n_334;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_116;
wire n_211;
wire n_175;
wire n_117;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_346;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_251;
wire n_120;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_61),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_69),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_39),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_28),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_13),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_35),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_21),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_48),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_81),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_30),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_33),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_86),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_32),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_31),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_41),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_57),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_5),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_37),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_40),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_54),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_43),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_55),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_46),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_11),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_66),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_59),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_53),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_50),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_0),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_20),
.B(n_19),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_1),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_2),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_3),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_4),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_104),
.A2(n_6),
.B(n_7),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_7),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_23),
.B(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_106),
.B(n_24),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_10),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_10),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_112),
.A2(n_11),
.B(n_12),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_13),
.B(n_14),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_139),
.B(n_15),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_15),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_125),
.A2(n_128),
.B(n_126),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_26),
.B(n_25),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_109),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_164),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_148),
.B(n_143),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_215),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_159),
.Y(n_233)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_152),
.B(n_149),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_177),
.B1(n_169),
.B2(n_183),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_175),
.Y(n_239)
);

NAND2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_193),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_207),
.B(n_180),
.C(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_181),
.Y(n_243)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_212),
.C(n_192),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_181),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_193),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_212),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_176),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_189),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_156),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_182),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_113),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_240),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_171),
.B(n_213),
.C(n_187),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_199),
.B1(n_200),
.B2(n_186),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_204),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_199),
.B1(n_200),
.B2(n_186),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_208),
.B1(n_160),
.B2(n_161),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_250),
.B(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_229),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_254),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_210),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_214),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_116),
.B1(n_117),
.B2(n_114),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_197),
.B(n_196),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_197),
.B(n_201),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_209),
.B(n_205),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_118),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_217),
.B(n_211),
.C(n_236),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_122),
.B(n_120),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_124),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

NAND2x1p5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_184),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_158),
.B(n_140),
.C(n_141),
.Y(n_295)
);

AO21x2_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_277),
.B(n_279),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

AO21x2_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_274),
.B(n_275),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_150),
.B(n_147),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

BUFx4f_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

AO21x2_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_269),
.B(n_278),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AO21x2_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_157),
.B(n_151),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_163),
.B(n_58),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_60),
.B(n_101),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_282),
.B(n_286),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g318 ( 
.A(n_316),
.B(n_307),
.Y(n_318)
);

AO31x2_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_300),
.A3(n_306),
.B(n_296),
.Y(n_319)
);

AO31x2_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_298),
.A3(n_305),
.B(n_303),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

OR2x6_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_49),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_313),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_314),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_65),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

AND2x4_ASAP7_75t_SL g337 ( 
.A(n_332),
.B(n_330),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_333),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_334),
.Y(n_339)
);

AND2x4_ASAP7_75t_SL g340 ( 
.A(n_332),
.B(n_330),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_339),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_342),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_337),
.B1(n_340),
.B2(n_335),
.Y(n_347)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_70),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_351),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_341),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_72),
.B(n_73),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_76),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_357)
);

NOR2x1_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_90),
.Y(n_358)
);

OAI22x1_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_359)
);


endmodule