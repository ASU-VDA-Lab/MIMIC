module real_jpeg_26051_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_1),
.B(n_104),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_51),
.C(n_54),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_151),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_1),
.B(n_82),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_1),
.A2(n_87),
.B1(n_91),
.B2(n_227),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_32),
.B1(n_54),
.B2(n_55),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_3),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_31),
.B1(n_41),
.B2(n_58),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_58),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_7),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_148),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_148),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_148),
.Y(n_288)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_9),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_155),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_155),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_155),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_67),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_67),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_14),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_146),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_146),
.Y(n_220)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_15),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_19),
.B(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_83),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_20),
.A2(n_70),
.B1(n_71),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_20),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_42),
.B2(n_43),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_21),
.A2(n_22),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_44),
.C(n_60),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_33),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_23),
.A2(n_100),
.B1(n_154),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_24),
.A2(n_27),
.B(n_152),
.C(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_25),
.B(n_26),
.C(n_38),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_26),
.A2(n_27),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_L g243 ( 
.A(n_26),
.B(n_49),
.C(n_63),
.Y(n_243)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HAxp5_ASAP7_75t_SL g242 ( 
.A(n_27),
.B(n_151),
.CON(n_242),
.SN(n_242)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_29),
.Y(n_117)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_34),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_35),
.B(n_151),
.Y(n_152)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_38),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_39),
.A2(n_104),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_39),
.A2(n_104),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_39),
.A2(n_104),
.B1(n_161),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_44),
.A2(n_45),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B(n_56),
.Y(n_45)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_46),
.A2(n_53),
.B1(n_203),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_46),
.A2(n_73),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_48),
.A2(n_64),
.B(n_241),
.C(n_243),
.Y(n_240)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_49),
.B(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_78),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_53),
.A2(n_75),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_53),
.B(n_151),
.Y(n_225)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_55),
.B(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_76),
.B(n_97),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_68),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_66),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_61),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_82),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_61),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_61),
.A2(n_82),
.B1(n_189),
.B2(n_242),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_61),
.A2(n_68),
.B(n_113),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_65),
.A2(n_164),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_65),
.A2(n_81),
.B(n_114),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g315 ( 
.A1(n_71),
.A2(n_72),
.B(n_79),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_74),
.A2(n_76),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_74),
.A2(n_76),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_74),
.A2(n_76),
.B1(n_95),
.B2(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_83),
.B(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_98),
.B(n_99),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_84),
.A2(n_85),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_86),
.A2(n_93),
.B1(n_98),
.B2(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_86),
.A2(n_98),
.B1(n_99),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_92),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_87),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_87),
.A2(n_220),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_87),
.A2(n_92),
.B(n_136),
.Y(n_245)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_88),
.A2(n_135),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_88),
.B(n_137),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_88),
.A2(n_183),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_90),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_92),
.Y(n_209)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_93),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_99),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_103),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_100),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_102),
.B(n_104),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_116),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_326),
.B(n_331),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_311),
.B(n_325),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_292),
.B(n_310),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_191),
.B(n_274),
.C(n_291),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_175),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_130),
.B(n_175),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_156),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_142),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_132),
.B(n_142),
.C(n_156),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_133),
.B(n_140),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_138),
.Y(n_228)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_151),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_141),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.C(n_149),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_177),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_165),
.B2(n_174),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_159),
.B(n_162),
.C(n_174),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_167),
.B1(n_172),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_182),
.B(n_184),
.Y(n_181)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_178),
.B(n_180),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_187),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_184),
.B(n_207),
.Y(n_280)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_187),
.B(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_273),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_268),
.B(n_272),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_253),
.B(n_267),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_236),
.B(n_252),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_216),
.B(n_235),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_204),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_200),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_211),
.C(n_214),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_234),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_222),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_229),
.B(n_233),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_251),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_247),
.C(n_248),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_244),
.B2(n_245),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_255),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_263),
.C(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_271),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_290),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_284),
.C(n_290),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_283),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_283),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_287),
.C(n_289),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_293),
.B(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_309),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_298),
.B1(n_307),
.B2(n_308),
.Y(n_295)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_308),
.C(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_304),
.C(n_306),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_312),
.B(n_313),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_315),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_320),
.C(n_324),
.Y(n_327)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_322),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);


endmodule