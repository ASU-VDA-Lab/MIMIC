module fake_jpeg_1760_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_51),
.Y(n_82)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_22),
.A2(n_39),
.B1(n_37),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_106)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_22),
.B(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_52),
.B(n_63),
.Y(n_105)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_68),
.Y(n_87)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_16),
.B(n_1),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_19),
.B(n_3),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_79),
.Y(n_95)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_41),
.Y(n_77)
);

NOR2xp67_ASAP7_75t_R g119 ( 
.A(n_77),
.B(n_14),
.Y(n_119)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_38),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_88),
.B1(n_90),
.B2(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_40),
.C(n_36),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_120),
.C(n_98),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_38),
.B1(n_33),
.B2(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_106),
.B1(n_114),
.B2(n_45),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_118),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_79),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_14),
.B(n_9),
.C(n_13),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_121),
.B(n_104),
.C(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_50),
.B(n_13),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_107),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_59),
.C(n_61),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_64),
.A3(n_67),
.B1(n_48),
.B2(n_57),
.C1(n_42),
.C2(n_44),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_129),
.C(n_132),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_48),
.B1(n_118),
.B2(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_123),
.A2(n_125),
.B1(n_127),
.B2(n_145),
.Y(n_182)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_105),
.B1(n_83),
.B2(n_92),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_120),
.B1(n_91),
.B2(n_82),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_114),
.Y(n_129)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_130),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_87),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_107),
.B1(n_81),
.B2(n_110),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_158),
.B1(n_154),
.B2(n_149),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_96),
.B1(n_99),
.B2(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_100),
.A2(n_110),
.B1(n_112),
.B2(n_84),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_82),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_97),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_134),
.B(n_131),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_174),
.B(n_166),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_184),
.C(n_168),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_145),
.B1(n_137),
.B2(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_125),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_186),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_128),
.B(n_138),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_129),
.B(n_132),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_136),
.B(n_130),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_141),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_190),
.B(n_195),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_150),
.B1(n_140),
.B2(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_126),
.C(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_162),
.C(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_174),
.B1(n_160),
.B2(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_182),
.B1(n_176),
.B2(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_201),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_177),
.B(n_171),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_205),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_161),
.B1(n_179),
.B2(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_178),
.B1(n_180),
.B2(n_170),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_168),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_203),
.B1(n_193),
.B2(n_206),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_162),
.B(n_178),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_220),
.B(n_207),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_188),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_194),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_190),
.C(n_204),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_195),
.C(n_200),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_222),
.CI(n_197),
.CON(n_229),
.SN(n_229)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_224),
.C(n_225),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_215),
.C(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_230),
.C(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_220),
.B(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_199),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_217),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_231),
.B(n_211),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_210),
.B(n_226),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_232),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_225),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_210),
.B1(n_208),
.B2(n_229),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_224),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_243),
.C(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_247),
.A3(n_229),
.B1(n_214),
.B2(n_213),
.C1(n_223),
.C2(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_255),
.C(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_239),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_259),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_260),
.A2(n_256),
.B(n_214),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_257),
.C(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);


endmodule