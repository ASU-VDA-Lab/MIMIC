module fake_jpeg_6216_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_15),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_60),
.Y(n_77)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AND2x4_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_20),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_26),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_17),
.B(n_20),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_26),
.C(n_23),
.Y(n_79)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_91)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_27),
.B1(n_16),
.B2(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_86),
.B1(n_89),
.B2(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_27),
.B1(n_16),
.B2(n_31),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_47),
.B1(n_27),
.B2(n_16),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_97),
.B1(n_108),
.B2(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_48),
.B(n_69),
.C(n_39),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_113),
.B1(n_71),
.B2(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_72),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_66),
.B1(n_68),
.B2(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_68),
.B1(n_39),
.B2(n_38),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_46),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_77),
.B1(n_86),
.B2(n_21),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_17),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_17),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_80),
.B(n_79),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_29),
.B(n_74),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_114),
.C(n_100),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_126),
.C(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_132),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_77),
.C(n_93),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_94),
.B1(n_96),
.B2(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_130),
.B1(n_95),
.B2(n_97),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_138),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_143),
.C(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_140),
.B1(n_92),
.B2(n_88),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_44),
.B1(n_92),
.B2(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_74),
.C(n_72),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_28),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_105),
.B1(n_103),
.B2(n_106),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_157),
.B1(n_132),
.B2(n_28),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_169),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_148),
.B(n_9),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_99),
.B(n_31),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_123),
.B(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_153),
.B(n_155),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_154),
.A2(n_161),
.B(n_19),
.Y(n_194)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_158),
.B1(n_131),
.B2(n_143),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_108),
.B1(n_44),
.B2(n_111),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_160),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_25),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_17),
.B(n_18),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_25),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_164),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_104),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_104),
.C(n_38),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_168),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_51),
.B1(n_49),
.B2(n_30),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_141),
.B1(n_130),
.B2(n_145),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_119),
.C(n_33),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_33),
.A3(n_19),
.B1(n_28),
.B2(n_4),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_176),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_175),
.B(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_196),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_182),
.B(n_184),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_132),
.B1(n_126),
.B2(n_33),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_153),
.B1(n_168),
.B2(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_33),
.B1(n_19),
.B2(n_3),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_8),
.C(n_14),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_178),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_220),
.B1(n_3),
.B2(n_4),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_146),
.B1(n_171),
.B2(n_149),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_210),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_175),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_159),
.C(n_162),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_174),
.C(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_226),
.C(n_238),
.Y(n_248)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_234),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_183),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_229),
.B(n_230),
.Y(n_256)
);

FAx1_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_194),
.CI(n_195),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_198),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_181),
.B(n_183),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_164),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_206),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_172),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_249),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_238),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_228),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_197),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_200),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_235),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_206),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_224),
.C(n_222),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_254),
.C(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_216),
.C(n_219),
.Y(n_254)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_229),
.B1(n_233),
.B2(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_232),
.C(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_202),
.B(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_5),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_214),
.B(n_239),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_204),
.B(n_4),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_269),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_241),
.B(n_261),
.Y(n_270)
);

O2A1O1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_267),
.B(n_266),
.C(n_258),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_255),
.B(n_244),
.C(n_8),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_260),
.C(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_7),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_278),
.B(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_285),
.B(n_286),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_278),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_276),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_10),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_296),
.B(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_280),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_284),
.B(n_282),
.Y(n_298)
);

NAND2x1_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_292),
.B(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_302),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_291),
.B(n_14),
.C(n_15),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_13),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_15),
.Y(n_307)
);


endmodule