module fake_ariane_758_n_1220 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1220);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1220;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1209;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_1214;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_183;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_1029;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_1167;
wire n_690;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_940;
wire n_756;
wire n_466;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_1131;
wire n_765;
wire n_1187;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_1217;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_207;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_731;
wire n_779;
wire n_336;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_315;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_553;
wire n_446;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_557;
wire n_405;
wire n_1201;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_600;
wire n_433;
wire n_481;
wire n_721;
wire n_840;
wire n_1084;
wire n_1053;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_928;
wire n_839;
wire n_1099;
wire n_218;
wire n_1153;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_478;
wire n_703;
wire n_222;
wire n_1207;
wire n_748;
wire n_1212;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_1074;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_206;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_977;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_1216;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_1218;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_1213;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_181;
wire n_1142;
wire n_658;
wire n_616;
wire n_705;
wire n_630;
wire n_617;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_209;
wire n_743;
wire n_1194;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_1210;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_673;
wire n_452;
wire n_1114;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_571;
wire n_680;
wire n_414;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_609;
wire n_1164;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_872;
wire n_407;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_664;
wire n_629;
wire n_215;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_216;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_213;
wire n_895;
wire n_862;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_204;
wire n_996;
wire n_521;
wire n_1211;
wire n_963;
wire n_873;
wire n_1139;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_289;
wire n_548;
wire n_815;
wire n_542;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1215;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_211;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_119),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_11),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_25),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_89),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_16),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_8),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_125),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_101),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_30),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_152),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_122),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_10),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_4),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_92),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_83),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_72),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_91),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_6),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_29),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_161),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_16),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_114),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_124),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_82),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_44),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_11),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_81),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_178),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_188),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_197),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_198),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_202),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_203),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_225),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_189),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_191),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_192),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_193),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_196),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_199),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_200),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_201),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_254),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_256),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_238),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_236),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_236),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_245),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_264),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_246),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_247),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_237),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_250),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_249),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_251),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_252),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_252),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_235),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_265),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_266),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_291),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_277),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_297),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_294),
.Y(n_338)
);

INVx4_ASAP7_75t_R g339 ( 
.A(n_292),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_294),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_301),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_295),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_303),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_303),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_301),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_267),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_267),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_278),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_318),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_332),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_322),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_325),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_340),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_279),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_343),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_328),
.Y(n_377)
);

NAND2xp33_ASAP7_75t_R g378 ( 
.A(n_343),
.B(n_279),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_356),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_356),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_346),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_346),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_357),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_354),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_354),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_337),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_338),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_338),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_283),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_280),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_393),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_381),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

BUFx8_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_342),
.B1(n_352),
.B2(n_344),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_285),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_280),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_374),
.A2(n_352),
.B1(n_286),
.B2(n_287),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_290),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_349),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_396),
.A2(n_355),
.B1(n_286),
.B2(n_287),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_396),
.A2(n_293),
.B1(n_304),
.B2(n_283),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_350),
.Y(n_425)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_281),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_293),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_378),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_395),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_379),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_368),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_348),
.B(n_347),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_387),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_304),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_390),
.B(n_351),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_394),
.B(n_353),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_358),
.A2(n_305),
.B1(n_313),
.B2(n_314),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_288),
.Y(n_450)
);

AOI22x1_ASAP7_75t_SL g451 ( 
.A1(n_387),
.A2(n_337),
.B1(n_313),
.B2(n_314),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_360),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_289),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_361),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_358),
.B(n_305),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_360),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_358),
.B(n_290),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_366),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_358),
.B(n_290),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_358),
.A2(n_296),
.B1(n_300),
.B2(n_290),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_360),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_358),
.B(n_310),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_434),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_401),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_430),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_430),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_467),
.B(n_290),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_408),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_408),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_326),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_411),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_411),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_327),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_408),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_R g490 ( 
.A(n_434),
.B(n_327),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_440),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g492 ( 
.A(n_459),
.B(n_208),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_440),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_400),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_440),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_413),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_416),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

OA21x2_ASAP7_75t_L g499 ( 
.A1(n_461),
.A2(n_345),
.B(n_186),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_416),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_451),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_413),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_467),
.B(n_208),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_451),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_425),
.B(n_339),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_462),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_462),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_454),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_454),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_458),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_456),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_425),
.B(n_179),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_457),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_490),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_507),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_475),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_475),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_469),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_511),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_511),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_519),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_469),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_496),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_504),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_510),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_508),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_470),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_478),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_470),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_471),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_471),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_472),
.B(n_449),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_486),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_500),
.B(n_438),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_478),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_489),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_468),
.B(n_421),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_489),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_494),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_484),
.B(n_418),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_493),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_495),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_491),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_491),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_514),
.B(n_424),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_402),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_545),
.A2(n_492),
.B1(n_505),
.B2(n_480),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_536),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_538),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_528),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_555),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_524),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_528),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_480),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_538),
.B(n_442),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_534),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_546),
.Y(n_573)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_551),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_533),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_546),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_526),
.Y(n_577)
);

AOI22x1_ASAP7_75t_L g578 ( 
.A1(n_522),
.A2(n_427),
.B1(n_424),
.B2(n_421),
.Y(n_578)
);

BUFx6f_ASAP7_75t_SL g579 ( 
.A(n_546),
.Y(n_579)
);

HAxp5_ASAP7_75t_SL g580 ( 
.A(n_522),
.B(n_437),
.CON(n_580),
.SN(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_542),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_559),
.B(n_465),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_535),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_531),
.B(n_516),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_532),
.B(n_494),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_547),
.A2(n_480),
.B1(n_438),
.B2(n_439),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_553),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_542),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_529),
.B(n_463),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_537),
.A2(n_439),
.B1(n_506),
.B2(n_502),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_539),
.B(n_442),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_543),
.B(n_485),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_544),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_525),
.B(n_497),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_497),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_527),
.B(n_423),
.C(n_417),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_527),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_540),
.B(n_422),
.C(n_446),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_556),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_540),
.B(n_485),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_512),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_552),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_549),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_558),
.B(n_485),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_512),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_558),
.B(n_426),
.C(n_420),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_550),
.B(n_443),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_554),
.B(n_443),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_554),
.B(n_513),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_546),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_554),
.A2(n_439),
.B1(n_437),
.B2(n_518),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_528),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_559),
.B(n_485),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_521),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_538),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_538),
.B(n_513),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_521),
.B(n_439),
.Y(n_623)
);

OAI22xp33_ASAP7_75t_L g624 ( 
.A1(n_554),
.A2(n_439),
.B1(n_506),
.B2(n_502),
.Y(n_624)
);

INVx8_ASAP7_75t_L g625 ( 
.A(n_534),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_534),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_528),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_546),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_528),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_546),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_554),
.A2(n_427),
.B1(n_444),
.B2(n_508),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_521),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_528),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_559),
.B(n_485),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_538),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_528),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_528),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_521),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_521),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_528),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

BUFx4f_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_444),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_622),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_562),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_625),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_625),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_561),
.A2(n_518),
.B1(n_448),
.B2(n_436),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_564),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_606),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_597),
.B(n_473),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_567),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_563),
.B(n_431),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_580),
.B(n_455),
.C(n_450),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_568),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_520),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_602),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_574),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_560),
.A2(n_455),
.B1(n_450),
.B2(n_431),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_560),
.B(n_520),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_613),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_602),
.B(n_445),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_605),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_619),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_578),
.B(n_455),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_625),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_594),
.B(n_429),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_597),
.B(n_473),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_594),
.B(n_429),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_596),
.B(n_428),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_596),
.B(n_447),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_572),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_621),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_632),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_606),
.Y(n_679)
);

BUFx6f_ASAP7_75t_SL g680 ( 
.A(n_606),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_622),
.B(n_487),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_570),
.B(n_518),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_622),
.B(n_487),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_640),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_621),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_600),
.B(n_445),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_610),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_593),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_622),
.Y(n_690)
);

INVx6_ASAP7_75t_L g691 ( 
.A(n_572),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_631),
.A2(n_436),
.B1(n_448),
.B2(n_409),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_641),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_565),
.B(n_473),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_580),
.A2(n_433),
.B1(n_410),
.B2(n_415),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_624),
.B(n_433),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_643),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_621),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_588),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_600),
.B(n_433),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_637),
.B(n_481),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_584),
.B(n_433),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_561),
.A2(n_448),
.B1(n_441),
.B2(n_477),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_612),
.B(n_433),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_586),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_614),
.B(n_476),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_644),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_612),
.B(n_476),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_581),
.B(n_481),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_623),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_566),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_598),
.B(n_432),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_573),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_626),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_644),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_566),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_604),
.B(n_441),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_569),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_572),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_569),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_608),
.B(n_435),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_611),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_575),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_581),
.B(n_582),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_575),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_589),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_591),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_571),
.B(n_479),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_615),
.B(n_487),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_646),
.B(n_581),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_663),
.B(n_603),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_699),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_660),
.B(n_590),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_705),
.B(n_603),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_647),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_709),
.B(n_607),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_708),
.B(n_607),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_651),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_713),
.B(n_571),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_666),
.B(n_590),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_657),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_648),
.B(n_609),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_661),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_646),
.B(n_581),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_689),
.B(n_587),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_724),
.B(n_595),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_704),
.B(n_595),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_646),
.B(n_582),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_658),
.B(n_599),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_664),
.B(n_668),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_678),
.B(n_616),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_685),
.B(n_616),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_648),
.B(n_582),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_658),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_693),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_697),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_667),
.B(n_583),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_711),
.B(n_587),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_655),
.B(n_618),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_723),
.B(n_718),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_730),
.B(n_706),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_688),
.B(n_618),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_684),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_690),
.B(n_582),
.Y(n_766)
);

AO221x1_ASAP7_75t_L g767 ( 
.A1(n_695),
.A2(n_592),
.B1(n_630),
.B2(n_615),
.C(n_636),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_684),
.B(n_635),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_700),
.B(n_635),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_715),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_694),
.B(n_628),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_717),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_SL g773 ( 
.A(n_652),
.B(n_579),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_701),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_726),
.B(n_589),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_691),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_701),
.B(n_628),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_658),
.B(n_576),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_712),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_671),
.B(n_673),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_707),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_674),
.B(n_630),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_691),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_720),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_653),
.B(n_636),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_722),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_669),
.B(n_601),
.C(n_692),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_653),
.B(n_583),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_672),
.B(n_435),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_687),
.B(n_579),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_672),
.B(n_617),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_702),
.B(n_617),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_682),
.B(n_576),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_727),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_728),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_725),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_721),
.B(n_679),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_670),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_714),
.B(n_620),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_710),
.B(n_576),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_714),
.B(n_620),
.Y(n_801)
);

INVxp33_ASAP7_75t_L g802 ( 
.A(n_707),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_698),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_698),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_719),
.B(n_627),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_719),
.B(n_627),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_731),
.B(n_629),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_798),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_798),
.B(n_676),
.Y(n_809)
);

OAI221xp5_ASAP7_75t_L g810 ( 
.A1(n_787),
.A2(n_656),
.B1(n_662),
.B2(n_696),
.C(n_231),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_732),
.B(n_746),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_762),
.B(n_715),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_740),
.Y(n_813)
);

NAND3x1_ASAP7_75t_L g814 ( 
.A(n_790),
.B(n_645),
.C(n_675),
.Y(n_814)
);

NAND3x1_ASAP7_75t_L g815 ( 
.A(n_790),
.B(n_649),
.C(n_680),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_744),
.B(n_729),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_745),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_745),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_780),
.B(n_707),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_752),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_734),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_787),
.A2(n_703),
.B1(n_650),
.B2(n_658),
.Y(n_822)
);

OAI221xp5_ASAP7_75t_L g823 ( 
.A1(n_751),
.A2(n_759),
.B1(n_217),
.B2(n_735),
.C(n_742),
.Y(n_823)
);

AO22x2_ASAP7_75t_L g824 ( 
.A1(n_737),
.A2(n_633),
.B1(n_634),
.B2(n_629),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_757),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_743),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_763),
.B(n_758),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_779),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_796),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_781),
.B(n_716),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_781),
.B(n_716),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_772),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_770),
.B(n_665),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_784),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_736),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_781),
.Y(n_836)
);

BUFx6f_ASAP7_75t_SL g837 ( 
.A(n_781),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_738),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_733),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_786),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_765),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_756),
.B(n_677),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_756),
.B(n_681),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_775),
.B(n_681),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_739),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_794),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_778),
.B(n_726),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_759),
.B(n_731),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_795),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_774),
.B(n_765),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_761),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_764),
.B(n_731),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_775),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_735),
.A2(n_686),
.B1(n_677),
.B2(n_654),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_791),
.Y(n_855)
);

BUFx6f_ASAP7_75t_SL g856 ( 
.A(n_776),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_775),
.B(n_681),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_747),
.A2(n_441),
.B1(n_716),
.B2(n_405),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_742),
.A2(n_686),
.B1(n_659),
.B2(n_576),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_778),
.B(n_681),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_783),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_792),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_748),
.B(n_710),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_L g864 ( 
.A(n_773),
.B(n_683),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_755),
.B(n_487),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_782),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_804),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_753),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_754),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_807),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_799),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_741),
.B(n_801),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_760),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_805),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_797),
.Y(n_875)
);

OAI221xp5_ASAP7_75t_L g876 ( 
.A1(n_789),
.A2(n_234),
.B1(n_180),
.B2(n_233),
.C(n_229),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_806),
.B(n_731),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_768),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_797),
.B(n_683),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_749),
.B(n_683),
.Y(n_880)
);

INVx6_ASAP7_75t_L g881 ( 
.A(n_793),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_788),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_771),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_785),
.B(n_0),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_777),
.Y(n_885)
);

INVx6_ASAP7_75t_L g886 ( 
.A(n_802),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_769),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_839),
.B(n_767),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_808),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_823),
.B(n_766),
.C(n_800),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_845),
.B(n_766),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_835),
.B(n_800),
.Y(n_892)
);

AND2x6_ASAP7_75t_SL g893 ( 
.A(n_809),
.B(n_184),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_808),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_823),
.A2(n_209),
.B(n_212),
.C(n_185),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_870),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_810),
.A2(n_683),
.B1(n_746),
.B2(n_732),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_808),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_836),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_811),
.B(n_750),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_836),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_817),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_866),
.B(n_802),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_818),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_824),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_824),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_838),
.B(n_750),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_811),
.B(n_487),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_878),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_844),
.B(n_498),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_871),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_875),
.B(n_0),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_844),
.B(n_498),
.Y(n_913)
);

CKINVDCx6p67_ASAP7_75t_R g914 ( 
.A(n_856),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_853),
.B(n_633),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_821),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_857),
.B(n_498),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_850),
.B(n_634),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_SL g919 ( 
.A(n_861),
.B(n_509),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_874),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_872),
.B(n_638),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_847),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_857),
.B(n_479),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_867),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_829),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_825),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_810),
.B(n_206),
.C(n_182),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_872),
.B(n_642),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_SL g929 ( 
.A(n_856),
.B(n_498),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_886),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_867),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_851),
.B(n_642),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_841),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_876),
.A2(n_419),
.B(n_221),
.C(n_186),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_812),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_833),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_813),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_820),
.B(n_816),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_822),
.A2(n_474),
.B1(n_419),
.B2(n_482),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_883),
.B(n_639),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_886),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_868),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_847),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_853),
.B(n_498),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_900),
.A2(n_864),
.B(n_876),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_900),
.A2(n_848),
.B(n_880),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_908),
.A2(n_848),
.B(n_880),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_905),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_902),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_890),
.A2(n_814),
.B(n_884),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_942),
.B(n_885),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_943),
.B(n_933),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_897),
.A2(n_852),
.B1(n_877),
.B2(n_854),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_888),
.B(n_852),
.C(n_877),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_908),
.A2(n_854),
.B(n_863),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_914),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_912),
.A2(n_895),
.B(n_934),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_924),
.B(n_887),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_929),
.A2(n_913),
.B(n_910),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_910),
.A2(n_917),
.B(n_913),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_917),
.A2(n_859),
.B(n_819),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_891),
.A2(n_859),
.B(n_827),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_L g963 ( 
.A(n_927),
.B(n_834),
.C(n_828),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_892),
.A2(n_827),
.B(n_860),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_893),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_L g966 ( 
.A1(n_938),
.A2(n_869),
.B(n_873),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_922),
.B(n_860),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_905),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_912),
.A2(n_938),
.B(n_934),
.C(n_922),
.Y(n_969)
);

AO32x2_ASAP7_75t_L g970 ( 
.A1(n_924),
.A2(n_862),
.A3(n_855),
.B1(n_882),
.B2(n_826),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_944),
.A2(n_843),
.B(n_879),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_904),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_944),
.A2(n_843),
.B(n_842),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_936),
.B(n_881),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_931),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_907),
.A2(n_842),
.B(n_853),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_931),
.A2(n_815),
.B(n_830),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_894),
.B(n_881),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_919),
.B(n_903),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_916),
.B(n_847),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_935),
.B(n_836),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_889),
.B(n_215),
.C(n_213),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_926),
.A2(n_831),
.B(n_858),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_921),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_906),
.A2(n_221),
.B(n_226),
.C(n_224),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_928),
.A2(n_840),
.B(n_832),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_930),
.B(n_847),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_896),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_899),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_889),
.A2(n_849),
.B(n_846),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_481),
.C(n_452),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_930),
.B(n_941),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_941),
.B(n_865),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_940),
.A2(n_183),
.B(n_195),
.C(n_181),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_932),
.A2(n_837),
.B(n_499),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_898),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_937),
.A2(n_499),
.B(n_837),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_899),
.A2(n_464),
.B1(n_466),
.B2(n_460),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_899),
.B(n_639),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_899),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_909),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_918),
.B(n_499),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_901),
.A2(n_499),
.B(n_483),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_911),
.B(n_1),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_901),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_909),
.A2(n_638),
.B(n_483),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_925),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_920),
.A2(n_181),
.B(n_406),
.C(n_460),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_901),
.A2(n_482),
.B(n_466),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_901),
.A2(n_464),
.B(n_488),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_979),
.B(n_915),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_987),
.B(n_915),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_SL g1013 ( 
.A(n_952),
.B(n_923),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_963),
.B(n_923),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_956),
.B(n_1005),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_987),
.B(n_939),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_SL g1017 ( 
.A(n_996),
.B(n_923),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_967),
.B(n_923),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_967),
.B(n_923),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_977),
.B(n_181),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_962),
.B(n_410),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_989),
.B(n_975),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_955),
.B(n_410),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_989),
.B(n_410),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_989),
.B(n_410),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_959),
.B(n_961),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_978),
.B(n_1),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_964),
.B(n_414),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_960),
.B(n_414),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_951),
.B(n_2),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_974),
.B(n_992),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_946),
.B(n_414),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_1018),
.B(n_945),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1026),
.B(n_1030),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_950),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1027),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_1020),
.A2(n_957),
.B(n_994),
.C(n_969),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1014),
.A2(n_954),
.B1(n_980),
.B2(n_953),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1021),
.B(n_949),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_1018),
.B(n_965),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_SL g1041 ( 
.A(n_1019),
.B(n_981),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_SL g1042 ( 
.A1(n_1023),
.A2(n_1011),
.B(n_1016),
.C(n_993),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_SL g1043 ( 
.A1(n_1022),
.A2(n_1000),
.B(n_982),
.C(n_983),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_1019),
.B(n_1000),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1032),
.A2(n_971),
.B1(n_947),
.B2(n_973),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1012),
.B(n_972),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1028),
.A2(n_976),
.B1(n_958),
.B2(n_985),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_1024),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1029),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_1015),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1025),
.B(n_984),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1013),
.B(n_966),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_1017),
.B(n_998),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1026),
.A2(n_1004),
.B(n_1008),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_1015),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_1027),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1026),
.A2(n_991),
.B1(n_999),
.B2(n_995),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1031),
.B(n_990),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_1044),
.A2(n_968),
.B(n_948),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_990),
.B1(n_1009),
.B2(n_1007),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_1035),
.A2(n_1001),
.A3(n_988),
.B(n_1010),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_1036),
.A2(n_986),
.B(n_997),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_1056),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_L g1064 ( 
.A(n_1043),
.B(n_1002),
.C(n_1003),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_1056),
.B(n_1006),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_1063),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_1063),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_1067),
.B(n_1034),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_1066),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1068),
.A2(n_1059),
.B(n_1033),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1069),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1071),
.A2(n_1050),
.B1(n_1052),
.B2(n_1056),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1071),
.B(n_1054),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1073),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1072),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_1067),
.Y(n_1076)
);

BUFx4f_ASAP7_75t_SL g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AOI222xp33_ASAP7_75t_L g1078 ( 
.A1(n_1074),
.A2(n_1070),
.B1(n_1037),
.B2(n_1066),
.C1(n_1067),
.C2(n_1065),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1076),
.B(n_1055),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1078),
.B(n_1066),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_1077),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_R g1082 ( 
.A(n_1081),
.B(n_1040),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_1046),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1083),
.B(n_1079),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1082),
.B(n_1080),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_1041),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1086),
.A2(n_1064),
.B1(n_1062),
.B2(n_1060),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1087),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1089),
.B(n_1061),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1088),
.A2(n_1057),
.B1(n_1049),
.B2(n_1047),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1090),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1091),
.A2(n_1042),
.B(n_1038),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_206),
.C(n_182),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_1093),
.B(n_227),
.C(n_207),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1092),
.A2(n_1053),
.B1(n_1048),
.B2(n_1045),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_3),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_1051),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1094),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1098),
.B(n_1048),
.Y(n_1100)
);

NAND2x1_ASAP7_75t_L g1101 ( 
.A(n_1097),
.B(n_1048),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_SL g1102 ( 
.A(n_1100),
.B(n_1099),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1101),
.B(n_1039),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1102),
.B(n_3),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1103),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1104),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_970),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1106),
.Y(n_1108)
);

NAND4xp25_ASAP7_75t_L g1109 ( 
.A(n_1107),
.B(n_5),
.C(n_7),
.D(n_8),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_L g1110 ( 
.A(n_1108),
.B(n_5),
.C(n_7),
.D(n_9),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1109),
.B(n_9),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1111),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_227),
.B(n_207),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1111),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1114),
.B(n_10),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1112),
.B(n_12),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1113),
.B(n_12),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_1116),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1115),
.B(n_13),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_1118),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1119),
.B(n_1117),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_232),
.B(n_211),
.Y(n_1122)
);

OAI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_232),
.B(n_216),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1123),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1122),
.B(n_14),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1124),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1125),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1126),
.B(n_219),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_1127),
.B(n_218),
.C(n_204),
.Y(n_1129)
);

AO22x2_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_1130)
);

NAND4xp25_ASAP7_75t_L g1131 ( 
.A(n_1128),
.B(n_15),
.C(n_17),
.D(n_18),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_L g1132 ( 
.A(n_1129),
.B(n_219),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_R g1133 ( 
.A(n_1132),
.B(n_18),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1130),
.Y(n_1134)
);

AOI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_1131),
.A2(n_222),
.B1(n_223),
.B2(n_219),
.C(n_230),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1134),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_1135),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1136),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1137),
.A2(n_1133),
.B(n_230),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1138),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1139),
.A2(n_230),
.B1(n_405),
.B2(n_407),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1140),
.B(n_19),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1141),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1143),
.Y(n_1144)
);

NAND4xp75_ASAP7_75t_L g1145 ( 
.A(n_1142),
.B(n_19),
.C(n_20),
.D(n_21),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1144),
.Y(n_1146)
);

AND4x2_ASAP7_75t_L g1147 ( 
.A(n_1145),
.B(n_20),
.C(n_21),
.D(n_22),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_R g1148 ( 
.A(n_1146),
.B(n_22),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1147),
.B(n_23),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1146),
.B(n_230),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1149),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1148),
.B(n_23),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1150),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1153)
);

AO22x1_ASAP7_75t_L g1154 ( 
.A1(n_1151),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1152),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1155),
.A2(n_1153),
.B1(n_28),
.B2(n_29),
.Y(n_1156)
);

AO21x2_ASAP7_75t_L g1157 ( 
.A1(n_1154),
.A2(n_27),
.B(n_30),
.Y(n_1157)
);

OR5x1_ASAP7_75t_L g1158 ( 
.A(n_1156),
.B(n_31),
.C(n_32),
.D(n_33),
.E(n_34),
.Y(n_1158)
);

NAND4xp75_ASAP7_75t_L g1159 ( 
.A(n_1157),
.B(n_32),
.C(n_33),
.D(n_34),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_1159),
.B(n_35),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1158),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1160),
.B(n_35),
.C(n_37),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1161),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1163),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1162),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1164),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_1166)
);

XNOR2xp5_ASAP7_75t_L g1167 ( 
.A(n_1165),
.B(n_43),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1164),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1167),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1166),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1168),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1171)
);

AOI31xp33_ASAP7_75t_L g1172 ( 
.A1(n_1169),
.A2(n_54),
.A3(n_55),
.B(n_56),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1171),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1173),
.A2(n_1170),
.B1(n_61),
.B2(n_63),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1172),
.Y(n_1175)
);

XNOR2xp5_ASAP7_75t_L g1176 ( 
.A(n_1173),
.B(n_60),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1175),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1176),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1174),
.Y(n_1179)
);

OAI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1177),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_1180)
);

OAI222xp33_ASAP7_75t_L g1181 ( 
.A1(n_1179),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.C1(n_74),
.C2(n_75),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1178),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1182),
.A2(n_1181),
.B(n_1180),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_1182),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1182),
.B(n_76),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1182),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1186)
);

AOI221xp5_ASAP7_75t_L g1187 ( 
.A1(n_1182),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.C(n_86),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1182),
.A2(n_87),
.B(n_88),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1182),
.B(n_90),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1182),
.B(n_93),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1182),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_1191)
);

INVxp33_ASAP7_75t_L g1192 ( 
.A(n_1182),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1182),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1182),
.A2(n_104),
.B(n_105),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_1182),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.C(n_111),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1192),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_1196)
);

XNOR2xp5_ASAP7_75t_L g1197 ( 
.A(n_1184),
.B(n_116),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1183),
.A2(n_117),
.B(n_118),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1194),
.A2(n_1187),
.B1(n_1195),
.B2(n_1191),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1186),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1188),
.A2(n_1193),
.B(n_1190),
.Y(n_1201)
);

AO21x2_ASAP7_75t_L g1202 ( 
.A1(n_1185),
.A2(n_120),
.B(n_121),
.Y(n_1202)
);

OAI221xp5_ASAP7_75t_L g1203 ( 
.A1(n_1189),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.C(n_129),
.Y(n_1203)
);

XOR2xp5_ASAP7_75t_L g1204 ( 
.A(n_1192),
.B(n_130),
.Y(n_1204)
);

XOR2x2_ASAP7_75t_L g1205 ( 
.A(n_1201),
.B(n_134),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1199),
.B(n_135),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1202),
.B(n_137),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1200),
.A2(n_138),
.B(n_139),
.Y(n_1208)
);

XNOR2xp5_ASAP7_75t_L g1209 ( 
.A(n_1198),
.B(n_140),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1197),
.Y(n_1210)
);

AOI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1204),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1210),
.A2(n_1203),
.B1(n_1196),
.B2(n_147),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1206),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_1213)
);

AOI322xp5_ASAP7_75t_L g1214 ( 
.A1(n_1212),
.A2(n_1205),
.A3(n_1207),
.B1(n_1208),
.B2(n_1211),
.C1(n_1209),
.C2(n_158),
.Y(n_1214)
);

OA22x2_ASAP7_75t_L g1215 ( 
.A1(n_1214),
.A2(n_1213),
.B1(n_151),
.B2(n_153),
.Y(n_1215)
);

OAI221xp5_ASAP7_75t_R g1216 ( 
.A1(n_1215),
.A2(n_150),
.B1(n_155),
.B2(n_157),
.C(n_159),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1216),
.A2(n_160),
.B(n_163),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1217),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_1218)
);

AOI211xp5_ASAP7_75t_L g1219 ( 
.A1(n_1218),
.A2(n_168),
.B(n_169),
.C(n_172),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_173),
.B(n_175),
.C(n_176),
.Y(n_1220)
);


endmodule