module fake_jpeg_2365_n_378 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_4),
.B(n_1),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_10),
.B(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_46),
.Y(n_123)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_21),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_17),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_0),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_24),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_24),
.A2(n_2),
.B(n_3),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_40),
.C(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_79),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_2),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_3),
.Y(n_122)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_86),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_64),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_36),
.B1(n_34),
.B2(n_37),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_19),
.B1(n_105),
.B2(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_36),
.B1(n_34),
.B2(n_28),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_43),
.B1(n_50),
.B2(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_19),
.B1(n_36),
.B2(n_31),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_41),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_109),
.B(n_114),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_45),
.A2(n_17),
.B1(n_31),
.B2(n_26),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_56),
.B1(n_77),
.B2(n_60),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_47),
.B(n_35),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_115),
.B(n_127),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_19),
.B1(n_31),
.B2(n_33),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_125),
.B1(n_71),
.B2(n_73),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_SL g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_25),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_43),
.A2(n_15),
.B1(n_30),
.B2(n_25),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_15),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_131),
.A2(n_161),
.B1(n_166),
.B2(n_172),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_145),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_175),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_54),
.B1(n_30),
.B2(n_33),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_134),
.A2(n_146),
.B1(n_110),
.B2(n_144),
.Y(n_207)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_55),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_138),
.B(n_150),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_107),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_94),
.B1(n_125),
.B2(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_140),
.A2(n_155),
.B1(n_110),
.B2(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_141),
.B(n_164),
.Y(n_190)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_49),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_102),
.A2(n_112),
.B(n_95),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_148),
.A2(n_151),
.B(n_138),
.Y(n_212)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

OR2x4_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_111),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_26),
.B(n_65),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_59),
.B1(n_66),
.B2(n_87),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_162),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_29),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_165),
.C(n_177),
.Y(n_182)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_4),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_168),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_84),
.A2(n_26),
.B1(n_29),
.B2(n_6),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_83),
.B(n_4),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_29),
.C(n_5),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_84),
.A2(n_98),
.B1(n_87),
.B2(n_103),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_4),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_6),
.C(n_7),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_171),
.Y(n_194)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_81),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_106),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_96),
.B(n_7),
.C(n_8),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_85),
.B(n_9),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_10),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_180),
.B(n_219),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_85),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_185),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_148),
.A2(n_130),
.B1(n_118),
.B2(n_106),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_195),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_191),
.A2(n_220),
.B(n_215),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_10),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_204),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_118),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_107),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_142),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_208),
.B(n_212),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_110),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_209),
.B(n_211),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_140),
.A2(n_135),
.B1(n_139),
.B2(n_147),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_210),
.A2(n_211),
.B1(n_216),
.B2(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_150),
.B1(n_151),
.B2(n_133),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_153),
.A2(n_156),
.B1(n_163),
.B2(n_174),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_137),
.B1(n_162),
.B2(n_145),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_132),
.B(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_187),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_133),
.A2(n_165),
.B1(n_149),
.B2(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_152),
.B(n_143),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_241),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_225),
.A2(n_217),
.B1(n_203),
.B2(n_193),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_227),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_244),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_173),
.B1(n_159),
.B2(n_167),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_246),
.B1(n_203),
.B2(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_242),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_209),
.B(n_188),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_182),
.B(n_136),
.C(n_137),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_238),
.C(n_249),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_137),
.C(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_245),
.B(n_247),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_208),
.A2(n_212),
.B1(n_220),
.B2(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_186),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_199),
.B(n_184),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_205),
.B(n_209),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_188),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_189),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_251),
.A2(n_252),
.B1(n_209),
.B2(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_188),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_253),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_198),
.C(n_190),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_255),
.A2(n_256),
.B(n_260),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_213),
.B1(n_185),
.B2(n_205),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_263),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_194),
.B(n_213),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_269),
.B1(n_273),
.B2(n_283),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_194),
.B(n_191),
.Y(n_267)
);

AOI221xp5_ASAP7_75t_L g302 ( 
.A1(n_267),
.A2(n_280),
.B1(n_255),
.B2(n_282),
.C(n_257),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_226),
.A2(n_218),
.B(n_193),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_274),
.C(n_277),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_246),
.A2(n_198),
.B1(n_190),
.B2(n_201),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_201),
.C(n_238),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_228),
.A2(n_201),
.B1(n_241),
.B2(n_221),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_278),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_254),
.C(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_227),
.B1(n_224),
.B2(n_236),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_236),
.A2(n_242),
.B(n_223),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_247),
.B1(n_244),
.B2(n_222),
.Y(n_283)
);

AO22x1_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_234),
.B1(n_243),
.B2(n_251),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_262),
.B(n_231),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_259),
.A2(n_231),
.B1(n_230),
.B2(n_235),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_291),
.A2(n_295),
.B1(n_297),
.B2(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_229),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_292),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_274),
.C(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_296),
.C(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_232),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_232),
.C(n_239),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_270),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_299),
.A2(n_305),
.B(n_304),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_240),
.C(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_303),
.A2(n_275),
.B1(n_261),
.B2(n_284),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_281),
.Y(n_304)
);

XOR2x2_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_308),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_266),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_257),
.B(n_261),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_263),
.A3(n_260),
.B1(n_267),
.B2(n_275),
.C(n_264),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_268),
.C(n_258),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

AO22x1_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_284),
.B1(n_276),
.B2(n_280),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_313),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_273),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_314),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_325),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_317),
.C(n_310),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_291),
.A2(n_260),
.B1(n_269),
.B2(n_300),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_286),
.B1(n_290),
.B2(n_297),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_287),
.C(n_296),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_323),
.C(n_311),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_288),
.B(n_300),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_307),
.C(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_298),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_329),
.A2(n_343),
.B1(n_331),
.B2(n_332),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_285),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_333),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_285),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_336),
.C(n_341),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_335),
.A2(n_329),
.B1(n_330),
.B2(n_336),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_303),
.C(n_312),
.Y(n_336)
);

OA21x2_ASAP7_75t_SL g337 ( 
.A1(n_322),
.A2(n_319),
.B(n_327),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_337),
.B(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_340),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_315),
.C(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_333),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_345),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_338),
.B(n_321),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_334),
.B(n_326),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_348),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_328),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_354),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_350),
.A2(n_339),
.B(n_351),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_353),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_341),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_355),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_355),
.B(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_363),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_357),
.A2(n_362),
.B(n_352),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_354),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_352),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_367),
.C(n_368),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_359),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_364),
.C(n_360),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_372),
.A2(n_346),
.B(n_349),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_360),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_373),
.B(n_350),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_374),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_370),
.C(n_371),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_375),
.Y(n_378)
);


endmodule