module fake_jpeg_284_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_29),
.B(n_26),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_72),
.Y(n_79)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_85),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_61),
.B1(n_54),
.B2(n_62),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_59),
.B1(n_66),
.B2(n_57),
.Y(n_92)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_55),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_63),
.C(n_61),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_64),
.B1(n_54),
.B2(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_98),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_83),
.B1(n_78),
.B2(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_96),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_59),
.B1(n_56),
.B2(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_1),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_58),
.C(n_19),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_58),
.C(n_24),
.Y(n_130)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_20),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_4),
.B(n_5),
.C(n_7),
.D(n_8),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_97),
.B(n_58),
.C(n_22),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_112),
.B(n_11),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.C(n_35),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_135),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_28),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_111),
.C(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_118),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_121),
.B(n_120),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_150),
.B(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_157),
.B1(n_134),
.B2(n_125),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_123),
.B1(n_16),
.B2(n_18),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_123),
.B1(n_31),
.B2(n_32),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_15),
.B1(n_36),
.B2(n_37),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_157),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_151),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_153),
.C(n_149),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_158),
.C(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_162),
.B1(n_154),
.B2(n_152),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_162),
.C(n_170),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_169),
.B1(n_166),
.B2(n_44),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_175),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_176),
.B(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_39),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_40),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_45),
.Y(n_186)
);


endmodule