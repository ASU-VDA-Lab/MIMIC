module real_jpeg_30481_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_4;
wire n_12;
wire n_8;
wire n_11;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

INVx4_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_10),
.Y(n_11)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx1_ASAP7_75t_L g3 ( 
.A(n_4),
.Y(n_3)
);

OAI22xp33_ASAP7_75t_SL g4 ( 
.A1(n_5),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_4)
);

INVx1_ASAP7_75t_L g5 ( 
.A(n_6),
.Y(n_5)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_10),
.B(n_11),
.Y(n_7)
);

INVx2_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);


endmodule