module fake_ibex_159_n_899 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_899);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_899;

wire n_151;
wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_280;
wire n_340;
wire n_708;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_136;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_141;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_139;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_137;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_135;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_164;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g135 ( 
.A(n_38),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_36),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_46),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_34),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_27),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_24),
.Y(n_152)
);

INVxp33_ASAP7_75t_SL g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_26),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_13),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_40),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_23),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_101),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_77),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_20),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_50),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_51),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_99),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_122),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_88),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_31),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_62),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_11),
.B(n_95),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_19),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_35),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_86),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_7),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_69),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_59),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_37),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_44),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_133),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_56),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_103),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_68),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_76),
.Y(n_209)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_127),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_12),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_79),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_92),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_89),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_85),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_125),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_48),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_108),
.B(n_128),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_52),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_25),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_29),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_78),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_146),
.B(n_43),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_163),
.B(n_0),
.Y(n_239)
);

BUFx8_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_45),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_161),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_1),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_152),
.B1(n_173),
.B2(n_182),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_2),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_139),
.B(n_4),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_156),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_168),
.B(n_5),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_167),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_170),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_180),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_144),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_144),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_153),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_194),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_216),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_186),
.B(n_49),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_169),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_153),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_180),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_144),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_139),
.B(n_14),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_192),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_192),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_137),
.B(n_151),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_183),
.B(n_15),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_144),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_174),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_183),
.B(n_17),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_135),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_196),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_217),
.B(n_17),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_155),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_155),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_136),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_217),
.B(n_18),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_138),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_140),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_141),
.B(n_18),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_142),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_143),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_145),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_196),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_181),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_147),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_137),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_255),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_148),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_234),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_149),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_213),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_154),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_288),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_257),
.B(n_158),
.Y(n_326)
);

BUFx4f_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_264),
.B(n_151),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

CKINVDCx8_ASAP7_75t_R g330 ( 
.A(n_267),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_266),
.B(n_210),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_266),
.B(n_171),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_235),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_235),
.B(n_159),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_234),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_240),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_252),
.B(n_160),
.Y(n_341)
);

BUFx6f_ASAP7_75t_SL g342 ( 
.A(n_234),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_252),
.B(n_162),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_244),
.B(n_164),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_220),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_266),
.B(n_220),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_223),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_234),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_293),
.B(n_165),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_261),
.B(n_223),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_309),
.B(n_166),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_240),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_262),
.B(n_227),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_309),
.B(n_197),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_254),
.B(n_202),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_241),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_234),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_249),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_254),
.B(n_232),
.C(n_172),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_249),
.Y(n_363)
);

AND2x6_ASAP7_75t_L g364 ( 
.A(n_310),
.B(n_175),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_254),
.B(n_218),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_258),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_258),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_234),
.B(n_291),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_270),
.B(n_179),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_176),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_295),
.B(n_177),
.Y(n_371)
);

INVx4_ASAP7_75t_SL g372 ( 
.A(n_300),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_288),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g374 ( 
.A(n_300),
.B(n_178),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_267),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_259),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_241),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_184),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g380 ( 
.A(n_294),
.B(n_208),
.C(n_187),
.Y(n_380)
);

INVx4_ASAP7_75t_SL g381 ( 
.A(n_302),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_281),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_237),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_250),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_265),
.Y(n_388)
);

BUFx8_ASAP7_75t_SL g389 ( 
.A(n_242),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_303),
.B(n_185),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_303),
.B(n_209),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_305),
.B(n_211),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_273),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_305),
.B(n_205),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_237),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_237),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_265),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_281),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_236),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_282),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_301),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_310),
.B(n_212),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_250),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_237),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_306),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_286),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_306),
.B(n_307),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_268),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_268),
.Y(n_409)
);

OAI22x1_ASAP7_75t_L g410 ( 
.A1(n_285),
.A2(n_229),
.B1(n_221),
.B2(n_222),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_307),
.B(n_201),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_269),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_245),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_287),
.B(n_190),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_290),
.B(n_219),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_236),
.B(n_204),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_269),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_271),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_236),
.B(n_198),
.Y(n_419)
);

NAND2x1p5_ASAP7_75t_L g420 ( 
.A(n_263),
.B(n_191),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_246),
.B(n_271),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_246),
.B(n_228),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_238),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_327),
.A2(n_263),
.B1(n_292),
.B2(n_283),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_313),
.B(n_285),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_389),
.Y(n_427)
);

BUFx12f_ASAP7_75t_L g428 ( 
.A(n_312),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_304),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_321),
.B(n_239),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_316),
.B(n_276),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_246),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_316),
.B(n_338),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_349),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_317),
.A2(n_292),
.B(n_283),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_378),
.B(n_276),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_420),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_329),
.B(n_331),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_378),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_338),
.Y(n_443)
);

AND2x6_ASAP7_75t_SL g444 ( 
.A(n_345),
.B(n_274),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_343),
.A2(n_315),
.B1(n_327),
.B2(n_355),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_343),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_375),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_308),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_L g450 ( 
.A1(n_398),
.A2(n_272),
.B1(n_280),
.B2(n_296),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_339),
.B(n_308),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_352),
.B(n_296),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_323),
.A2(n_326),
.B1(n_315),
.B2(n_341),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_392),
.Y(n_455)
);

NOR3xp33_ASAP7_75t_SL g456 ( 
.A(n_382),
.B(n_277),
.C(n_242),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_R g458 ( 
.A(n_312),
.B(n_274),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_330),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_320),
.A2(n_225),
.B1(n_200),
.B2(n_250),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_341),
.B(n_326),
.Y(n_461)
);

NOR3xp33_ASAP7_75t_SL g462 ( 
.A(n_311),
.B(n_365),
.C(n_358),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_368),
.A2(n_250),
.B(n_260),
.Y(n_464)
);

NOR2x1p5_ASAP7_75t_L g465 ( 
.A(n_314),
.B(n_200),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_343),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_412),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_415),
.B(n_19),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_332),
.B(n_279),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_325),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_320),
.A2(n_279),
.B1(n_260),
.B2(n_238),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_412),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_320),
.A2(n_324),
.B1(n_364),
.B2(n_390),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_360),
.B(n_260),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_314),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_360),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_320),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_323),
.Y(n_486)
);

OR2x2_ASAP7_75t_SL g487 ( 
.A(n_373),
.B(n_21),
.Y(n_487)
);

NOR3xp33_ASAP7_75t_SL g488 ( 
.A(n_380),
.B(n_24),
.C(n_25),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_393),
.B(n_27),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_400),
.A2(n_279),
.B1(n_238),
.B2(n_30),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_336),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_347),
.B(n_28),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_324),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_335),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_342),
.B(n_33),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_324),
.Y(n_498)
);

BUFx4f_ASAP7_75t_L g499 ( 
.A(n_324),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_318),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_348),
.B(n_39),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_379),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_364),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_418),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_322),
.B(n_41),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

OR2x6_ASAP7_75t_SL g507 ( 
.A(n_340),
.B(n_42),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_336),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_346),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_47),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_364),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_340),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_351),
.B(n_53),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_422),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_353),
.B(n_54),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_342),
.B(n_55),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_328),
.B(n_57),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_383),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_448),
.B(n_410),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_431),
.A2(n_317),
.B(n_319),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_333),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_440),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_442),
.B(n_374),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_451),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_430),
.A2(n_374),
.B1(n_390),
.B2(n_370),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_436),
.A2(n_361),
.B(n_367),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_426),
.B(n_371),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_486),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_458),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_439),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_439),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_467),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_482),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_433),
.A2(n_394),
.B(n_391),
.C(n_385),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_442),
.A2(n_362),
.B1(n_411),
.B2(n_419),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_432),
.Y(n_538)
);

OAI21xp33_ASAP7_75t_SL g539 ( 
.A1(n_445),
.A2(n_402),
.B(n_414),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_499),
.B(n_386),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_455),
.B(n_357),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_430),
.B(n_422),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_457),
.A2(n_374),
.B1(n_390),
.B2(n_344),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_441),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_461),
.B(n_416),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_434),
.A2(n_359),
.B(n_377),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_482),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_441),
.A2(n_374),
.B1(n_390),
.B2(n_344),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_464),
.A2(n_511),
.B(n_492),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_458),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_491),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_452),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_467),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_427),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_465),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_508),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_509),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_471),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_461),
.B(n_344),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_470),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_471),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_454),
.A2(n_344),
.B1(n_376),
.B2(n_366),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_482),
.B(n_361),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_444),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_409),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_453),
.B(n_367),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_480),
.B(n_366),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_509),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_450),
.A2(n_363),
.B1(n_408),
.B2(n_397),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_476),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_425),
.B(n_363),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

CKINVDCx8_ASAP7_75t_R g581 ( 
.A(n_513),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_425),
.B(n_485),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_493),
.B(n_403),
.Y(n_583)
);

A2O1A1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_505),
.A2(n_423),
.B(n_404),
.C(n_396),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_493),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_504),
.B(n_403),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_504),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_479),
.A2(n_387),
.B(n_404),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_462),
.B(n_483),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_487),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_452),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_483),
.B(n_498),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_506),
.A2(n_423),
.B1(n_404),
.B2(n_396),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_484),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_519),
.A2(n_423),
.B1(n_396),
.B2(n_395),
.Y(n_598)
);

CKINVDCx11_ASAP7_75t_R g599 ( 
.A(n_507),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_SL g601 ( 
.A1(n_501),
.A2(n_65),
.B(n_66),
.C(n_71),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_472),
.A2(n_395),
.B(n_384),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_512),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_449),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_512),
.A2(n_395),
.B(n_384),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_468),
.B(n_477),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_515),
.B(n_81),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_435),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_462),
.B(n_83),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_435),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_446),
.B(n_469),
.Y(n_611)
);

AO21x2_ASAP7_75t_L g612 ( 
.A1(n_584),
.A2(n_516),
.B(n_514),
.Y(n_612)
);

NAND4xp25_ASAP7_75t_L g613 ( 
.A(n_543),
.B(n_494),
.C(n_450),
.D(n_456),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_581),
.B(n_499),
.Y(n_614)
);

OA21x2_ASAP7_75t_L g615 ( 
.A1(n_584),
.A2(n_536),
.B(n_602),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_572),
.Y(n_616)
);

AO31x2_ASAP7_75t_L g617 ( 
.A1(n_536),
.A2(n_490),
.A3(n_505),
.B(n_518),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_567),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_569),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_569),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_527),
.A2(n_460),
.B(n_474),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_597),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_604),
.A2(n_456),
.B1(n_478),
.B2(n_488),
.C(n_424),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_545),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_589),
.B(n_498),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_553),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_574),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_546),
.B(n_528),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_522),
.A2(n_478),
.B(n_438),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_595),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_559),
.B(n_463),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_605),
.A2(n_496),
.B(n_500),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_588),
.A2(n_475),
.B(n_503),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_606),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_576),
.A2(n_473),
.B1(n_510),
.B2(n_497),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_582),
.A2(n_539),
.B(n_579),
.C(n_520),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_522),
.B(n_510),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_561),
.A2(n_503),
.B1(n_512),
.B2(n_488),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_558),
.B(n_466),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_565),
.B(n_466),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_589),
.B(n_475),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_531),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_532),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_606),
.B(n_517),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_521),
.A2(n_517),
.B(n_497),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_532),
.A2(n_517),
.B(n_497),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_552),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_533),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_554),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_563),
.A2(n_447),
.B(n_443),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_578),
.A2(n_447),
.B(n_443),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_558),
.B(n_337),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_609),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_523),
.B(n_592),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_557),
.Y(n_658)
);

CKINVDCx11_ASAP7_75t_R g659 ( 
.A(n_555),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_577),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_537),
.A2(n_113),
.B(n_115),
.C(n_117),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_564),
.Y(n_662)
);

OA21x2_ASAP7_75t_L g663 ( 
.A1(n_580),
.A2(n_129),
.B(n_587),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_593),
.B(n_596),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_587),
.A2(n_568),
.B(n_598),
.Y(n_665)
);

BUFx2_ASAP7_75t_R g666 ( 
.A(n_530),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_573),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_603),
.Y(n_668)
);

AO31x2_ASAP7_75t_L g669 ( 
.A1(n_585),
.A2(n_524),
.A3(n_610),
.B(n_608),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_542),
.B(n_571),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_598),
.A2(n_594),
.B(n_610),
.Y(n_671)
);

AO21x2_ASAP7_75t_L g672 ( 
.A1(n_601),
.A2(n_550),
.B(n_566),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_571),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_534),
.B(n_570),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_599),
.A2(n_591),
.B1(n_526),
.B2(n_549),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_562),
.B(n_526),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_599),
.A2(n_549),
.B1(n_538),
.B2(n_544),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_583),
.A2(n_586),
.B(n_608),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_534),
.B(n_593),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_544),
.A2(n_607),
.B(n_594),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_611),
.B(n_538),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_540),
.A2(n_525),
.B(n_600),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_556),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_593),
.A2(n_560),
.B1(n_596),
.B2(n_575),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_541),
.A2(n_535),
.B(n_548),
.C(n_590),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_535),
.A2(n_548),
.B1(n_590),
.B2(n_551),
.Y(n_687)
);

CKINVDCx11_ASAP7_75t_R g688 ( 
.A(n_603),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_548),
.B(n_590),
.Y(n_689)
);

AO31x2_ASAP7_75t_L g690 ( 
.A1(n_603),
.A2(n_584),
.A3(n_536),
.B(n_582),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_546),
.B(n_448),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_536),
.A2(n_539),
.B(n_327),
.C(n_582),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_572),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_569),
.Y(n_694)
);

OA21x2_ASAP7_75t_L g695 ( 
.A1(n_584),
.A2(n_536),
.B(n_602),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_531),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_572),
.B(n_442),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_572),
.B(n_442),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_553),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_536),
.A2(n_522),
.B(n_547),
.Y(n_700)
);

AOI21xp33_ASAP7_75t_SL g701 ( 
.A1(n_592),
.A2(n_427),
.B(n_281),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_572),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_561),
.B(n_340),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_527),
.A2(n_436),
.B(n_602),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_527),
.A2(n_436),
.B(n_602),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_561),
.A2(n_267),
.B1(n_285),
.B2(n_281),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_558),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_527),
.A2(n_436),
.B(n_602),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_675),
.A2(n_619),
.B1(n_620),
.B2(n_694),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g710 ( 
.A1(n_691),
.A2(n_699),
.B1(n_614),
.B2(n_635),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_707),
.Y(n_711)
);

CKINVDCx10_ASAP7_75t_R g712 ( 
.A(n_659),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_628),
.B(n_706),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_692),
.A2(n_672),
.B(n_700),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_707),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_633),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_616),
.B(n_693),
.Y(n_717)
);

CKINVDCx11_ASAP7_75t_R g718 ( 
.A(n_659),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_619),
.A2(n_620),
.B1(n_694),
.B2(n_698),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_679),
.B(n_697),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_679),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_692),
.A2(n_672),
.B(n_645),
.Y(n_722)
);

AOI221xp5_ASAP7_75t_L g723 ( 
.A1(n_702),
.A2(n_627),
.B1(n_622),
.B2(n_618),
.C(n_637),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_679),
.A2(n_670),
.B1(n_623),
.B2(n_674),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_688),
.Y(n_725)
);

AOI222xp33_ASAP7_75t_L g726 ( 
.A1(n_630),
.A2(n_677),
.B1(n_624),
.B2(n_673),
.C1(n_703),
.C2(n_648),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_688),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_662),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_677),
.A2(n_636),
.B1(n_676),
.B2(n_703),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

AOI221xp5_ASAP7_75t_L g731 ( 
.A1(n_637),
.A2(n_701),
.B1(n_636),
.B2(n_626),
.C(n_629),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_657),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_638),
.A2(n_681),
.B1(n_642),
.B2(n_625),
.Y(n_733)
);

OA21x2_ASAP7_75t_L g734 ( 
.A1(n_704),
.A2(n_708),
.B(n_705),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_612),
.A2(n_615),
.B(n_695),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_662),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_666),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_SL g738 ( 
.A1(n_639),
.A2(n_656),
.B1(n_661),
.B2(n_687),
.C(n_683),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_681),
.A2(n_625),
.B1(n_631),
.B2(n_664),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_641),
.B(n_685),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_664),
.A2(n_646),
.B1(n_684),
.B2(n_647),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_651),
.B(n_653),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_643),
.B(n_696),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_661),
.A2(n_680),
.B(n_686),
.C(n_678),
.Y(n_744)
);

OAI221xp5_ASAP7_75t_L g745 ( 
.A1(n_644),
.A2(n_696),
.B1(n_650),
.B2(n_649),
.C(n_615),
.Y(n_745)
);

OAI211xp5_ASAP7_75t_SL g746 ( 
.A1(n_667),
.A2(n_689),
.B(n_644),
.C(n_650),
.Y(n_746)
);

BUFx12f_ASAP7_75t_L g747 ( 
.A(n_640),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_665),
.B(n_621),
.C(n_632),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_669),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_L g750 ( 
.A1(n_655),
.A2(n_663),
.B1(n_668),
.B2(n_617),
.C(n_690),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_668),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_669),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_617),
.A2(n_690),
.B1(n_669),
.B2(n_654),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_634),
.B(n_671),
.Y(n_754)
);

INVx5_ASAP7_75t_SL g755 ( 
.A(n_669),
.Y(n_755)
);

OAI211xp5_ASAP7_75t_SL g756 ( 
.A1(n_617),
.A2(n_456),
.B(n_706),
.C(n_599),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_690),
.A2(n_652),
.B1(n_288),
.B2(n_281),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_690),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_613),
.A2(n_327),
.B1(n_599),
.B2(n_675),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_613),
.A2(n_327),
.B1(n_599),
.B2(n_675),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_628),
.B(n_448),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_691),
.A2(n_288),
.B1(n_281),
.B2(n_285),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_675),
.A2(n_327),
.B1(n_620),
.B2(n_619),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_613),
.A2(n_327),
.B1(n_599),
.B2(n_675),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_691),
.B(n_628),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_675),
.A2(n_327),
.B1(n_620),
.B2(n_619),
.Y(n_766)
);

AOI32xp33_ASAP7_75t_L g767 ( 
.A1(n_691),
.A2(n_450),
.A3(n_231),
.B1(n_242),
.B2(n_274),
.Y(n_767)
);

AND2x4_ASAP7_75t_SL g768 ( 
.A(n_679),
.B(n_534),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_679),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_635),
.B(n_660),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_613),
.A2(n_327),
.B1(n_599),
.B2(n_675),
.Y(n_771)
);

OAI211xp5_ASAP7_75t_SL g772 ( 
.A1(n_706),
.A2(n_456),
.B(n_599),
.C(n_330),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_633),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_613),
.B(n_325),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_742),
.B(n_719),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_749),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_765),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_747),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_743),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_752),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_719),
.B(n_763),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_713),
.B(n_761),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_768),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_770),
.B(n_723),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_734),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_770),
.B(n_723),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_716),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_773),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_732),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_715),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_758),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_711),
.B(n_720),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_763),
.B(n_766),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_766),
.B(n_717),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_729),
.B(n_709),
.Y(n_795)
);

AOI211xp5_ASAP7_75t_L g796 ( 
.A1(n_724),
.A2(n_756),
.B(n_709),
.C(n_772),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_730),
.Y(n_797)
);

OAI33xp33_ASAP7_75t_L g798 ( 
.A1(n_757),
.A2(n_753),
.A3(n_746),
.B1(n_744),
.B2(n_767),
.B3(n_774),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_726),
.B(n_731),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_745),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_731),
.B(n_714),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_751),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_753),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_755),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_769),
.B(n_748),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_755),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_721),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_755),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_759),
.B(n_771),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_793),
.B(n_735),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_785),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_775),
.B(n_725),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_793),
.B(n_741),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_784),
.B(n_764),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_775),
.B(n_725),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_780),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_804),
.Y(n_817)
);

OAI221xp5_ASAP7_75t_L g818 ( 
.A1(n_799),
.A2(n_760),
.B1(n_710),
.B2(n_733),
.C(n_762),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_781),
.B(n_750),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_803),
.B(n_754),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_776),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_791),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_791),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_805),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_806),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_786),
.B(n_722),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_792),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_792),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_779),
.Y(n_829)
);

AOI221xp5_ASAP7_75t_L g830 ( 
.A1(n_818),
.A2(n_798),
.B1(n_799),
.B2(n_782),
.C(n_777),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_810),
.B(n_803),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_814),
.B(n_797),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_818),
.A2(n_781),
.B(n_795),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_810),
.B(n_794),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_821),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_821),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_813),
.B(n_794),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_829),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_829),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_812),
.B(n_800),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_816),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_811),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_841),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_837),
.B(n_822),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_841),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_840),
.B(n_820),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_831),
.B(n_813),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_842),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_838),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_836),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_837),
.B(n_822),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_831),
.B(n_820),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_834),
.B(n_823),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_847),
.B(n_834),
.Y(n_854)
);

AOI32xp33_ASAP7_75t_L g855 ( 
.A1(n_852),
.A2(n_830),
.A3(n_847),
.B1(n_796),
.B2(n_737),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_846),
.B(n_840),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_846),
.B(n_836),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_852),
.B(n_839),
.Y(n_858)
);

OAI32xp33_ASAP7_75t_L g859 ( 
.A1(n_844),
.A2(n_812),
.A3(n_815),
.B1(n_789),
.B2(n_833),
.Y(n_859)
);

AOI222xp33_ASAP7_75t_L g860 ( 
.A1(n_849),
.A2(n_833),
.B1(n_809),
.B2(n_832),
.C1(n_814),
.C2(n_819),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_853),
.B(n_820),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_850),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_850),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_860),
.B(n_851),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_857),
.Y(n_865)
);

NOR3x1_ASAP7_75t_L g866 ( 
.A(n_858),
.B(n_783),
.C(n_815),
.Y(n_866)
);

AOI21xp33_ASAP7_75t_SL g867 ( 
.A1(n_855),
.A2(n_778),
.B(n_783),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_856),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_863),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_861),
.A2(n_819),
.B1(n_796),
.B2(n_809),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_859),
.A2(n_835),
.B(n_790),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_854),
.B(n_848),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_862),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_867),
.A2(n_862),
.B(n_802),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_864),
.B(n_845),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_868),
.A2(n_827),
.B1(n_828),
.B2(n_824),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_865),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_SL g878 ( 
.A1(n_871),
.A2(n_740),
.B(n_808),
.C(n_738),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_872),
.B(n_848),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_875),
.A2(n_870),
.B(n_873),
.Y(n_880)
);

OAI221xp5_ASAP7_75t_SL g881 ( 
.A1(n_874),
.A2(n_865),
.B1(n_866),
.B2(n_727),
.C(n_795),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_879),
.B(n_869),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_877),
.B(n_869),
.Y(n_883)
);

OAI211xp5_ASAP7_75t_L g884 ( 
.A1(n_878),
.A2(n_718),
.B(n_728),
.C(n_736),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_881),
.A2(n_876),
.B(n_801),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_883),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_880),
.B(n_843),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_882),
.B(n_826),
.Y(n_888)
);

OR4x2_ASAP7_75t_L g889 ( 
.A(n_885),
.B(n_712),
.C(n_882),
.D(n_884),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_886),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_SL g891 ( 
.A(n_887),
.B(n_728),
.C(n_739),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_891),
.B(n_888),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_890),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_889),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_893),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_895),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_896),
.A2(n_894),
.B1(n_892),
.B2(n_891),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_897),
.A2(n_894),
.B1(n_825),
.B2(n_817),
.Y(n_898)
);

AOI222xp33_ASAP7_75t_L g899 ( 
.A1(n_898),
.A2(n_807),
.B1(n_787),
.B2(n_797),
.C1(n_788),
.C2(n_802),
.Y(n_899)
);


endmodule