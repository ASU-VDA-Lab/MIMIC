module fake_jpeg_28073_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_29),
.B1(n_34),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_57),
.B1(n_0),
.B2(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_25),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_27),
.B(n_33),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_71),
.C(n_35),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_18),
.B1(n_29),
.B2(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_56),
.B(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_65),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_28),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_25),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_85),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_82),
.B1(n_89),
.B2(n_92),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_40),
.B1(n_21),
.B2(n_35),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_96),
.B1(n_102),
.B2(n_106),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_98),
.B(n_5),
.C(n_6),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_80),
.B(n_91),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_19),
.B1(n_31),
.B2(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_90),
.B1(n_95),
.B2(n_101),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_88),
.Y(n_121)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_19),
.B1(n_31),
.B2(n_17),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_23),
.B1(n_31),
.B2(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_93),
.B(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_23),
.B(n_32),
.C(n_17),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_32),
.B1(n_31),
.B2(n_19),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_15),
.B(n_14),
.C(n_13),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_32),
.B1(n_14),
.B2(n_10),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_32),
.B1(n_14),
.B2(n_10),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_10),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_63),
.C(n_64),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_50),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_104),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_58),
.B1(n_49),
.B2(n_53),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_121),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_58),
.B1(n_53),
.B2(n_66),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_136),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_122),
.B1(n_109),
.B2(n_101),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_66),
.B1(n_48),
.B2(n_5),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_48),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_77),
.B1(n_81),
.B2(n_98),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_79),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_48),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_6),
.C(n_7),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_105),
.C(n_108),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_111),
.B(n_122),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_152),
.B1(n_115),
.B2(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_144),
.B(n_151),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_84),
.B1(n_86),
.B2(n_110),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_84),
.B1(n_86),
.B2(n_100),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_119),
.B1(n_123),
.B2(n_137),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_105),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_97),
.B1(n_90),
.B2(n_108),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_170),
.B(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_97),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_158),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_130),
.C(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_159),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_75),
.CI(n_83),
.CON(n_159),
.SN(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_83),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_7),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_74),
.B1(n_72),
.B2(n_9),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_112),
.B(n_8),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_113),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_136),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_8),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_182),
.B(n_187),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_200),
.C(n_202),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_189),
.B(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_115),
.B1(n_129),
.B2(n_136),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_197),
.B1(n_172),
.B2(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_190),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_127),
.B(n_123),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_192),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_201),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_162),
.B1(n_169),
.B2(n_153),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_145),
.A2(n_172),
.B(n_141),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_180),
.B1(n_179),
.B2(n_183),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_124),
.C(n_119),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_187),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_172),
.B1(n_142),
.B2(n_152),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_221),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_222),
.Y(n_234)
);

XOR2x1_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_143),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_220),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_156),
.C(n_158),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_217),
.C(n_218),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_159),
.B1(n_143),
.B2(n_168),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_215),
.B1(n_223),
.B2(n_187),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_159),
.B1(n_165),
.B2(n_154),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_167),
.C(n_151),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_137),
.C(n_161),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_124),
.C(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_127),
.C(n_170),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_183),
.A3(n_174),
.B1(n_194),
.B2(n_189),
.C1(n_187),
.C2(n_193),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_204),
.C(n_196),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_224),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_179),
.B(n_190),
.C(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_245),
.B1(n_193),
.B2(n_225),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_246),
.B(n_248),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_209),
.B1(n_205),
.B2(n_214),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_186),
.B(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_185),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_220),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_207),
.C(n_212),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_253),
.C(n_265),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_249),
.C(n_237),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_258),
.B1(n_264),
.B2(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_215),
.B1(n_173),
.B2(n_221),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_236),
.B1(n_245),
.B2(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_203),
.B1(n_208),
.B2(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_266),
.B1(n_238),
.B2(n_236),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_217),
.C(n_206),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_227),
.B1(n_181),
.B2(n_165),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_233),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_195),
.B(n_196),
.Y(n_283)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_245),
.B1(n_236),
.B2(n_235),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_238),
.B(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_181),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_178),
.Y(n_288)
);

NAND4xp25_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_259),
.C(n_250),
.D(n_195),
.Y(n_282)
);

OAI21x1_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_291),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_252),
.B(n_265),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_280),
.B(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_253),
.C(n_262),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_276),
.C(n_275),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_178),
.B(n_146),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_291),
.B1(n_283),
.B2(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_268),
.B1(n_271),
.B2(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_298),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_286),
.C(n_290),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_275),
.C(n_279),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_268),
.C(n_270),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_270),
.B1(n_178),
.B2(n_146),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_146),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_293),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_307),
.C(n_302),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_296),
.B(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_303),
.CI(n_301),
.CON(n_309),
.SN(n_309)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_72),
.A3(n_74),
.B1(n_128),
.B2(n_308),
.C1(n_309),
.C2(n_306),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_309),
.B(n_128),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_309),
.Y(n_313)
);


endmodule