module fake_jpeg_22121_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_33),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_62),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_59),
.Y(n_91)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_35),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_46),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_42),
.B1(n_23),
.B2(n_26),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_84),
.B1(n_85),
.B2(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_51),
.Y(n_113)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_43),
.B1(n_23),
.B2(n_36),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_93),
.B1(n_69),
.B2(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_21),
.B1(n_16),
.B2(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_21),
.B1(n_16),
.B2(n_31),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_49),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_88),
.C(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_43),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_21),
.B(n_30),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_94),
.B(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_34),
.B1(n_30),
.B2(n_19),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_57),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_68),
.B1(n_69),
.B2(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_114),
.B1(n_93),
.B2(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_78),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_98),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_79),
.B(n_72),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_110),
.B(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_61),
.B(n_54),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_117),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_34),
.B1(n_25),
.B2(n_19),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_20),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_25),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_20),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_131),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_88),
.B1(n_77),
.B2(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_125),
.B1(n_130),
.B2(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_102),
.B1(n_103),
.B2(n_101),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_127),
.A2(n_113),
.B(n_107),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_74),
.B1(n_73),
.B2(n_84),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_135),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_148),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_156),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_80),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_133),
.B(n_112),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_97),
.B1(n_112),
.B2(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_120),
.B1(n_130),
.B2(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_86),
.C(n_115),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_152),
.C(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_153),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_86),
.C(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_80),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_106),
.CI(n_117),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_128),
.Y(n_155)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_106),
.C(n_118),
.D(n_112),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_125),
.B1(n_127),
.B2(n_126),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_163),
.B1(n_83),
.B2(n_90),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_170),
.C(n_154),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_162),
.B(n_168),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_149),
.C(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_22),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_175),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_154),
.B(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_142),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.C(n_167),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_89),
.B(n_87),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_180),
.B(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_168),
.B1(n_83),
.B2(n_81),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_166),
.A2(n_22),
.B(n_89),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_188),
.B1(n_58),
.B2(n_28),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_170),
.C(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.C(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_180),
.B(n_169),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_159),
.B(n_164),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_187),
.B1(n_174),
.B2(n_178),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_194),
.A3(n_183),
.B1(n_10),
.B2(n_11),
.C1(n_8),
.C2(n_9),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_192),
.B(n_193),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_3),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_3),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_12),
.C1(n_13),
.C2(n_193),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_192),
.B(n_5),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_180),
.B(n_128),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_200),
.A2(n_197),
.B(n_5),
.C(n_7),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.CI(n_199),
.CON(n_204),
.SN(n_204)
);


endmodule