module real_aes_8706_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g503 ( .A1(n_0), .A2(n_167), .B(n_504), .C(n_507), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_1), .B(n_499), .Y(n_508) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g165 ( .A(n_3), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_4), .B(n_168), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_5), .A2(n_467), .B(n_543), .Y(n_542) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_6), .A2(n_175), .B(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_7), .A2(n_35), .B1(n_155), .B2(n_203), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_8), .B(n_175), .Y(n_183) );
AND2x6_ASAP7_75t_L g170 ( .A(n_9), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_10), .A2(n_170), .B(n_472), .C(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_11), .B(n_36), .Y(n_123) );
INVx1_ASAP7_75t_L g149 ( .A(n_12), .Y(n_149) );
INVx1_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_14), .B(n_151), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_15), .B(n_168), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_16), .B(n_142), .Y(n_249) );
AO32x2_ASAP7_75t_L g219 ( .A1(n_17), .A2(n_141), .A3(n_175), .B1(n_194), .B2(n_220), .Y(n_219) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_18), .A2(n_39), .B1(n_126), .B2(n_745), .C1(n_746), .C2(n_748), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_19), .B(n_155), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_20), .B(n_142), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_21), .A2(n_53), .B1(n_155), .B2(n_203), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_22), .A2(n_79), .B1(n_151), .B2(n_155), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_23), .B(n_155), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_24), .A2(n_194), .B(n_472), .C(n_490), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_25), .A2(n_194), .B(n_472), .C(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_26), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_27), .B(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_28), .A2(n_467), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_29), .B(n_196), .Y(n_237) );
INVx2_ASAP7_75t_L g153 ( .A(n_30), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_31), .A2(n_470), .B(n_474), .C(n_480), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_32), .B(n_155), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_33), .B(n_196), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_34), .B(n_214), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_36), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_37), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_38), .Y(n_520) );
INVx1_ASAP7_75t_L g745 ( .A(n_39), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_40), .B(n_168), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_41), .B(n_467), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_42), .A2(n_129), .B1(n_130), .B2(n_451), .Y(n_128) );
INVx1_ASAP7_75t_L g451 ( .A(n_42), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_42), .A2(n_44), .B1(n_451), .B2(n_757), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_43), .A2(n_470), .B(n_480), .C(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_44), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_45), .B(n_155), .Y(n_178) );
INVx1_ASAP7_75t_L g505 ( .A(n_46), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_47), .A2(n_89), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g536 ( .A(n_48), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_49), .B(n_155), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_50), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_51), .B(n_467), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_52), .B(n_163), .Y(n_182) );
AOI22xp33_ASAP7_75t_SL g247 ( .A1(n_54), .A2(n_58), .B1(n_151), .B2(n_155), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_55), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_56), .B(n_155), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_57), .B(n_155), .Y(n_211) );
INVx1_ASAP7_75t_L g171 ( .A(n_59), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_60), .B(n_467), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_61), .B(n_499), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_62), .A2(n_157), .B(n_163), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_63), .B(n_155), .Y(n_166) );
INVx1_ASAP7_75t_L g145 ( .A(n_64), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_66), .B(n_168), .Y(n_478) );
AO32x2_ASAP7_75t_L g200 ( .A1(n_67), .A2(n_175), .A3(n_194), .B1(n_201), .B2(n_206), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_68), .B(n_169), .Y(n_517) );
INVx1_ASAP7_75t_L g190 ( .A(n_69), .Y(n_190) );
INVx1_ASAP7_75t_L g232 ( .A(n_70), .Y(n_232) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_71), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_72), .B(n_477), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_73), .A2(n_472), .B(n_480), .C(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_74), .B(n_151), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_75), .Y(n_544) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_77), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_78), .B(n_476), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_80), .B(n_203), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_81), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_82), .B(n_151), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_83), .A2(n_101), .B1(n_112), .B2(n_758), .Y(n_100) );
INVx2_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_85), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_86), .B(n_193), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_87), .B(n_151), .Y(n_179) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_88), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g454 ( .A(n_88), .B(n_122), .Y(n_454) );
INVx2_ASAP7_75t_L g458 ( .A(n_88), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_90), .A2(n_99), .B1(n_151), .B2(n_152), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_91), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g475 ( .A(n_92), .Y(n_475) );
INVxp67_ASAP7_75t_L g547 ( .A(n_93), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_94), .B(n_151), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g513 ( .A(n_96), .Y(n_513) );
INVx1_ASAP7_75t_L g571 ( .A(n_97), .Y(n_571) );
AND2x2_ASAP7_75t_L g538 ( .A(n_98), .B(n_196), .Y(n_538) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx5_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_104), .Y(n_759) );
OR2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
AND2x2_ASAP7_75t_L g122 ( .A(n_108), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_125), .B1(n_751), .B2(n_753), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g752 ( .A(n_117), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_118), .A2(n_120), .B(n_754), .Y(n_753) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_124), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_121), .B(n_458), .Y(n_750) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g457 ( .A(n_122), .B(n_458), .Y(n_457) );
OAI22x1_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_452), .B1(n_455), .B2(n_459), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_128), .A2(n_452), .B1(n_457), .B2(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_129), .A2(n_130), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_417), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_321), .C(n_405), .Y(n_131) );
NAND4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_264), .C(n_286), .D(n_302), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_197), .B1(n_223), .B2(n_242), .C(n_250), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_173), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_136), .B(n_242), .Y(n_276) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_136), .B(n_304), .C(n_317), .D(n_319), .Y(n_316) );
INVxp67_ASAP7_75t_L g433 ( .A(n_136), .Y(n_433) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g315 ( .A(n_137), .B(n_253), .Y(n_315) );
AND2x2_ASAP7_75t_L g339 ( .A(n_137), .B(n_173), .Y(n_339) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g306 ( .A(n_138), .B(n_241), .Y(n_306) );
AND2x2_ASAP7_75t_L g346 ( .A(n_138), .B(n_327), .Y(n_346) );
AND2x2_ASAP7_75t_L g363 ( .A(n_138), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_138), .B(n_174), .Y(n_387) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g240 ( .A(n_139), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g258 ( .A(n_139), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g270 ( .A(n_139), .B(n_174), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_139), .B(n_184), .Y(n_292) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_147), .B(n_172), .Y(n_139) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_140), .A2(n_185), .B(n_195), .Y(n_184) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_141), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_143), .B(n_144), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_161), .B(n_170), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_157), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_150), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_150), .A2(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g156 ( .A(n_153), .Y(n_156) );
INVx1_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
INVx3_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_155), .Y(n_573) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
AND2x6_ASAP7_75t_L g472 ( .A(n_156), .B(n_473), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_157), .A2(n_571), .B(n_572), .C(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_158), .A2(n_235), .B(n_236), .Y(n_234) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g477 ( .A(n_159), .Y(n_477) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g169 ( .A(n_160), .Y(n_169) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx1_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
AND2x2_ASAP7_75t_L g468 ( .A(n_160), .B(n_164), .Y(n_468) );
INVx1_ASAP7_75t_L g473 ( .A(n_160), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_166), .C(n_167), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g189 ( .A1(n_162), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_162), .A2(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_167), .A2(n_181), .B(n_182), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_167), .A2(n_193), .B1(n_221), .B2(n_222), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_167), .A2(n_193), .B1(n_246), .B2(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_168), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_168), .A2(n_187), .B(n_188), .Y(n_186) );
O2A1O1Ixp5_ASAP7_75t_SL g230 ( .A1(n_168), .A2(n_231), .B(n_232), .C(n_233), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_168), .B(n_547), .Y(n_546) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g201 ( .A1(n_169), .A2(n_193), .B1(n_202), .B2(n_205), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_170), .A2(n_177), .B(n_180), .Y(n_176) );
BUFx3_ASAP7_75t_L g194 ( .A(n_170), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_170), .A2(n_210), .B(n_215), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_170), .A2(n_230), .B(n_234), .Y(n_229) );
AND2x4_ASAP7_75t_L g467 ( .A(n_170), .B(n_468), .Y(n_467) );
INVx4_ASAP7_75t_SL g481 ( .A(n_170), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_170), .B(n_468), .Y(n_514) );
AND2x2_ASAP7_75t_L g273 ( .A(n_173), .B(n_274), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_173), .A2(n_323), .B1(n_326), .B2(n_328), .C(n_332), .Y(n_322) );
AND2x2_ASAP7_75t_L g381 ( .A(n_173), .B(n_346), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_173), .B(n_363), .Y(n_415) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_184), .Y(n_173) );
INVx3_ASAP7_75t_L g241 ( .A(n_174), .Y(n_241) );
AND2x2_ASAP7_75t_L g290 ( .A(n_174), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g344 ( .A(n_174), .B(n_259), .Y(n_344) );
AND2x2_ASAP7_75t_L g402 ( .A(n_174), .B(n_403), .Y(n_402) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_183), .Y(n_174) );
INVx4_ASAP7_75t_L g244 ( .A(n_175), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_175), .A2(n_523), .B(n_524), .Y(n_522) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_175), .Y(n_541) );
AND2x2_ASAP7_75t_L g242 ( .A(n_184), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
INVx1_ASAP7_75t_L g314 ( .A(n_184), .Y(n_314) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_184), .Y(n_320) );
AND2x2_ASAP7_75t_L g365 ( .A(n_184), .B(n_241), .Y(n_365) );
OR2x2_ASAP7_75t_L g404 ( .A(n_184), .B(n_243), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_189), .B(n_194), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_192), .A2(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx4_ASAP7_75t_L g506 ( .A(n_193), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_194), .B(n_244), .C(n_245), .Y(n_263) );
INVx2_ASAP7_75t_L g206 ( .A(n_196), .Y(n_206) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_196), .A2(n_209), .B(n_218), .Y(n_208) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_196), .A2(n_229), .B(n_237), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_196), .A2(n_466), .B(n_469), .Y(n_465) );
INVx1_ASAP7_75t_L g496 ( .A(n_196), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_196), .A2(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_197), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
AND2x2_ASAP7_75t_L g400 ( .A(n_198), .B(n_397), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_198), .B(n_382), .Y(n_432) );
BUFx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g331 ( .A(n_199), .B(n_255), .Y(n_331) );
AND2x2_ASAP7_75t_L g380 ( .A(n_199), .B(n_226), .Y(n_380) );
INVx1_ASAP7_75t_L g426 ( .A(n_199), .Y(n_426) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
AND2x2_ASAP7_75t_L g281 ( .A(n_200), .B(n_255), .Y(n_281) );
INVx1_ASAP7_75t_L g298 ( .A(n_200), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_200), .B(n_219), .Y(n_304) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_204), .Y(n_479) );
INVx2_ASAP7_75t_L g507 ( .A(n_204), .Y(n_507) );
INVx1_ASAP7_75t_L g493 ( .A(n_206), .Y(n_493) );
AND2x2_ASAP7_75t_L g372 ( .A(n_207), .B(n_280), .Y(n_372) );
INVx2_ASAP7_75t_L g437 ( .A(n_207), .Y(n_437) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
AND2x2_ASAP7_75t_L g254 ( .A(n_208), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g267 ( .A(n_208), .B(n_227), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_208), .B(n_226), .Y(n_295) );
INVx1_ASAP7_75t_L g301 ( .A(n_208), .Y(n_301) );
INVx1_ASAP7_75t_L g318 ( .A(n_208), .Y(n_318) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_208), .Y(n_330) );
INVx2_ASAP7_75t_L g398 ( .A(n_208), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g255 ( .A(n_219), .Y(n_255) );
BUFx2_ASAP7_75t_L g352 ( .A(n_219), .Y(n_352) );
AND2x2_ASAP7_75t_L g397 ( .A(n_219), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_238), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_225), .B(n_334), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_225), .A2(n_396), .B(n_410), .Y(n_420) );
AND2x2_ASAP7_75t_L g445 ( .A(n_225), .B(n_331), .Y(n_445) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g367 ( .A(n_227), .Y(n_367) );
AND2x2_ASAP7_75t_L g396 ( .A(n_227), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_228), .Y(n_280) );
INVx2_ASAP7_75t_L g299 ( .A(n_228), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_228), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g253 ( .A(n_239), .Y(n_253) );
OR2x2_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g334 ( .A(n_239), .B(n_330), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_239), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g435 ( .A(n_239), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_239), .B(n_372), .Y(n_447) );
AND2x2_ASAP7_75t_L g326 ( .A(n_240), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g349 ( .A(n_240), .B(n_242), .Y(n_349) );
INVx2_ASAP7_75t_L g261 ( .A(n_241), .Y(n_261) );
AND2x2_ASAP7_75t_L g289 ( .A(n_241), .B(n_262), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_241), .B(n_314), .Y(n_370) );
AND2x2_ASAP7_75t_L g284 ( .A(n_242), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g431 ( .A(n_242), .Y(n_431) );
AND2x2_ASAP7_75t_L g443 ( .A(n_242), .B(n_306), .Y(n_443) );
AND2x2_ASAP7_75t_L g269 ( .A(n_243), .B(n_259), .Y(n_269) );
INVx1_ASAP7_75t_L g364 ( .A(n_243), .Y(n_364) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_248), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_244), .B(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g499 ( .A(n_244), .Y(n_499) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_244), .A2(n_512), .B(n_519), .Y(n_511) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_244), .A2(n_568), .B(n_575), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_244), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g262 ( .A(n_249), .B(n_263), .Y(n_262) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_256), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_253), .B(n_300), .Y(n_309) );
OR2x2_ASAP7_75t_L g441 ( .A(n_253), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g358 ( .A(n_254), .B(n_299), .Y(n_358) );
AND2x2_ASAP7_75t_L g366 ( .A(n_254), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g425 ( .A(n_254), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g449 ( .A(n_254), .B(n_296), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_255), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g436 ( .A(n_255), .B(n_299), .Y(n_436) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x2_ASAP7_75t_L g288 ( .A(n_258), .B(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g450 ( .A(n_258), .Y(n_450) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g285 ( .A(n_261), .Y(n_285) );
AND2x2_ASAP7_75t_L g336 ( .A(n_261), .B(n_269), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_261), .B(n_404), .Y(n_430) );
INVx2_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
INVx3_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
OR2x2_ASAP7_75t_L g355 ( .A(n_262), .B(n_356), .Y(n_355) );
AOI311xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .A3(n_270), .B(n_271), .C(n_282), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_265), .A2(n_303), .B(n_305), .C(n_307), .Y(n_302) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g287 ( .A(n_267), .Y(n_287) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g305 ( .A(n_269), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_269), .B(n_285), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_269), .B(n_270), .Y(n_438) );
AND2x2_ASAP7_75t_L g360 ( .A(n_270), .B(n_274), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_277), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g418 ( .A(n_274), .B(n_306), .Y(n_418) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_275), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g312 ( .A(n_275), .Y(n_312) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g303 ( .A(n_279), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g348 ( .A(n_281), .Y(n_348) );
AND2x4_ASAP7_75t_L g410 ( .A(n_281), .B(n_379), .Y(n_410) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_284), .A2(n_350), .B1(n_362), .B2(n_366), .C1(n_368), .C2(n_372), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_290), .C(n_293), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_287), .B(n_331), .Y(n_354) );
INVx1_ASAP7_75t_L g376 ( .A(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
OR2x2_ASAP7_75t_L g375 ( .A(n_292), .B(n_376), .Y(n_375) );
OAI21xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_300), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g311 ( .A(n_294), .B(n_312), .C(n_313), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_294), .A2(n_331), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_299), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g408 ( .A(n_299), .Y(n_408) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_299), .Y(n_424) );
INVx2_ASAP7_75t_L g382 ( .A(n_300), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_304), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_310), .B1(n_311), .B2(n_315), .C(n_316), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_310), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g444 ( .A(n_310), .Y(n_444) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g325 ( .A(n_317), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_317), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g383 ( .A(n_317), .B(n_331), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_317), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g416 ( .A(n_317), .B(n_351), .Y(n_416) );
BUFx3_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND5xp2_ASAP7_75t_L g321 ( .A(n_322), .B(n_340), .C(n_361), .D(n_373), .E(n_388), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI32xp33_ASAP7_75t_L g413 ( .A1(n_325), .A2(n_352), .A3(n_368), .B1(n_414), .B2(n_416), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_327), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g337 ( .A(n_331), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_353), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g412 ( .A(n_344), .B(n_363), .Y(n_412) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_349), .A2(n_410), .B1(n_428), .B2(n_433), .C(n_434), .Y(n_427) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_L g393 ( .A(n_352), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_357), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g371 ( .A(n_363), .Y(n_371) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_384), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_382), .A2(n_429), .B1(n_431), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B(n_401), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B(n_411), .C(n_413), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_421), .C(n_446), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_418), .Y(n_422) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B(n_427), .C(n_439), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B(n_438), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g747 ( .A(n_459), .Y(n_747) );
OR3x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_659), .C(n_702), .Y(n_459) );
NAND5xp2_ASAP7_75t_L g460 ( .A(n_461), .B(n_586), .C(n_616), .D(n_633), .E(n_648), .Y(n_460) );
AOI221xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_509), .B1(n_549), .B2(n_555), .C(n_559), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_484), .Y(n_462) );
OR2x2_ASAP7_75t_L g564 ( .A(n_463), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g603 ( .A(n_463), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g621 ( .A(n_463), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_463), .B(n_557), .Y(n_638) );
OR2x2_ASAP7_75t_L g650 ( .A(n_463), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_463), .B(n_609), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_463), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_463), .B(n_587), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_463), .B(n_595), .Y(n_701) );
AND2x2_ASAP7_75t_L g733 ( .A(n_463), .B(n_497), .Y(n_733) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_463), .Y(n_741) );
INVx5_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_464), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g561 ( .A(n_464), .B(n_539), .Y(n_561) );
BUFx2_ASAP7_75t_L g583 ( .A(n_464), .Y(n_583) );
AND2x2_ASAP7_75t_L g612 ( .A(n_464), .B(n_485), .Y(n_612) );
AND2x2_ASAP7_75t_L g667 ( .A(n_464), .B(n_565), .Y(n_667) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_482), .Y(n_464) );
BUFx2_ASAP7_75t_L g488 ( .A(n_467), .Y(n_488) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_471), .A2(n_481), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_471), .A2(n_481), .B(n_544), .C(n_545), .Y(n_543) );
INVx5_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_478), .C(n_479), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_476), .A2(n_479), .B(n_536), .C(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_484), .B(n_621), .Y(n_630) );
OAI32xp33_ASAP7_75t_L g644 ( .A1(n_484), .A2(n_580), .A3(n_645), .B1(n_646), .B2(n_647), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_484), .B(n_646), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_484), .B(n_564), .Y(n_687) );
INVx1_ASAP7_75t_SL g716 ( .A(n_484), .Y(n_716) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_484), .B(n_511), .C(n_667), .D(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_497), .Y(n_484) );
INVx5_ASAP7_75t_L g558 ( .A(n_485), .Y(n_558) );
AND2x2_ASAP7_75t_L g587 ( .A(n_485), .B(n_498), .Y(n_587) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_485), .Y(n_666) );
AND2x2_ASAP7_75t_L g736 ( .A(n_485), .B(n_683), .Y(n_736) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_489), .B(n_493), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
AND2x4_ASAP7_75t_L g609 ( .A(n_497), .B(n_558), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_497), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g643 ( .A(n_497), .B(n_565), .Y(n_643) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g557 ( .A(n_498), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g595 ( .A(n_498), .B(n_567), .Y(n_595) );
AND2x2_ASAP7_75t_L g604 ( .A(n_498), .B(n_566), .Y(n_604) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B(n_508), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_509), .A2(n_673), .B1(n_675), .B2(n_677), .C1(n_680), .C2(n_681), .Y(n_672) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_528), .Y(n_509) );
AND2x2_ASAP7_75t_L g605 ( .A(n_510), .B(n_606), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g722 ( .A(n_510), .B(n_583), .C(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
INVx5_ASAP7_75t_SL g554 ( .A(n_511), .Y(n_554) );
OAI322xp33_ASAP7_75t_L g559 ( .A1(n_511), .A2(n_560), .A3(n_562), .B1(n_563), .B2(n_577), .C1(n_580), .C2(n_582), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_511), .B(n_552), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_511), .B(n_540), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
INVx2_ASAP7_75t_L g552 ( .A(n_521), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_521), .B(n_530), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_528), .B(n_590), .Y(n_645) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g624 ( .A(n_529), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_539), .Y(n_529) );
OR2x2_ASAP7_75t_L g553 ( .A(n_530), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_530), .B(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g592 ( .A(n_530), .B(n_540), .Y(n_592) );
AND2x2_ASAP7_75t_L g615 ( .A(n_530), .B(n_552), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_530), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g631 ( .A(n_530), .B(n_590), .Y(n_631) );
AND2x2_ASAP7_75t_L g639 ( .A(n_530), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_530), .B(n_599), .Y(n_689) );
INVx5_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g579 ( .A(n_531), .B(n_554), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_531), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g606 ( .A(n_531), .B(n_540), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_531), .B(n_653), .Y(n_694) );
OR2x2_ASAP7_75t_L g710 ( .A(n_531), .B(n_654), .Y(n_710) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_531), .B(n_671), .Y(n_717) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_531), .Y(n_724) );
OR2x6_ASAP7_75t_L g531 ( .A(n_532), .B(n_538), .Y(n_531) );
AND2x2_ASAP7_75t_L g578 ( .A(n_539), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g628 ( .A(n_539), .B(n_552), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_539), .B(n_554), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_539), .B(n_590), .Y(n_712) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_540), .B(n_554), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_540), .B(n_552), .Y(n_600) );
OR2x2_ASAP7_75t_L g654 ( .A(n_540), .B(n_552), .Y(n_654) );
AND2x2_ASAP7_75t_L g671 ( .A(n_540), .B(n_551), .Y(n_671) );
INVxp67_ASAP7_75t_L g693 ( .A(n_540), .Y(n_693) );
AND2x2_ASAP7_75t_L g720 ( .A(n_540), .B(n_590), .Y(n_720) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_540), .Y(n_727) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_548), .Y(n_540) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_551), .B(n_601), .Y(n_674) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g590 ( .A(n_552), .B(n_554), .Y(n_590) );
OR2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
OR2x2_ASAP7_75t_L g662 ( .A(n_553), .B(n_654), .Y(n_662) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g562 ( .A(n_557), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_557), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g563 ( .A(n_558), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_558), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_558), .B(n_565), .Y(n_597) );
INVx2_ASAP7_75t_L g642 ( .A(n_558), .Y(n_642) );
AND2x2_ASAP7_75t_L g655 ( .A(n_558), .B(n_595), .Y(n_655) );
AND2x2_ASAP7_75t_L g680 ( .A(n_558), .B(n_604), .Y(n_680) );
INVx1_ASAP7_75t_L g632 ( .A(n_563), .Y(n_632) );
INVx2_ASAP7_75t_SL g619 ( .A(n_564), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_565), .Y(n_622) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_566), .Y(n_585) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_L g683 ( .A(n_567), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_574), .Y(n_568) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g652 ( .A(n_579), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g658 ( .A(n_579), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_579), .A2(n_661), .B1(n_663), .B2(n_668), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_579), .B(n_671), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_580), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g614 ( .A(n_581), .Y(n_614) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
OR2x2_ASAP7_75t_L g596 ( .A(n_583), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_583), .B(n_587), .Y(n_647) );
AND2x2_ASAP7_75t_L g670 ( .A(n_583), .B(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g646 ( .A(n_585), .Y(n_646) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_593), .C(n_607), .Y(n_586) );
INVx1_ASAP7_75t_L g610 ( .A(n_587), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g718 ( .A1(n_587), .A2(n_719), .B1(n_721), .B2(n_722), .C(n_725), .Y(n_718) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g737 ( .A(n_590), .Y(n_737) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g686 ( .A(n_592), .B(n_625), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B(n_598), .C(n_602), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OAI32xp33_ASAP7_75t_L g711 ( .A1(n_600), .A2(n_601), .A3(n_664), .B1(n_701), .B2(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
AND2x2_ASAP7_75t_L g743 ( .A(n_603), .B(n_642), .Y(n_743) );
AND2x2_ASAP7_75t_L g690 ( .A(n_604), .B(n_642), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_604), .B(n_612), .Y(n_708) );
AOI31xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_610), .A3(n_611), .B(n_613), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_609), .B(n_621), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_609), .B(n_619), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_609), .A2(n_639), .B1(n_729), .B2(n_732), .C(n_734), .Y(n_728) );
CKINVDCx16_ASAP7_75t_R g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g634 ( .A(n_614), .B(n_635), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_623), .B1(n_626), .B2(n_629), .C1(n_631), .C2(n_632), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g699 ( .A(n_618), .Y(n_699) );
INVx1_ASAP7_75t_L g721 ( .A(n_621), .Y(n_721) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_624), .A2(n_735), .B1(n_737), .B2(n_738), .Y(n_734) );
INVx1_ASAP7_75t_L g640 ( .A(n_625), .Y(n_640) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B1(n_639), .B2(n_641), .C(n_644), .Y(n_633) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g678 ( .A(n_636), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g730 ( .A(n_636), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g705 ( .A(n_641), .Y(n_705) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g669 ( .A(n_642), .Y(n_669) );
INVx1_ASAP7_75t_L g651 ( .A(n_643), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_646), .B(n_733), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B1(n_655), .B2(n_656), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g742 ( .A(n_655), .Y(n_742) );
INVxp33_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_657), .B(n_701), .Y(n_700) );
OAI32xp33_ASAP7_75t_L g691 ( .A1(n_658), .A2(n_692), .A3(n_693), .B1(n_694), .B2(n_695), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_672), .C(n_684), .D(n_696), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NAND2xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_667), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_681), .A2(n_697), .B1(n_714), .B2(n_717), .C(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g732 ( .A(n_683), .B(n_733), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_693), .B(n_724), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_700), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_713), .C(n_728), .D(n_739), .Y(n_702) );
O2A1O1Ixp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B(n_709), .C(n_711), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g744 ( .A(n_731), .Y(n_744) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B(n_744), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
endmodule