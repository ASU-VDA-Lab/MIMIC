module fake_netlist_6_2639_n_2261 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2261);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2261;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_1371;
wire n_383;
wire n_1285;
wire n_873;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1624;
wire n_1124;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1317;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_1767;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_1207;
wire n_683;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1397;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_1303;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_924;
wire n_475;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g361 ( 
.A(n_45),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_197),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_54),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_248),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_252),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_19),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_300),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_33),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_169),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_282),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_88),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_307),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_196),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_247),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_94),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_336),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_238),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_115),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_77),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_16),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_102),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_101),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_214),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_69),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_270),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_44),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_105),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_116),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_293),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_161),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_311),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_358),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_152),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_233),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_134),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_257),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_343),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_172),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_350),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_72),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_181),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_200),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_135),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_189),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_277),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_91),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_16),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_174),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_301),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_299),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_12),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_76),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_310),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_256),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_148),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_58),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_27),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_22),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_260),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_262),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_242),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_188),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_42),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_258),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_268),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_333),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_332),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_30),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_84),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g436 ( 
.A(n_55),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_150),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_226),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_72),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_133),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_88),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_244),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_79),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_109),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_251),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_100),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_212),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_65),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_344),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_356),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_209),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_265),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_55),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_261),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_29),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_198),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_204),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_89),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_229),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_278),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_43),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_14),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_92),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_125),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_329),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_237),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_306),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_354),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_129),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_11),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_58),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_230),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_243),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_295),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_180),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_304),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_309),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_30),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_201),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_118),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_47),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_91),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_193),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_57),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_234),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_297),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_239),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_285),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_246),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_217),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_283),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_206),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_3),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_76),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_302),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_60),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_328),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_71),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_123),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_281),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_357),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_98),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_317),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_253),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_223),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_162),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_353),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_225),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_78),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_179),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_314),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_227),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_177),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_119),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_323),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_46),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_351),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_280),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_218),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_97),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_324),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_275),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_111),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_81),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_112),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_17),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_271),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_32),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_136),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_160),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_34),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_138),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_349),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_70),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_80),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_4),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_340),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_326),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_308),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_286),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_56),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_54),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_48),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_132),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_173),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_166),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_287),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_335),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_73),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_185),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_231),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_236),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_266),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_288),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_8),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_235),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_205),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_352),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_273),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_19),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_59),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_178),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_291),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_67),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_319),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_195),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_4),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_144),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_345),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_182),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_71),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_84),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_215),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_296),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_359),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_87),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_290),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_59),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_274),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_325),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_43),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_149),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_62),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_341),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_318),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_154),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_330),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_294),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_292),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_241),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_339),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_210),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_21),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_232),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_3),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_222),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_216),
.Y(n_598)
);

BUFx5_ASAP7_75t_L g599 ( 
.A(n_86),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_35),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_156),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_183),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_8),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_35),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_312),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_66),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_186),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_272),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_240),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_263),
.Y(n_610)
);

INVxp33_ASAP7_75t_SL g611 ( 
.A(n_5),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_192),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_52),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_316),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_202),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_249),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_220),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_22),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_184),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_38),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_83),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_305),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_27),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_11),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_211),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_34),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_334),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_213),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_42),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_224),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_199),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_167),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_41),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_321),
.Y(n_634)
);

CKINVDCx14_ASAP7_75t_R g635 ( 
.A(n_320),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_303),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_315),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_28),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_110),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_86),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_269),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_327),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_194),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_171),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_95),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_94),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_208),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_190),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_68),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_342),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_355),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_255),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_276),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_203),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_284),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_164),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_176),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_191),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_37),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_347),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_187),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_87),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_289),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_113),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_348),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_130),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_73),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_170),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_47),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_39),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_29),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_64),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_52),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_228),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_207),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_65),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_267),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_81),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_45),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_9),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_221),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_31),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_219),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_41),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_13),
.Y(n_685)
);

BUFx5_ASAP7_75t_L g686 ( 
.A(n_298),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_92),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_250),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_313),
.Y(n_689)
);

BUFx5_ASAP7_75t_L g690 ( 
.A(n_245),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_259),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_279),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_254),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_367),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_436),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_363),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_436),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_436),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_436),
.Y(n_699)
);

CKINVDCx16_ASAP7_75t_R g700 ( 
.A(n_366),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_375),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_454),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_436),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_436),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_599),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_532),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_365),
.Y(n_707)
);

INVxp67_ASAP7_75t_SL g708 ( 
.A(n_649),
.Y(n_708)
);

INVxp33_ASAP7_75t_L g709 ( 
.A(n_382),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_599),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_377),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_679),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_599),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_378),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_599),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_649),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_599),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_372),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_649),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_472),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_599),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_462),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_462),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_649),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_685),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_685),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_685),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_379),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_685),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_386),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_435),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_439),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_497),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_529),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_543),
.Y(n_735)
);

INVxp33_ASAP7_75t_L g736 ( 
.A(n_544),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_562),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_369),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_361),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_565),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_402),
.Y(n_741)
);

INVxp33_ASAP7_75t_SL g742 ( 
.A(n_380),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_568),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_577),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_607),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_381),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_595),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_387),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_579),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_584),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

INVxp33_ASAP7_75t_L g752 ( 
.A(n_603),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_361),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_604),
.Y(n_754)
);

INVxp33_ASAP7_75t_SL g755 ( 
.A(n_388),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_620),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_662),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_389),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_676),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_678),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_424),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_373),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_373),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_493),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_390),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_493),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_408),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_540),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_686),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_540),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_635),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_393),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_424),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_607),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_567),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_567),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_569),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_569),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_664),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_664),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_635),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_674),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_674),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_364),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_495),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_612),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_536),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_368),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_371),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_374),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_536),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_383),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_391),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_537),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_392),
.Y(n_795)
);

INVxp33_ASAP7_75t_SL g796 ( 
.A(n_403),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_537),
.Y(n_797)
);

INVxp33_ASAP7_75t_SL g798 ( 
.A(n_410),
.Y(n_798)
);

CKINVDCx16_ASAP7_75t_R g799 ( 
.A(n_495),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_395),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_396),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_495),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_397),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_405),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_407),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_409),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_417),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_394),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_425),
.Y(n_809)
);

CKINVDCx14_ASAP7_75t_R g810 ( 
.A(n_500),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_406),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_432),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_406),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_486),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_406),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_426),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_612),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_451),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_486),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_453),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_458),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_399),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_460),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_468),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_474),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_471),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_469),
.Y(n_827)
);

INVxp33_ASAP7_75t_SL g828 ( 
.A(n_411),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_473),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_534),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_370),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_477),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_370),
.B(n_0),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_487),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_574),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_621),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_488),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_491),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_385),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_508),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_630),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_513),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_514),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_519),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_400),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_686),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_528),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_545),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_549),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_686),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_686),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_415),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_557),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_630),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_686),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_558),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_560),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_563),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_406),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_564),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_418),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_570),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_581),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_422),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_583),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_509),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_585),
.Y(n_867)
);

BUFx2_ASAP7_75t_SL g868 ( 
.A(n_440),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_376),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_385),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_591),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_401),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_592),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_423),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_404),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_446),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_597),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_602),
.Y(n_878)
);

INVxp33_ASAP7_75t_SL g879 ( 
.A(n_434),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_429),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_605),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_609),
.Y(n_882)
);

INVxp33_ASAP7_75t_SL g883 ( 
.A(n_441),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_622),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_686),
.Y(n_885)
);

INVxp33_ASAP7_75t_L g886 ( 
.A(n_546),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_631),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_636),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_464),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_644),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_647),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_650),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_658),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_661),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_665),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_668),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_484),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_590),
.Y(n_898)
);

INVxp33_ASAP7_75t_SL g899 ( 
.A(n_443),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_677),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_484),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_448),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_688),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_686),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_550),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_693),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_588),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_588),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_653),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_456),
.B(n_0),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_653),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_594),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_691),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_691),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_690),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_416),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_613),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_416),
.Y(n_918)
);

INVxp33_ASAP7_75t_SL g919 ( 
.A(n_459),
.Y(n_919)
);

CKINVDCx16_ASAP7_75t_R g920 ( 
.A(n_687),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_416),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_463),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_416),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_467),
.Y(n_924)
);

CKINVDCx14_ASAP7_75t_R g925 ( 
.A(n_615),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_479),
.Y(n_926)
);

XOR2xp5_ASAP7_75t_L g927 ( 
.A(n_465),
.B(n_1),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_482),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_467),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_467),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_467),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_690),
.Y(n_932)
);

INVxp33_ASAP7_75t_L g933 ( 
.A(n_465),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_506),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_506),
.Y(n_935)
);

BUFx2_ASAP7_75t_SL g936 ( 
.A(n_571),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_506),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_413),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_414),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_506),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_419),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_643),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_643),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_643),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_643),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_483),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_485),
.Y(n_947)
);

INVxp33_ASAP7_75t_SL g948 ( 
.A(n_494),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_362),
.Y(n_949)
);

INVxp33_ASAP7_75t_L g950 ( 
.A(n_611),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_384),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_499),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_510),
.Y(n_953)
);

INVxp33_ASAP7_75t_SL g954 ( 
.A(n_517),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_420),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_421),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_505),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_525),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_427),
.Y(n_959)
);

INVxp33_ASAP7_75t_SL g960 ( 
.A(n_527),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_535),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_542),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_556),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_428),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_398),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_561),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_852),
.B(n_593),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_694),
.B(n_430),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_811),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_724),
.Y(n_970)
);

AND2x6_ASAP7_75t_L g971 ( 
.A(n_695),
.B(n_412),
.Y(n_971)
);

BUFx8_ASAP7_75t_L g972 ( 
.A(n_738),
.Y(n_972)
);

CKINVDCx6p67_ASAP7_75t_R g973 ( 
.A(n_841),
.Y(n_973)
);

INVx6_ASAP7_75t_L g974 ( 
.A(n_745),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_927),
.A2(n_706),
.B1(n_836),
.B2(n_826),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_SL g976 ( 
.A(n_826),
.B(n_572),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_836),
.A2(n_582),
.B1(n_596),
.B2(n_573),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_771),
.B(n_457),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_811),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_700),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_725),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_726),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_708),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_712),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_852),
.B(n_478),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_811),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_933),
.B(n_496),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_874),
.B(n_586),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_815),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_805),
.B(n_639),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_781),
.B(n_431),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_701),
.B(n_433),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_697),
.A2(n_438),
.B(n_437),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_815),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_708),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_727),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_SL g998 ( 
.A1(n_950),
.A2(n_886),
.B1(n_854),
.B2(n_802),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_861),
.B(n_442),
.Y(n_999)
);

OA21x2_ASAP7_75t_L g1000 ( 
.A1(n_698),
.A2(n_445),
.B(n_444),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_859),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_949),
.B(n_606),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_874),
.B(n_447),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_859),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_711),
.B(n_449),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_774),
.Y(n_1006)
);

BUFx8_ASAP7_75t_SL g1007 ( 
.A(n_707),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_716),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_716),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_786),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_714),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_859),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_876),
.B(n_450),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_817),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_825),
.B(n_618),
.Y(n_1015)
);

BUFx8_ASAP7_75t_L g1016 ( 
.A(n_922),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_946),
.B(n_452),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_719),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_813),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_813),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_956),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_813),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_813),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_719),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_729),
.Y(n_1025)
);

BUFx8_ASAP7_75t_SL g1026 ( 
.A(n_741),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_729),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_710),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_728),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_785),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_699),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_SL g1032 ( 
.A1(n_869),
.A2(n_917),
.B1(n_920),
.B2(n_889),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_916),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_964),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_703),
.Y(n_1035)
);

AOI22x1_ASAP7_75t_SL g1036 ( 
.A1(n_767),
.A2(n_624),
.B1(n_626),
.B2(n_623),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_918),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_746),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_921),
.Y(n_1039)
);

BUFx8_ASAP7_75t_SL g1040 ( 
.A(n_812),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_718),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_704),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_748),
.B(n_692),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_861),
.B(n_455),
.Y(n_1044)
);

AO22x1_ASAP7_75t_L g1045 ( 
.A1(n_814),
.A2(n_633),
.B1(n_638),
.B2(n_629),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_923),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_924),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_880),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_758),
.B(n_461),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_905),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_864),
.B(n_466),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_765),
.Y(n_1052)
);

BUFx8_ASAP7_75t_SL g1053 ( 
.A(n_830),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_747),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_705),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_929),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_814),
.B(n_819),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_947),
.B(n_470),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_930),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_772),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_713),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_952),
.B(n_475),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_931),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_934),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_808),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_822),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_935),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_937),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_951),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_953),
.B(n_476),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_696),
.A2(n_645),
.B1(n_646),
.B2(n_640),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_866),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_940),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_833),
.B(n_690),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_912),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_715),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_845),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_942),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_872),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_864),
.B(n_480),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_717),
.A2(n_690),
.B(n_489),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_944),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_721),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_945),
.A2(n_490),
.B(n_481),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_731),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_732),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_733),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_769),
.A2(n_690),
.B(n_498),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_734),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_735),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_737),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_762),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_740),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_875),
.B(n_492),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_846),
.A2(n_690),
.B(n_502),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_743),
.Y(n_1097)
);

BUFx8_ASAP7_75t_SL g1098 ( 
.A(n_835),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_938),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_744),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_850),
.A2(n_690),
.B(n_503),
.Y(n_1101)
);

BUFx8_ASAP7_75t_SL g1102 ( 
.A(n_898),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_939),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_750),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_902),
.B(n_501),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_751),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_754),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_763),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_965),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_756),
.Y(n_1110)
);

BUFx8_ASAP7_75t_SL g1111 ( 
.A(n_941),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_958),
.B(n_504),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_757),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_759),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_955),
.B(n_689),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_959),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_760),
.Y(n_1117)
);

BUFx8_ASAP7_75t_SL g1118 ( 
.A(n_961),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_696),
.A2(n_667),
.B1(n_669),
.B2(n_659),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_851),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_722),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_855),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_723),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_907),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_742),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_885),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_819),
.B(n_507),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_904),
.A2(n_512),
.B(n_511),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_908),
.A2(n_516),
.B(n_515),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_909),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_755),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_902),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_915),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_911),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_868),
.B(n_518),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_926),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_913),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_932),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_739),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_914),
.A2(n_521),
.B(n_520),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_926),
.B(n_522),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_784),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_788),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_789),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_739),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_790),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_936),
.B(n_523),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_910),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_983),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_1041),
.Y(n_1150)
);

INVx6_ASAP7_75t_L g1151 ( 
.A(n_974),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_988),
.B(n_796),
.Y(n_1152)
);

OA21x2_ASAP7_75t_L g1153 ( 
.A1(n_1089),
.A2(n_839),
.B(n_831),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1048),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1081),
.A2(n_793),
.B(n_792),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_969),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_983),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_996),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_995),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_1033),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1007),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1008),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_968),
.B(n_795),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1009),
.B(n_962),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1026),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1009),
.B(n_963),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1018),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1050),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1018),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1024),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_991),
.B(n_928),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1057),
.B(n_957),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1057),
.B(n_798),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1024),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1025),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1075),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1069),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_969),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_SL g1179 ( 
.A1(n_975),
.A2(n_810),
.B1(n_925),
.B2(n_799),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1040),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_1053),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1069),
.B(n_828),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_1098),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1025),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1027),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_974),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1021),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1027),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1121),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1127),
.B(n_879),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1069),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1111),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1029),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1121),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1121),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_967),
.B(n_957),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1096),
.A2(n_801),
.B(n_800),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_969),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_979),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1020),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1123),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1123),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_979),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1109),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1012),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1019),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_967),
.B(n_831),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1142),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1020),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1142),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1109),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1038),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_993),
.B(n_883),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1093),
.B(n_1108),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1144),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1101),
.A2(n_804),
.B(n_803),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_979),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1103),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1144),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_987),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1116),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1005),
.B(n_899),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1144),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1132),
.B(n_928),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1031),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1035),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1109),
.B(n_966),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_987),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1077),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1034),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1139),
.B(n_764),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1043),
.B(n_919),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1020),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_999),
.B(n_839),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1079),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1139),
.B(n_766),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_987),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1032),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1099),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1042),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_990),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1145),
.B(n_768),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1128),
.A2(n_897),
.B(n_870),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1125),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1013),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_990),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1032),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1049),
.B(n_948),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1095),
.B(n_954),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_990),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1131),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1001),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1055),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1001),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1044),
.B(n_870),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_980),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1066),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1061),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1076),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1001),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1051),
.B(n_897),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1011),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1084),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1086),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_984),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1086),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1004),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1011),
.Y(n_1269)
);

AND2x6_ASAP7_75t_L g1270 ( 
.A(n_1074),
.B(n_770),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1052),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_1023),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1004),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1052),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1087),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_976),
.A2(n_671),
.B1(n_672),
.B2(n_670),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1004),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1087),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1091),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1072),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1060),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_976),
.B(n_960),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1054),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1023),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_1148),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1091),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1113),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1113),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1136),
.B(n_775),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1033),
.Y(n_1290)
);

CKINVDCx8_ASAP7_75t_R g1291 ( 
.A(n_1054),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1060),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1102),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1033),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1114),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1145),
.B(n_776),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_985),
.B(n_524),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1054),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1114),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1056),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1065),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1143),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1150),
.B(n_1002),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1235),
.B(n_985),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1149),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1173),
.B(n_989),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1265),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1267),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1227),
.Y(n_1310)
);

NAND2xp33_ASAP7_75t_L g1311 ( 
.A(n_1270),
.B(n_971),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1275),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1278),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1206),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1241),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1151),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1152),
.B(n_1015),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1154),
.B(n_989),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1200),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1254),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1279),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1193),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1172),
.A2(n_971),
.B1(n_901),
.B2(n_994),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1259),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1256),
.B(n_971),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_L g1326 ( 
.A(n_1270),
.B(n_971),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1176),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1200),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1262),
.B(n_1028),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1187),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1286),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1260),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1196),
.A2(n_975),
.B1(n_1119),
.B2(n_702),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1171),
.B(n_1030),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1287),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1264),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1288),
.Y(n_1337)
);

NOR2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1295),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1168),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1215),
.Y(n_1341)
);

INVxp67_ASAP7_75t_SL g1342 ( 
.A(n_1157),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1299),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1225),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1151),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1284),
.Y(n_1346)
);

AND2x6_ASAP7_75t_L g1347 ( 
.A(n_1228),
.B(n_1017),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1302),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1246),
.B(n_1003),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1159),
.Y(n_1350)
);

AND3x2_ASAP7_75t_L g1351 ( 
.A(n_1257),
.B(n_702),
.C(n_1006),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1186),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1158),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1266),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1162),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1209),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1167),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1163),
.B(n_1190),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1213),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1169),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1289),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1284),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1214),
.A2(n_1003),
.B1(n_1105),
.B2(n_1080),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1170),
.A2(n_901),
.B1(n_1000),
.B2(n_994),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1207),
.A2(n_1119),
.B1(n_736),
.B2(n_752),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1174),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1175),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1184),
.B(n_1120),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1185),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1188),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1219),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1160),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1223),
.B(n_1065),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1205),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1284),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1258),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1233),
.B(n_1115),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1231),
.Y(n_1378)
);

OAI21xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1282),
.A2(n_978),
.B(n_1140),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1164),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1163),
.B(n_1017),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1234),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1215),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1166),
.B(n_1122),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1166),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1234),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1249),
.B(n_1058),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1155),
.A2(n_1141),
.B(n_1135),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1218),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1250),
.B(n_1062),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1229),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1297),
.B(n_1070),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1242),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1232),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1270),
.B(n_1138),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1232),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1251),
.Y(n_1397)
);

AND2x6_ASAP7_75t_L g1398 ( 
.A(n_1237),
.B(n_1070),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1253),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1237),
.B(n_1112),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1243),
.B(n_1112),
.Y(n_1401)
);

NAND2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1179),
.B(n_673),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1243),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1268),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1296),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1197),
.A2(n_1217),
.B(n_1210),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1276),
.A2(n_749),
.B1(n_730),
.B2(n_682),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1296),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1160),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1273),
.Y(n_1410)
);

NOR2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1271),
.B(n_973),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1277),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1280),
.B(n_1010),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1290),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1300),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1274),
.B(n_1147),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1156),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1208),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1156),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1156),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1178),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1270),
.B(n_1000),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1211),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1216),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1178),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1281),
.B(n_992),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1220),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1224),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1178),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1177),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1222),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1198),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1204),
.Y(n_1434)
);

BUFx10_ASAP7_75t_L g1435 ( 
.A(n_1192),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1353),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1377),
.B(n_1292),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1390),
.B(n_1363),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1304),
.B(n_1301),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1390),
.B(n_1245),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1366),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1377),
.B(n_1252),
.Y(n_1442)
);

NAND2xp33_ASAP7_75t_L g1443 ( 
.A(n_1347),
.B(n_1212),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1305),
.B(n_1189),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1327),
.B(n_1191),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1325),
.B(n_1276),
.C(n_1129),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1369),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1334),
.B(n_1014),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1305),
.B(n_1194),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1342),
.B(n_1195),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1370),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1373),
.B(n_1182),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1304),
.B(n_1291),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1308),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1309),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1338),
.B(n_1283),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_L g1457 ( 
.A(n_1347),
.B(n_1198),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1312),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1342),
.B(n_1201),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1307),
.B(n_1298),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1318),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1367),
.B(n_1202),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1344),
.B(n_1230),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1344),
.B(n_1236),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1313),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1346),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1321),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1331),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1307),
.B(n_1240),
.Y(n_1469)
);

AOI22x1_ASAP7_75t_SL g1470 ( 
.A1(n_1322),
.A2(n_1248),
.B1(n_1239),
.B2(n_1165),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1367),
.B(n_1129),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1329),
.B(n_1045),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1329),
.B(n_1085),
.Y(n_1473)
);

NAND2xp33_ASAP7_75t_L g1474 ( 
.A(n_1347),
.B(n_1198),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1358),
.B(n_1285),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1358),
.B(n_1285),
.Y(n_1476)
);

NOR2xp67_ASAP7_75t_L g1477 ( 
.A(n_1359),
.B(n_1161),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1335),
.Y(n_1478)
);

BUFx2_ASAP7_75t_R g1479 ( 
.A(n_1371),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1317),
.B(n_972),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1317),
.B(n_972),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1355),
.B(n_1272),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1357),
.B(n_1126),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1360),
.B(n_1126),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1337),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1346),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1339),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1343),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1368),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1368),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1325),
.B(n_1133),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1384),
.B(n_1361),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1384),
.B(n_1133),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1387),
.B(n_998),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1303),
.B(n_1180),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1413),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1361),
.B(n_1244),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_SL g1498 ( 
.A(n_1376),
.B(n_977),
.C(n_1293),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1380),
.B(n_1244),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1385),
.B(n_1199),
.Y(n_1500)
);

BUFx5_ASAP7_75t_L g1501 ( 
.A(n_1347),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1354),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1340),
.B(n_1016),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1349),
.B(n_1118),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1431),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1392),
.A2(n_1400),
.B(n_1401),
.C(n_1379),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1349),
.B(n_1400),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1434),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1433),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1401),
.B(n_1016),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1394),
.Y(n_1511)
);

NOR2xp67_ASAP7_75t_L g1512 ( 
.A(n_1432),
.B(n_1392),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1347),
.B(n_1199),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1396),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1323),
.B(n_1153),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1323),
.B(n_1199),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1403),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1427),
.B(n_1181),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1398),
.B(n_1203),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1378),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1398),
.B(n_1203),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1405),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1314),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1398),
.B(n_1203),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1346),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1311),
.B(n_1153),
.C(n_1074),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1326),
.B(n_1046),
.C(n_1039),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1316),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1398),
.B(n_1221),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1333),
.A2(n_807),
.B1(n_809),
.B2(n_806),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1306),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1437),
.B(n_1417),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1502),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1528),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_L g1535 ( 
.A(n_1477),
.B(n_1330),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1458),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1492),
.B(n_1376),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1448),
.Y(n_1538)
);

AO22x2_ASAP7_75t_L g1539 ( 
.A1(n_1438),
.A2(n_1407),
.B1(n_1036),
.B2(n_1071),
.Y(n_1539)
);

AO22x2_ASAP7_75t_L g1540 ( 
.A1(n_1480),
.A2(n_1407),
.B1(n_1071),
.B2(n_1333),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1467),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1454),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1506),
.A2(n_1364),
.B1(n_1381),
.B2(n_1433),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1455),
.Y(n_1544)
);

AO22x2_ASAP7_75t_L g1545 ( 
.A1(n_1481),
.A2(n_977),
.B1(n_1423),
.B2(n_1427),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1465),
.Y(n_1546)
);

AND2x6_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1423),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1452),
.A2(n_1381),
.B1(n_1398),
.B2(n_1417),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1468),
.Y(n_1549)
);

AO22x2_ASAP7_75t_L g1550 ( 
.A1(n_1446),
.A2(n_1408),
.B1(n_1383),
.B2(n_1341),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1466),
.B(n_1345),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1490),
.B(n_1365),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1466),
.B(n_1352),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1478),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1485),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1461),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1487),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1439),
.B(n_1365),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1488),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1496),
.B(n_1411),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1439),
.B(n_1310),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1445),
.B(n_1505),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1514),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1517),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1472),
.B(n_1315),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1494),
.A2(n_1320),
.B1(n_1332),
.B2(n_1324),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1436),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1442),
.B(n_1336),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1441),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1451),
.B(n_1348),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1440),
.B(n_1183),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1445),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1447),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1507),
.B(n_1419),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1528),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1444),
.Y(n_1578)
);

OAI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1475),
.A2(n_684),
.B1(n_680),
.B2(n_720),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1449),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1508),
.Y(n_1581)
);

AO22x2_ASAP7_75t_L g1582 ( 
.A1(n_1446),
.A2(n_1402),
.B1(n_1425),
.B2(n_1424),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_L g1583 ( 
.A(n_1501),
.B(n_1466),
.Y(n_1583)
);

AO22x2_ASAP7_75t_L g1584 ( 
.A1(n_1476),
.A2(n_1510),
.B1(n_1498),
.B2(n_1453),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1470),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1486),
.B(n_1372),
.Y(n_1586)
);

AO22x2_ASAP7_75t_L g1587 ( 
.A1(n_1516),
.A2(n_1429),
.B1(n_1428),
.B2(n_1395),
.Y(n_1587)
);

BUFx8_ASAP7_75t_L g1588 ( 
.A(n_1531),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1450),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1460),
.B(n_1435),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1543),
.A2(n_1515),
.B(n_1474),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1583),
.A2(n_1515),
.B(n_1457),
.Y(n_1593)
);

AOI33xp33_ASAP7_75t_L g1594 ( 
.A1(n_1570),
.A2(n_1530),
.A3(n_1351),
.B1(n_1110),
.B2(n_1097),
.B3(n_1117),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1578),
.B(n_1509),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1537),
.B(n_1495),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1536),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1548),
.A2(n_1443),
.B(n_1473),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1580),
.A2(n_1471),
.B(n_1526),
.Y(n_1600)
);

AO22x1_ASAP7_75t_L g1601 ( 
.A1(n_1588),
.A2(n_1504),
.B1(n_1518),
.B2(n_1520),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1532),
.B(n_1463),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1558),
.B(n_1445),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1541),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1559),
.B(n_1523),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1590),
.A2(n_1464),
.B1(n_1469),
.B2(n_1456),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1538),
.B(n_1486),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1560),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1589),
.B(n_1497),
.Y(n_1609)
);

NOR3xp33_ASAP7_75t_L g1610 ( 
.A(n_1579),
.B(n_1503),
.C(n_720),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1562),
.A2(n_1526),
.B(n_1409),
.Y(n_1611)
);

OR2x6_ASAP7_75t_SL g1612 ( 
.A(n_1552),
.B(n_1500),
.Y(n_1612)
);

AOI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1587),
.A2(n_1491),
.B(n_1499),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1540),
.B(n_1479),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1586),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1459),
.Y(n_1616)
);

NOR2x1_ASAP7_75t_L g1617 ( 
.A(n_1535),
.B(n_1527),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1556),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1573),
.B(n_1435),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1576),
.A2(n_1527),
.B(n_1493),
.C(n_1482),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1550),
.A2(n_1513),
.B(n_1519),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1572),
.B(n_1486),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1581),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1574),
.B(n_1374),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1571),
.A2(n_1483),
.B(n_1484),
.C(n_1462),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1547),
.B(n_1364),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1564),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1540),
.A2(n_1388),
.B(n_1406),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1550),
.A2(n_1524),
.B(n_1521),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1592),
.A2(n_1547),
.B(n_1567),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1598),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1591),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1599),
.A2(n_1582),
.B(n_1529),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1610),
.A2(n_1563),
.B(n_730),
.C(n_749),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1602),
.A2(n_1563),
.B(n_1544),
.C(n_1546),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1594),
.A2(n_1542),
.B(n_1554),
.C(n_1549),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1618),
.B(n_1557),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1619),
.A2(n_1584),
.B1(n_1539),
.B2(n_1561),
.Y(n_1641)
);

OAI22x1_ASAP7_75t_L g1642 ( 
.A1(n_1606),
.A2(n_1614),
.B1(n_1617),
.B2(n_1603),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1584),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1612),
.B(n_1575),
.Y(n_1645)
);

BUFx8_ASAP7_75t_L g1646 ( 
.A(n_1624),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1628),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1605),
.B(n_1545),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1598),
.B(n_1588),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1595),
.A2(n_1539),
.B1(n_1545),
.B2(n_1623),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1600),
.A2(n_1582),
.B(n_1388),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1611),
.A2(n_1406),
.B(n_1525),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1605),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1593),
.A2(n_1525),
.B(n_1501),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1608),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1601),
.B(n_1568),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1595),
.A2(n_1569),
.B1(n_1565),
.B2(n_1553),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1625),
.A2(n_1630),
.B(n_1621),
.C(n_1620),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1551),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1609),
.B(n_1351),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1350),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1613),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1615),
.B(n_1534),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1626),
.A2(n_1501),
.B(n_1395),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1607),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1622),
.B(n_1094),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1615),
.B(n_1577),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1627),
.Y(n_1668)
);

AND2x6_ASAP7_75t_SL g1669 ( 
.A(n_1627),
.B(n_1585),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_1420),
.B1(n_1421),
.B2(n_1418),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1629),
.A2(n_709),
.B1(n_761),
.B2(n_753),
.Y(n_1671)
);

NAND3x1_ASAP7_75t_L g1672 ( 
.A(n_1641),
.B(n_778),
.C(n_777),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1636),
.B(n_1629),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1658),
.A2(n_1501),
.B(n_1362),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1650),
.A2(n_1635),
.B1(n_1644),
.B2(n_1645),
.C(n_1660),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1652),
.A2(n_1501),
.B(n_1362),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1654),
.A2(n_1651),
.B(n_1634),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1655),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1649),
.B(n_1422),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1633),
.B(n_1094),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1671),
.A2(n_1415),
.B(n_1414),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1637),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_R g1683 ( 
.A(n_1667),
.B(n_1399),
.Y(n_1683)
);

CKINVDCx16_ASAP7_75t_R g1684 ( 
.A(n_1667),
.Y(n_1684)
);

O2A1O1Ixp5_ASAP7_75t_SL g1685 ( 
.A1(n_1657),
.A2(n_818),
.B(n_820),
.C(n_816),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1631),
.A2(n_1391),
.B(n_1389),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1656),
.A2(n_1362),
.B(n_1346),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1663),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1664),
.A2(n_1375),
.B(n_1362),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1663),
.Y(n_1690)
);

AO22x1_ASAP7_75t_L g1691 ( 
.A1(n_1646),
.A2(n_761),
.B1(n_753),
.B2(n_530),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1659),
.B(n_779),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1638),
.B(n_1632),
.C(n_1639),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1640),
.B(n_782),
.C(n_780),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1662),
.A2(n_1375),
.B(n_1328),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1648),
.B(n_1393),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1632),
.Y(n_1698)
);

NOR2xp67_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1397),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1642),
.A2(n_1092),
.B1(n_1106),
.B2(n_783),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1404),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1647),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1670),
.A2(n_1375),
.B(n_1356),
.Y(n_1703)
);

AO31x2_ASAP7_75t_L g1704 ( 
.A1(n_1666),
.A2(n_823),
.A3(n_824),
.B(n_821),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1653),
.A2(n_1416),
.B(n_1356),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1653),
.B(n_1410),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1646),
.Y(n_1707)
);

AO32x2_ASAP7_75t_L g1708 ( 
.A1(n_1669),
.A2(n_5),
.A3(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1665),
.B(n_1146),
.Y(n_1709)
);

AO21x1_ASAP7_75t_L g1710 ( 
.A1(n_1650),
.A2(n_829),
.B(n_827),
.Y(n_1710)
);

AOI211x1_ASAP7_75t_L g1711 ( 
.A1(n_1660),
.A2(n_834),
.B(n_837),
.C(n_832),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1636),
.B(n_1399),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1682),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1675),
.B(n_970),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1673),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1695),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1684),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1677),
.A2(n_787),
.B(n_773),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1678),
.B(n_773),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1674),
.A2(n_1319),
.B(n_1412),
.Y(n_1720)
);

NAND2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1688),
.B(n_1426),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1693),
.A2(n_840),
.B1(n_842),
.B2(n_838),
.Y(n_1722)
);

CKINVDCx12_ASAP7_75t_R g1723 ( 
.A(n_1679),
.Y(n_1723)
);

OA21x2_ASAP7_75t_L g1724 ( 
.A1(n_1696),
.A2(n_791),
.B(n_787),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1702),
.B(n_1697),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1701),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1676),
.A2(n_1386),
.B(n_1382),
.Y(n_1728)
);

AOI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1710),
.A2(n_844),
.B(n_843),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_SL g1730 ( 
.A1(n_1712),
.A2(n_1430),
.B(n_847),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1704),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1699),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1698),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1692),
.A2(n_794),
.B(n_797),
.C(n_791),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1704),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1694),
.A2(n_849),
.B(n_853),
.C(n_848),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1704),
.Y(n_1737)
);

INVx6_ASAP7_75t_L g1738 ( 
.A(n_1690),
.Y(n_1738)
);

AO21x2_ASAP7_75t_L g1739 ( 
.A1(n_1687),
.A2(n_857),
.B(n_856),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1705),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1685),
.A2(n_1046),
.B(n_1039),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1707),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1689),
.A2(n_1067),
.B(n_1064),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1708),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_2),
.Y(n_1745)
);

AND2x2_ASAP7_75t_SL g1746 ( 
.A(n_1708),
.B(n_858),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1679),
.B(n_1124),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_794),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1680),
.B(n_526),
.Y(n_1749)
);

AO21x2_ASAP7_75t_L g1750 ( 
.A1(n_1683),
.A2(n_862),
.B(n_860),
.Y(n_1750)
);

AOI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1691),
.A2(n_1681),
.B(n_1706),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1708),
.B(n_1686),
.Y(n_1752)
);

AO31x2_ASAP7_75t_L g1753 ( 
.A1(n_1703),
.A2(n_865),
.A3(n_867),
.B(n_863),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1711),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1672),
.Y(n_1755)
);

OAI21x1_ASAP7_75t_L g1756 ( 
.A1(n_1677),
.A2(n_1067),
.B(n_1064),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1707),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1675),
.B(n_981),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1682),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1672),
.A2(n_873),
.B(n_871),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1672),
.A2(n_878),
.B(n_877),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1684),
.A2(n_797),
.B1(n_882),
.B2(n_881),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1682),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_SL g1764 ( 
.A(n_1683),
.B(n_531),
.Y(n_1764)
);

NAND2x1p5_ASAP7_75t_L g1765 ( 
.A(n_1688),
.B(n_1221),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1684),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1678),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1682),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1672),
.A2(n_887),
.B(n_884),
.Y(n_1769)
);

BUFx5_ASAP7_75t_L g1770 ( 
.A(n_1678),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1684),
.A2(n_890),
.B1(n_891),
.B2(n_888),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1682),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1682),
.Y(n_1773)
);

OAI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1756),
.A2(n_1083),
.B(n_1073),
.Y(n_1774)
);

INVx6_ASAP7_75t_L g1775 ( 
.A(n_1738),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1713),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1713),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1716),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1716),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1759),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1759),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1726),
.B(n_892),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1738),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1722),
.A2(n_894),
.B(n_893),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1763),
.Y(n_1785)
);

CKINVDCx14_ASAP7_75t_R g1786 ( 
.A(n_1717),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1715),
.B(n_895),
.Y(n_1787)
);

BUFx2_ASAP7_75t_R g1788 ( 
.A(n_1766),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1767),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1763),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1768),
.Y(n_1791)
);

BUFx8_ASAP7_75t_SL g1792 ( 
.A(n_1742),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1768),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1773),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1772),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1772),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1726),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1770),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1770),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1746),
.A2(n_900),
.B1(n_903),
.B2(n_896),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1725),
.B(n_906),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1770),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1757),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1755),
.A2(n_538),
.B1(n_539),
.B2(n_533),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1727),
.B(n_982),
.Y(n_1805)
);

BUFx4f_ASAP7_75t_SL g1806 ( 
.A(n_1748),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1770),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1733),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1731),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1770),
.Y(n_1810)
);

BUFx12f_ASAP7_75t_L g1811 ( 
.A(n_1719),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1740),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1735),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1737),
.Y(n_1814)
);

INVx4_ASAP7_75t_L g1815 ( 
.A(n_1747),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1755),
.B(n_6),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1754),
.A2(n_547),
.B1(n_548),
.B2(n_541),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1744),
.Y(n_1818)
);

AOI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1751),
.A2(n_997),
.B(n_1124),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1752),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1732),
.Y(n_1821)
);

OAI22x1_ASAP7_75t_SL g1822 ( 
.A1(n_1803),
.A2(n_1723),
.B1(n_552),
.B2(n_553),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1806),
.A2(n_1745),
.B1(n_1730),
.B2(n_1749),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1806),
.A2(n_1758),
.B1(n_1714),
.B2(n_1750),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1808),
.Y(n_1825)
);

OAI222xp33_ASAP7_75t_L g1826 ( 
.A1(n_1800),
.A2(n_1747),
.B1(n_1771),
.B2(n_1762),
.C1(n_1765),
.C2(n_1721),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1792),
.Y(n_1827)
);

BUFx12f_ASAP7_75t_L g1828 ( 
.A(n_1782),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1811),
.A2(n_1764),
.B1(n_1729),
.B2(n_1739),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1792),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1800),
.A2(n_1761),
.B1(n_1769),
.B2(n_1760),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1820),
.B(n_1718),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1779),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1787),
.B(n_1718),
.C(n_1734),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1786),
.B(n_1736),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1797),
.A2(n_1724),
.B1(n_1741),
.B2(n_1743),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1786),
.A2(n_1724),
.B1(n_1728),
.B2(n_1720),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1815),
.A2(n_554),
.B1(n_555),
.B2(n_551),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1779),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1791),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1791),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1815),
.A2(n_566),
.B1(n_575),
.B2(n_559),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1804),
.A2(n_578),
.B(n_576),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1787),
.A2(n_587),
.B1(n_589),
.B2(n_580),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1817),
.A2(n_601),
.B(n_598),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1776),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1777),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1821),
.A2(n_610),
.B(n_608),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1778),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1818),
.B(n_1753),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1802),
.B(n_1807),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_R g1852 ( 
.A(n_1827),
.B(n_1775),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1808),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_R g1854 ( 
.A(n_1827),
.B(n_1775),
.Y(n_1854)
);

BUFx12f_ASAP7_75t_L g1855 ( 
.A(n_1830),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1825),
.B(n_1808),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1828),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_R g1858 ( 
.A(n_1830),
.B(n_1775),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1825),
.B(n_1808),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1847),
.B(n_1794),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_R g1861 ( 
.A(n_1828),
.B(n_1788),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1833),
.B(n_1780),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1841),
.B(n_1781),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1847),
.B(n_1849),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1839),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1839),
.B(n_1840),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1835),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1849),
.B(n_1789),
.Y(n_1868)
);

OR2x6_ASAP7_75t_L g1869 ( 
.A(n_1834),
.B(n_1783),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1846),
.B(n_1785),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1840),
.B(n_1790),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1846),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1832),
.B(n_1793),
.Y(n_1873)
);

NAND2xp33_ASAP7_75t_R g1874 ( 
.A(n_1851),
.B(n_1816),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1851),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1850),
.B(n_1795),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1852),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1873),
.B(n_1832),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1876),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1876),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1875),
.B(n_1850),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1862),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1856),
.B(n_1859),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1866),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1866),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1855),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1869),
.B(n_1801),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1869),
.B(n_1853),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1853),
.B(n_1783),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1872),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1857),
.B(n_1783),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1865),
.B(n_1796),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1865),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1867),
.Y(n_1894)
);

INVxp67_ASAP7_75t_SL g1895 ( 
.A(n_1874),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1864),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1862),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1863),
.B(n_1783),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1871),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1863),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1854),
.B(n_1809),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1858),
.B(n_1861),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1870),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1860),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1868),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1852),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1876),
.B(n_1809),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1876),
.B(n_1798),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1893),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1883),
.B(n_1788),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1894),
.Y(n_1911)
);

AND2x4_ASAP7_75t_SL g1912 ( 
.A(n_1894),
.B(n_1823),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1893),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1895),
.B(n_1805),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1894),
.Y(n_1915)
);

NAND2x1_ASAP7_75t_L g1916 ( 
.A(n_1900),
.B(n_1799),
.Y(n_1916)
);

INVx5_ASAP7_75t_L g1917 ( 
.A(n_1886),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1894),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1896),
.B(n_1813),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1899),
.B(n_1824),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1883),
.B(n_1810),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1892),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1892),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1904),
.B(n_1814),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1890),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1890),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1905),
.B(n_1812),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1905),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1894),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1889),
.B(n_1829),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1914),
.B(n_1882),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1929),
.B(n_1906),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1910),
.B(n_1906),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1909),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1917),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1917),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1928),
.B(n_1903),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1929),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1930),
.B(n_1902),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1913),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1920),
.B(n_1878),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1917),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1917),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1922),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1911),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1923),
.B(n_1903),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1931),
.B(n_1915),
.Y(n_1947)
);

AND2x4_ASAP7_75t_SL g1948 ( 
.A(n_1932),
.B(n_1886),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1933),
.B(n_1902),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1932),
.B(n_1918),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1938),
.Y(n_1951)
);

AND2x4_ASAP7_75t_SL g1952 ( 
.A(n_1939),
.B(n_1886),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1935),
.B(n_1877),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1936),
.B(n_1877),
.Y(n_1954)
);

NAND2x1_ASAP7_75t_L g1955 ( 
.A(n_1943),
.B(n_1888),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1951),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1948),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1949),
.B(n_1912),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1952),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1953),
.B(n_1942),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1947),
.Y(n_1961)
);

NOR2xp67_ASAP7_75t_L g1962 ( 
.A(n_1950),
.B(n_1943),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1961),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1956),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1960),
.B(n_1955),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1962),
.B(n_1954),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1962),
.Y(n_1967)
);

AOI21xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1966),
.A2(n_1965),
.B(n_1957),
.Y(n_1968)
);

XNOR2xp5_ASAP7_75t_L g1969 ( 
.A(n_1963),
.B(n_1958),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1967),
.B(n_1957),
.Y(n_1970)
);

XNOR2xp5_ASAP7_75t_L g1971 ( 
.A(n_1969),
.B(n_1959),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1970),
.A2(n_1955),
.B(n_1964),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1971),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1972),
.B(n_1944),
.Y(n_1974)
);

NOR2x1_ASAP7_75t_L g1975 ( 
.A(n_1973),
.B(n_1886),
.Y(n_1975)
);

NOR3x1_ASAP7_75t_L g1976 ( 
.A(n_1974),
.B(n_1968),
.C(n_1940),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1975),
.B(n_1886),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1976),
.B(n_1945),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1975),
.B(n_1945),
.C(n_1934),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1977),
.A2(n_1946),
.B(n_1941),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1979),
.A2(n_1946),
.B1(n_1937),
.B2(n_1925),
.C(n_1926),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1978),
.A2(n_1937),
.B1(n_1891),
.B2(n_1822),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1977),
.A2(n_1891),
.B1(n_1888),
.B2(n_1901),
.Y(n_1983)
);

AOI21x1_ASAP7_75t_L g1984 ( 
.A1(n_1980),
.A2(n_1916),
.B(n_1887),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_SL g1985 ( 
.A1(n_1983),
.A2(n_1900),
.B(n_1885),
.Y(n_1985)
);

O2A1O1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1981),
.A2(n_1843),
.B(n_1838),
.C(n_1842),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1984),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1985),
.Y(n_1988)
);

NAND4xp25_ASAP7_75t_L g1989 ( 
.A(n_1986),
.B(n_1982),
.C(n_1844),
.D(n_1845),
.Y(n_1989)
);

NOR2x1_ASAP7_75t_L g1990 ( 
.A(n_1986),
.B(n_1784),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1985),
.A2(n_1924),
.B(n_1919),
.Y(n_1991)
);

NOR2xp67_ASAP7_75t_L g1992 ( 
.A(n_1985),
.B(n_7),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1985),
.B(n_1090),
.C(n_1088),
.Y(n_1993)
);

NOR3x2_ASAP7_75t_L g1994 ( 
.A(n_1985),
.B(n_7),
.C(n_9),
.Y(n_1994)
);

INVx2_ASAP7_75t_SL g1995 ( 
.A(n_1985),
.Y(n_1995)
);

NAND3xp33_ASAP7_75t_L g1996 ( 
.A(n_1985),
.B(n_1090),
.C(n_1088),
.Y(n_1996)
);

NAND3xp33_ASAP7_75t_L g1997 ( 
.A(n_1985),
.B(n_1090),
.C(n_1088),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1985),
.B(n_1900),
.Y(n_1998)
);

AND4x2_ASAP7_75t_L g1999 ( 
.A(n_1985),
.B(n_13),
.C(n_10),
.D(n_12),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1994),
.Y(n_2000)
);

NOR2x1_ASAP7_75t_L g2001 ( 
.A(n_1988),
.B(n_1100),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1995),
.Y(n_2002)
);

NOR2x1_ASAP7_75t_L g2003 ( 
.A(n_1987),
.B(n_1100),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1992),
.A2(n_1998),
.B(n_1996),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1989),
.B(n_1990),
.Y(n_2005)
);

NOR2x1_ASAP7_75t_SL g2006 ( 
.A(n_1993),
.B(n_1901),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1999),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1991),
.B(n_1884),
.Y(n_2008)
);

NAND2x1p5_ASAP7_75t_L g2009 ( 
.A(n_1997),
.B(n_1100),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_R g2010 ( 
.A(n_1995),
.B(n_10),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1988),
.B(n_1104),
.Y(n_2011)
);

NOR3x2_ASAP7_75t_L g2012 ( 
.A(n_1999),
.B(n_14),
.C(n_15),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_SL g2013 ( 
.A(n_1992),
.B(n_1884),
.Y(n_2013)
);

NOR3x1_ASAP7_75t_L g2014 ( 
.A(n_1988),
.B(n_1848),
.C(n_1919),
.Y(n_2014)
);

NOR3x1_ASAP7_75t_L g2015 ( 
.A(n_1988),
.B(n_1924),
.C(n_1927),
.Y(n_2015)
);

NOR2xp67_ASAP7_75t_L g2016 ( 
.A(n_1995),
.B(n_15),
.Y(n_2016)
);

OAI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1998),
.A2(n_1885),
.B(n_1897),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1998),
.B(n_1897),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1998),
.B(n_1898),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1998),
.B(n_1889),
.Y(n_2020)
);

NOR2x1_ASAP7_75t_L g2021 ( 
.A(n_1988),
.B(n_1104),
.Y(n_2021)
);

NOR2x1_ASAP7_75t_L g2022 ( 
.A(n_1988),
.B(n_1104),
.Y(n_2022)
);

NOR2x1_ASAP7_75t_L g2023 ( 
.A(n_1988),
.B(n_1107),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1998),
.B(n_1898),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1998),
.B(n_1879),
.Y(n_2025)
);

NOR2xp67_ASAP7_75t_L g2026 ( 
.A(n_1995),
.B(n_17),
.Y(n_2026)
);

NOR2x1p5_ASAP7_75t_L g2027 ( 
.A(n_1989),
.B(n_1107),
.Y(n_2027)
);

OAI21xp33_ASAP7_75t_SL g2028 ( 
.A1(n_1992),
.A2(n_1921),
.B(n_1880),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1998),
.B(n_1879),
.Y(n_2029)
);

NAND4xp75_ASAP7_75t_L g2030 ( 
.A(n_1992),
.B(n_21),
.C(n_18),
.D(n_20),
.Y(n_2030)
);

AND2x2_ASAP7_75t_SL g2031 ( 
.A(n_1988),
.B(n_1107),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1992),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_L g2033 ( 
.A(n_1988),
.B(n_616),
.C(n_614),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1999),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1999),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_L g2036 ( 
.A(n_1988),
.B(n_18),
.Y(n_2036)
);

OAI21xp33_ASAP7_75t_L g2037 ( 
.A1(n_1998),
.A2(n_1880),
.B(n_1881),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_1988),
.B(n_20),
.Y(n_2038)
);

NAND4xp25_ASAP7_75t_L g2039 ( 
.A(n_2020),
.B(n_1831),
.C(n_25),
.D(n_23),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_L g2040 ( 
.A(n_2036),
.B(n_23),
.Y(n_2040)
);

NOR3xp33_ASAP7_75t_SL g2041 ( 
.A(n_2004),
.B(n_619),
.C(n_617),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_2012),
.Y(n_2042)
);

OAI31xp33_ASAP7_75t_L g2043 ( 
.A1(n_2034),
.A2(n_2035),
.A3(n_2007),
.B(n_2032),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_2002),
.B(n_627),
.C(n_625),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_L g2045 ( 
.A(n_2038),
.B(n_632),
.C(n_628),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2019),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2024),
.B(n_1881),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_R g2048 ( 
.A(n_2007),
.B(n_24),
.Y(n_2048)
);

NAND4xp25_ASAP7_75t_L g2049 ( 
.A(n_2005),
.B(n_2026),
.C(n_2016),
.D(n_2025),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_2029),
.B(n_1908),
.Y(n_2050)
);

BUFx2_ASAP7_75t_L g2051 ( 
.A(n_2010),
.Y(n_2051)
);

AOI211xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2000),
.A2(n_1826),
.B(n_26),
.C(n_24),
.Y(n_2052)
);

XOR2x1_ASAP7_75t_L g2053 ( 
.A(n_2027),
.B(n_25),
.Y(n_2053)
);

NAND4xp75_ASAP7_75t_L g2054 ( 
.A(n_2001),
.B(n_31),
.C(n_26),
.D(n_28),
.Y(n_2054)
);

NOR3xp33_ASAP7_75t_L g2055 ( 
.A(n_2030),
.B(n_637),
.C(n_634),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_L g2056 ( 
.A(n_2033),
.B(n_2021),
.C(n_2011),
.Y(n_2056)
);

NOR2x1_ASAP7_75t_L g2057 ( 
.A(n_2022),
.B(n_32),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_SL g2058 ( 
.A(n_2013),
.B(n_642),
.C(n_641),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_2008),
.B(n_2037),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2018),
.Y(n_2060)
);

AOI21xp33_ASAP7_75t_L g2061 ( 
.A1(n_2031),
.A2(n_33),
.B(n_36),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2017),
.B(n_36),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2023),
.B(n_37),
.Y(n_2063)
);

NOR3x1_ASAP7_75t_L g2064 ( 
.A(n_2014),
.B(n_38),
.C(n_39),
.Y(n_2064)
);

NOR2xp67_ASAP7_75t_L g2065 ( 
.A(n_2028),
.B(n_40),
.Y(n_2065)
);

OA21x2_ASAP7_75t_L g2066 ( 
.A1(n_2003),
.A2(n_40),
.B(n_44),
.Y(n_2066)
);

NAND5xp2_ASAP7_75t_L g2067 ( 
.A(n_2009),
.B(n_46),
.C(n_48),
.D(n_49),
.E(n_50),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_L g2068 ( 
.A(n_2015),
.B(n_651),
.C(n_648),
.Y(n_2068)
);

AOI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_2006),
.A2(n_1907),
.B1(n_1908),
.B2(n_1878),
.Y(n_2069)
);

CKINVDCx20_ASAP7_75t_R g2070 ( 
.A(n_2010),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2012),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_2010),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_R g2073 ( 
.A(n_2007),
.B(n_49),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2020),
.A2(n_1907),
.B1(n_652),
.B2(n_683),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_SL g2075 ( 
.A(n_2010),
.B(n_655),
.C(n_654),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_2030),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_2019),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2019),
.B(n_50),
.Y(n_2078)
);

BUFx4f_ASAP7_75t_SL g2079 ( 
.A(n_2002),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2012),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2019),
.B(n_51),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2013),
.A2(n_656),
.B1(n_657),
.B2(n_660),
.C(n_663),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2032),
.A2(n_675),
.B(n_666),
.Y(n_2083)
);

NAND4xp25_ASAP7_75t_L g2084 ( 
.A(n_2020),
.B(n_51),
.C(n_53),
.D(n_56),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2019),
.B(n_53),
.Y(n_2085)
);

AOI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_2020),
.A2(n_681),
.B1(n_60),
.B2(n_61),
.C(n_62),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2019),
.B(n_57),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2012),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2020),
.A2(n_1124),
.B1(n_1130),
.B2(n_1134),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_L g2090 ( 
.A(n_2036),
.B(n_61),
.Y(n_2090)
);

AOI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_2020),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.C(n_67),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2012),
.Y(n_2092)
);

NAND3xp33_ASAP7_75t_L g2093 ( 
.A(n_2043),
.B(n_1134),
.C(n_1130),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_SL g2094 ( 
.A(n_2072),
.B(n_63),
.C(n_68),
.Y(n_2094)
);

NAND3xp33_ASAP7_75t_L g2095 ( 
.A(n_2080),
.B(n_1134),
.C(n_1130),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_2042),
.B(n_1137),
.Y(n_2096)
);

XNOR2x1_ASAP7_75t_L g2097 ( 
.A(n_2054),
.B(n_69),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_R g2098 ( 
.A(n_2070),
.B(n_74),
.Y(n_2098)
);

NAND2xp33_ASAP7_75t_SL g2099 ( 
.A(n_2048),
.B(n_1137),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_R g2100 ( 
.A(n_2088),
.B(n_74),
.Y(n_2100)
);

NAND2xp33_ASAP7_75t_SL g2101 ( 
.A(n_2073),
.B(n_2071),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_SL g2102 ( 
.A(n_2092),
.B(n_1137),
.Y(n_2102)
);

NAND2xp33_ASAP7_75t_R g2103 ( 
.A(n_2066),
.B(n_75),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_2079),
.B(n_1221),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2087),
.B(n_75),
.Y(n_2105)
);

NAND2xp33_ASAP7_75t_SL g2106 ( 
.A(n_2078),
.B(n_77),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_R g2107 ( 
.A(n_2075),
.B(n_78),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_2040),
.A2(n_1774),
.B(n_1819),
.Y(n_2108)
);

XNOR2xp5_ASAP7_75t_L g2109 ( 
.A(n_2077),
.B(n_79),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_R g2110 ( 
.A(n_2060),
.B(n_80),
.Y(n_2110)
);

NAND2xp33_ASAP7_75t_SL g2111 ( 
.A(n_2081),
.B(n_82),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2050),
.B(n_82),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_2065),
.B(n_1238),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_2046),
.B(n_1238),
.Y(n_2114)
);

NOR3xp33_ASAP7_75t_SL g2115 ( 
.A(n_2049),
.B(n_83),
.C(n_85),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2050),
.B(n_89),
.Y(n_2116)
);

NAND2xp33_ASAP7_75t_SL g2117 ( 
.A(n_2085),
.B(n_90),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_R g2118 ( 
.A(n_2051),
.B(n_90),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_R g2119 ( 
.A(n_2058),
.B(n_93),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_R g2120 ( 
.A(n_2076),
.B(n_93),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_SL g2121 ( 
.A(n_2041),
.B(n_96),
.Y(n_2121)
);

NOR3xp33_ASAP7_75t_SL g2122 ( 
.A(n_2062),
.B(n_96),
.C(n_99),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_2059),
.B(n_103),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_2090),
.B(n_1238),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2047),
.B(n_2053),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_R g2126 ( 
.A(n_2064),
.B(n_104),
.Y(n_2126)
);

NAND2xp33_ASAP7_75t_SL g2127 ( 
.A(n_2067),
.B(n_2084),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2055),
.B(n_106),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2091),
.B(n_2086),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_R g2130 ( 
.A(n_2061),
.B(n_107),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_R g2131 ( 
.A(n_2057),
.B(n_108),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_R g2132 ( 
.A(n_2063),
.B(n_114),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_2074),
.B(n_1247),
.Y(n_2133)
);

NAND2xp33_ASAP7_75t_SL g2134 ( 
.A(n_2066),
.B(n_2039),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_R g2135 ( 
.A(n_2045),
.B(n_117),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_2044),
.B(n_1247),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2101),
.A2(n_2056),
.B1(n_2068),
.B2(n_2083),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2109),
.Y(n_2138)
);

INVxp67_ASAP7_75t_SL g2139 ( 
.A(n_2103),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2112),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2116),
.Y(n_2141)
);

INVxp67_ASAP7_75t_SL g2142 ( 
.A(n_2097),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2105),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2094),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2115),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2098),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2110),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2118),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2120),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2100),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2125),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2128),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2122),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2127),
.A2(n_2134),
.B1(n_2117),
.B2(n_2111),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2106),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2113),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2124),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2129),
.B(n_2089),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2126),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2093),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2131),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_2132),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2104),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2096),
.Y(n_2164)
);

AND2x4_ASAP7_75t_SL g2165 ( 
.A(n_2123),
.B(n_2069),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2114),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2130),
.Y(n_2167)
);

AO22x2_ASAP7_75t_L g2168 ( 
.A1(n_2095),
.A2(n_2136),
.B1(n_2133),
.B2(n_2099),
.Y(n_2168)
);

NOR2x1_ASAP7_75t_L g2169 ( 
.A(n_2102),
.B(n_2082),
.Y(n_2169)
);

NOR3xp33_ASAP7_75t_SL g2170 ( 
.A(n_2121),
.B(n_2052),
.C(n_120),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2107),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2108),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2135),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2139),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_2145),
.B(n_2119),
.Y(n_2175)
);

AOI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2151),
.A2(n_1261),
.B1(n_1255),
.B2(n_1247),
.Y(n_2176)
);

BUFx2_ASAP7_75t_L g2177 ( 
.A(n_2170),
.Y(n_2177)
);

AOI22x1_ASAP7_75t_L g2178 ( 
.A1(n_2142),
.A2(n_1261),
.B1(n_1255),
.B2(n_1037),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2165),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2144),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2148),
.Y(n_2181)
);

INVxp67_ASAP7_75t_L g2182 ( 
.A(n_2147),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2143),
.Y(n_2183)
);

XNOR2xp5_ASAP7_75t_L g2184 ( 
.A(n_2154),
.B(n_121),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2146),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2149),
.Y(n_2186)
);

NAND2xp33_ASAP7_75t_SL g2187 ( 
.A(n_2153),
.B(n_1255),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2162),
.Y(n_2188)
);

AO22x2_ASAP7_75t_L g2189 ( 
.A1(n_2150),
.A2(n_1078),
.B1(n_1068),
.B2(n_1047),
.Y(n_2189)
);

AOI22x1_ASAP7_75t_L g2190 ( 
.A1(n_2168),
.A2(n_1261),
.B1(n_1037),
.B2(n_1078),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2155),
.Y(n_2191)
);

AOI22x1_ASAP7_75t_L g2192 ( 
.A1(n_2168),
.A2(n_2159),
.B1(n_2138),
.B2(n_2167),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2140),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2141),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2161),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2171),
.Y(n_2196)
);

XOR2xp5_ASAP7_75t_L g2197 ( 
.A(n_2152),
.B(n_2173),
.Y(n_2197)
);

XNOR2x1_ASAP7_75t_L g2198 ( 
.A(n_2158),
.B(n_122),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2172),
.Y(n_2199)
);

XNOR2xp5_ASAP7_75t_L g2200 ( 
.A(n_2137),
.B(n_124),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2156),
.A2(n_1837),
.B1(n_1836),
.B2(n_1047),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2158),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2169),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2163),
.Y(n_2204)
);

OA22x2_ASAP7_75t_L g2205 ( 
.A1(n_2157),
.A2(n_1068),
.B1(n_1812),
.B2(n_128),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2164),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2200),
.Y(n_2207)
);

AO22x1_ASAP7_75t_L g2208 ( 
.A1(n_2202),
.A2(n_2160),
.B1(n_2166),
.B2(n_1082),
.Y(n_2208)
);

AOI221xp5_ASAP7_75t_SL g2209 ( 
.A1(n_2182),
.A2(n_1082),
.B1(n_1063),
.B2(n_1059),
.C(n_1056),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2198),
.Y(n_2210)
);

BUFx2_ASAP7_75t_SL g2211 ( 
.A(n_2183),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2205),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2184),
.B(n_126),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2174),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2179),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2191),
.A2(n_1082),
.B1(n_1063),
.B2(n_1059),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2206),
.Y(n_2217)
);

OAI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2204),
.A2(n_127),
.B(n_131),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2199),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2192),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2193),
.B(n_1753),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2188),
.Y(n_2222)
);

XNOR2x1_ASAP7_75t_L g2223 ( 
.A(n_2197),
.B(n_137),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2185),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2194),
.Y(n_2225)
);

OAI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_2215),
.A2(n_2203),
.B1(n_2181),
.B2(n_2186),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2223),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_2220),
.B(n_2180),
.Y(n_2228)
);

OAI22x1_ASAP7_75t_L g2229 ( 
.A1(n_2217),
.A2(n_2196),
.B1(n_2177),
.B2(n_2175),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2211),
.Y(n_2230)
);

AO211x2_ASAP7_75t_L g2231 ( 
.A1(n_2219),
.A2(n_2195),
.B(n_2189),
.C(n_2187),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2213),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2222),
.A2(n_2189),
.B(n_2190),
.Y(n_2233)
);

HB1xp67_ASAP7_75t_L g2234 ( 
.A(n_2224),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2214),
.A2(n_2176),
.B1(n_2201),
.B2(n_2178),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_2234),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_2226),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2230),
.A2(n_2225),
.B1(n_2207),
.B2(n_2212),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2229),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2227),
.B(n_2221),
.Y(n_2240)
);

CKINVDCx20_ASAP7_75t_R g2241 ( 
.A(n_2228),
.Y(n_2241)
);

OR2x6_ASAP7_75t_L g2242 ( 
.A(n_2232),
.B(n_2210),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2236),
.B(n_2237),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2238),
.A2(n_2233),
.B(n_2235),
.Y(n_2244)
);

AOI21xp33_ASAP7_75t_SL g2245 ( 
.A1(n_2239),
.A2(n_2208),
.B(n_2216),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2241),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2246),
.B(n_2243),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2244),
.A2(n_2242),
.B1(n_2240),
.B2(n_2218),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2245),
.A2(n_2242),
.B1(n_2231),
.B2(n_2209),
.Y(n_2249)
);

XOR2xp5_ASAP7_75t_L g2250 ( 
.A(n_2246),
.B(n_139),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2247),
.B(n_140),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2248),
.B(n_141),
.Y(n_2252)
);

NAND3xp33_ASAP7_75t_L g2253 ( 
.A(n_2249),
.B(n_1063),
.C(n_1059),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2253),
.A2(n_2250),
.B1(n_1056),
.B2(n_1023),
.Y(n_2254)
);

OAI221xp5_ASAP7_75t_L g2255 ( 
.A1(n_2252),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.C(n_146),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2254),
.A2(n_2251),
.B1(n_986),
.B2(n_1022),
.Y(n_2256)
);

AOI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_2255),
.A2(n_986),
.B1(n_1022),
.B2(n_153),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2257),
.B(n_147),
.Y(n_2258)
);

AOI221xp5_ASAP7_75t_L g2259 ( 
.A1(n_2256),
.A2(n_986),
.B1(n_155),
.B2(n_157),
.C(n_158),
.Y(n_2259)
);

AOI221xp5_ASAP7_75t_L g2260 ( 
.A1(n_2259),
.A2(n_151),
.B1(n_159),
.B2(n_163),
.C(n_165),
.Y(n_2260)
);

AOI211xp5_ASAP7_75t_L g2261 ( 
.A1(n_2260),
.A2(n_2258),
.B(n_168),
.C(n_175),
.Y(n_2261)
);


endmodule