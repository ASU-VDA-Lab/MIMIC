module real_aes_12416_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_47;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_0), .B(n_6), .C(n_22), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_1), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g38 ( .A(n_1), .B(n_39), .Y(n_38) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_2), .B(n_13), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_2), .B(n_30), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g45 ( .A(n_2), .Y(n_45) );
NAND2xp33_ASAP7_75t_R g47 ( .A(n_2), .B(n_13), .Y(n_47) );
NAND5xp2_ASAP7_75t_SL g18 ( .A(n_3), .B(n_5), .C(n_19), .D(n_24), .E(n_25), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_3), .Y(n_40) );
AOI322xp5_ASAP7_75t_R g32 ( .A1(n_4), .A2(n_8), .A3(n_26), .B1(n_33), .B2(n_38), .C1(n_42), .C2(n_46), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_5), .B(n_20), .Y(n_41) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_7), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_9), .Y(n_25) );
NAND3xp33_ASAP7_75t_SL g39 ( .A(n_9), .B(n_40), .C(n_41), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_10), .Y(n_31) );
INVx3_ASAP7_75t_L g37 ( .A(n_11), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_12), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_13), .Y(n_30) );
NOR2xp33_ASAP7_75t_R g44 ( .A(n_13), .B(n_45), .Y(n_44) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_14), .Y(n_22) );
OAI221xp5_ASAP7_75t_R g15 ( .A1(n_16), .A2(n_27), .B1(n_28), .B2(n_31), .C(n_32), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_17), .B(n_26), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g28 ( .A(n_17), .B(n_29), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_18), .B(n_43), .Y(n_42) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_18), .B(n_47), .Y(n_46) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g20 ( .A(n_21), .B(n_23), .Y(n_20) );
INVx1_ASAP7_75t_L g33 ( .A(n_34), .Y(n_33) );
BUFx3_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_37), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g43 ( .A(n_44), .Y(n_43) );
endmodule