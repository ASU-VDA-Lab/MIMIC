module fake_jpeg_26777_n_107 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_11),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_1),
.B(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_22),
.B(n_21),
.C(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_42),
.B1(n_15),
.B2(n_23),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_15),
.B1(n_11),
.B2(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_56),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_26),
.B1(n_32),
.B2(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_16),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_18),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_20),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_36),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_62),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_43),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_38),
.C(n_17),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_47),
.Y(n_72)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_80),
.B1(n_60),
.B2(n_70),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_58),
.B(n_46),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_50),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_61),
.C(n_66),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_35),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_71),
.C(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_74),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_62),
.C(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_7),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_86),
.C(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_68),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_57),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_35),
.B(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_90),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_9),
.B(n_6),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_5),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_97),
.Y(n_104)
);

OAI31xp33_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_2),
.A3(n_3),
.B(n_14),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_14),
.A3(n_27),
.B1(n_63),
.B2(n_101),
.C1(n_73),
.C2(n_93),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_105),
.C(n_102),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_63),
.Y(n_107)
);


endmodule