module real_aes_8422_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_1), .A2(n_146), .B(n_151), .C(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g258 ( .A(n_2), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_3), .A2(n_141), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_4), .B(n_218), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_5), .Y(n_124) );
AOI21xp33_ASAP7_75t_L g219 ( .A1(n_6), .A2(n_141), .B(n_220), .Y(n_219) );
AND2x6_ASAP7_75t_L g146 ( .A(n_7), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_8), .A2(n_140), .B(n_148), .Y(n_139) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_9), .B(n_40), .Y(n_123) );
INVx1_ASAP7_75t_L g553 ( .A(n_10), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_11), .B(n_190), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_12), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g225 ( .A(n_13), .Y(n_225) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
INVx1_ASAP7_75t_L g158 ( .A(n_15), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_16), .A2(n_159), .B(n_173), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_17), .B(n_218), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_18), .B(n_175), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_19), .B(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_20), .B(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_21), .A2(n_206), .B(n_232), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_22), .B(n_218), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_23), .B(n_190), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_24), .A2(n_155), .B(n_157), .C(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_25), .B(n_190), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_26), .Y(n_481) );
INVx1_ASAP7_75t_L g449 ( .A(n_27), .Y(n_449) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_28), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_29), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_30), .B(n_190), .Y(n_259) );
INVx1_ASAP7_75t_L g474 ( .A(n_31), .Y(n_474) );
INVx1_ASAP7_75t_L g237 ( .A(n_32), .Y(n_237) );
INVx2_ASAP7_75t_L g144 ( .A(n_33), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_34), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_35), .A2(n_206), .B(n_226), .C(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_L g475 ( .A(n_36), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_37), .A2(n_146), .B(n_151), .C(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_38), .A2(n_151), .B(n_448), .C(n_453), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g460 ( .A(n_39), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_40), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g235 ( .A(n_41), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_42), .A2(n_177), .B(n_223), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_43), .B(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_44), .A2(n_437), .B1(n_706), .B2(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_44), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_45), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_46), .Y(n_471) );
INVx1_ASAP7_75t_L g519 ( .A(n_47), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_48), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_49), .B(n_141), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_50), .A2(n_151), .B1(n_232), .B2(n_234), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_51), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_52), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_53), .A2(n_100), .B1(n_111), .B2(n_718), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_54), .A2(n_223), .B(n_224), .C(n_226), .Y(n_222) );
CKINVDCx14_ASAP7_75t_R g550 ( .A(n_55), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_56), .Y(n_194) );
INVx1_ASAP7_75t_L g221 ( .A(n_57), .Y(n_221) );
INVx1_ASAP7_75t_L g147 ( .A(n_58), .Y(n_147) );
INVx1_ASAP7_75t_L g137 ( .A(n_59), .Y(n_137) );
INVx1_ASAP7_75t_SL g463 ( .A(n_60), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_62), .B(n_218), .Y(n_523) );
INVx1_ASAP7_75t_L g484 ( .A(n_63), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_64), .A2(n_175), .B(n_226), .C(n_246), .Y(n_245) );
INVxp67_ASAP7_75t_L g247 ( .A(n_65), .Y(n_247) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_66), .A2(n_68), .B1(n_126), .B2(n_701), .C1(n_702), .C2(n_709), .Y(n_125) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
INVx1_ASAP7_75t_L g701 ( .A(n_68), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_69), .A2(n_141), .B(n_549), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_70), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_71), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_72), .A2(n_141), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g185 ( .A(n_73), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_74), .A2(n_140), .B(n_470), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_75), .Y(n_446) );
INVx1_ASAP7_75t_L g511 ( .A(n_76), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_77), .A2(n_146), .B(n_151), .C(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_78), .A2(n_141), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g514 ( .A(n_79), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_80), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx1_ASAP7_75t_L g503 ( .A(n_82), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_83), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_84), .A2(n_146), .B(n_151), .C(n_257), .Y(n_256) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_85), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g120 ( .A(n_85), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g436 ( .A(n_85), .Y(n_436) );
OR2x2_ASAP7_75t_L g700 ( .A(n_85), .B(n_122), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_86), .A2(n_151), .B(n_483), .C(n_487), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_87), .B(n_134), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_88), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_89), .A2(n_146), .B(n_151), .C(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_90), .Y(n_211) );
INVx1_ASAP7_75t_L g244 ( .A(n_91), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_92), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_93), .B(n_172), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_94), .B(n_163), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_95), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_97), .A2(n_141), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g522 ( .A(n_98), .Y(n_522) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx5_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g718 ( .A(n_103), .Y(n_718) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g122 ( .A(n_107), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AOI22x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_125), .B1(n_712), .B2(n_713), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_117), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g712 ( .A(n_115), .Y(n_712) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_117), .A2(n_714), .B(n_716), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_124), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g717 ( .A(n_120), .Y(n_717) );
NOR2x2_ASAP7_75t_L g711 ( .A(n_121), .B(n_436), .Y(n_711) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g435 ( .A(n_122), .B(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_435), .B1(n_437), .B2(n_700), .Y(n_126) );
INVx2_ASAP7_75t_SL g703 ( .A(n_127), .Y(n_703) );
OR4x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_331), .C(n_390), .D(n_417), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_273), .C(n_298), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_196), .B(n_216), .C(n_249), .Y(n_129) );
AOI211xp5_ASAP7_75t_SL g421 ( .A1(n_130), .A2(n_422), .B(n_424), .C(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
INVx1_ASAP7_75t_L g296 ( .A(n_131), .Y(n_296) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g271 ( .A(n_132), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g303 ( .A(n_132), .Y(n_303) );
AND2x2_ASAP7_75t_L g358 ( .A(n_132), .B(n_327), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_132), .B(n_214), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_132), .B(n_215), .Y(n_416) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g277 ( .A(n_133), .Y(n_277) );
AND2x2_ASAP7_75t_L g320 ( .A(n_133), .B(n_183), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_133), .B(n_215), .Y(n_338) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B(n_162), .Y(n_133) );
INVx1_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
INVx2_ASAP7_75t_L g200 ( .A(n_134), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_134), .A2(n_186), .B(n_446), .C(n_447), .Y(n_445) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_134), .A2(n_548), .B(n_554), .Y(n_547) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_L g164 ( .A(n_135), .B(n_136), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_142), .B(n_146), .Y(n_186) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g452 ( .A(n_143), .Y(n_452) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g233 ( .A(n_144), .Y(n_233) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx3_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
INVx4_ASAP7_75t_SL g161 ( .A(n_146), .Y(n_161) );
BUFx3_ASAP7_75t_L g453 ( .A(n_146), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_161), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_150), .A2(n_161), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_150), .A2(n_161), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_150), .A2(n_161), .B(n_460), .C(n_461), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_SL g470 ( .A1(n_150), .A2(n_161), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_150), .A2(n_161), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_150), .A2(n_161), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_150), .A2(n_161), .B(n_550), .C(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_155), .B(n_158), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_155), .A2(n_172), .B1(n_474), .B2(n_475), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_155), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_155), .B(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_156), .A2(n_235), .B1(n_236), .B2(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g236 ( .A(n_156), .Y(n_236) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g230 ( .A1(n_161), .A2(n_186), .B1(n_231), .B2(n_238), .Y(n_230) );
INVx1_ASAP7_75t_L g487 ( .A(n_161), .Y(n_487) );
INVx4_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_163), .A2(n_242), .B(n_248), .Y(n_241) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_163), .Y(n_457) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx4_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_165), .A2(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g406 ( .A(n_165), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_183), .Y(n_165) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
AND2x2_ASAP7_75t_L g275 ( .A(n_166), .B(n_215), .Y(n_275) );
OR2x2_ASAP7_75t_L g304 ( .A(n_166), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g318 ( .A(n_166), .Y(n_318) );
INVx3_ASAP7_75t_L g327 ( .A(n_166), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_166), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g370 ( .A(n_166), .B(n_276), .Y(n_370) );
AND2x2_ASAP7_75t_L g394 ( .A(n_166), .B(n_350), .Y(n_394) );
OR2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_180), .Y(n_166) );
AOI21xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_178), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_176), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_172), .A2(n_258), .B(n_259), .C(n_260), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_172), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_173), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_173), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_173), .B(n_553), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_176), .A2(n_189), .B(n_191), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_176), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
O2A1O1Ixp5_ASAP7_75t_L g502 ( .A1(n_176), .A2(n_485), .B(n_503), .C(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g192 ( .A(n_178), .Y(n_192) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_230), .B(n_239), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_179), .B(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_179), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx3_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_182), .B(n_455), .Y(n_454) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_182), .A2(n_480), .B(n_488), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_182), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
AND2x2_ASAP7_75t_L g430 ( .A(n_183), .B(n_272), .Y(n_430) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_192), .B(n_193), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_255), .B(n_256), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_186), .A2(n_481), .B(n_482), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_186), .A2(n_500), .B(n_501), .Y(n_499) );
INVx4_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
INVx2_ASAP7_75t_L g223 ( .A(n_190), .Y(n_223) );
INVx1_ASAP7_75t_L g468 ( .A(n_192), .Y(n_468) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_192), .A2(n_493), .B(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_195), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_195), .B(n_262), .Y(n_261) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_195), .A2(n_499), .B(n_505), .Y(n_498) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_212), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_198), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g350 ( .A(n_198), .B(n_338), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_198), .B(n_327), .Y(n_412) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
AND2x2_ASAP7_75t_L g276 ( .A(n_199), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g317 ( .A(n_199), .B(n_318), .Y(n_317) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
INVx1_ASAP7_75t_L g477 ( .A(n_200), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_200), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_209), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_206), .B(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g226 ( .A(n_208), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_212), .B(n_313), .Y(n_335) );
INVx1_ASAP7_75t_L g374 ( .A(n_212), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_212), .B(n_301), .Y(n_418) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g281 ( .A(n_213), .B(n_276), .Y(n_281) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_215), .B(n_272), .Y(n_305) );
INVx1_ASAP7_75t_L g384 ( .A(n_215), .Y(n_384) );
AOI322xp5_ASAP7_75t_L g408 ( .A1(n_216), .A2(n_323), .A3(n_383), .B1(n_409), .B2(n_411), .C1(n_413), .C2(n_415), .Y(n_408) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_217), .B(n_228), .Y(n_216) );
AND2x2_ASAP7_75t_L g263 ( .A(n_217), .B(n_241), .Y(n_263) );
INVx1_ASAP7_75t_SL g266 ( .A(n_217), .Y(n_266) );
AND2x2_ASAP7_75t_L g268 ( .A(n_217), .B(n_229), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_217), .B(n_285), .Y(n_291) );
INVx2_ASAP7_75t_L g310 ( .A(n_217), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_217), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g361 ( .A(n_217), .B(n_285), .Y(n_361) );
BUFx2_ASAP7_75t_L g378 ( .A(n_217), .Y(n_378) );
AND2x2_ASAP7_75t_L g392 ( .A(n_217), .B(n_252), .Y(n_392) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_228), .B(n_280), .Y(n_307) );
AND2x2_ASAP7_75t_L g434 ( .A(n_228), .B(n_310), .Y(n_434) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_241), .Y(n_228) );
OR2x2_ASAP7_75t_L g279 ( .A(n_229), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g285 ( .A(n_229), .Y(n_285) );
AND2x2_ASAP7_75t_L g330 ( .A(n_229), .B(n_253), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_229), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_229), .Y(n_414) );
INVx2_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g485 ( .A(n_236), .Y(n_485) );
AND2x2_ASAP7_75t_L g265 ( .A(n_241), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
BUFx2_ASAP7_75t_L g293 ( .A(n_241), .Y(n_293) );
AND2x2_ASAP7_75t_L g312 ( .A(n_241), .B(n_285), .Y(n_312) );
INVx3_ASAP7_75t_L g324 ( .A(n_241), .Y(n_324) );
OR2x2_ASAP7_75t_L g334 ( .A(n_241), .B(n_285), .Y(n_334) );
AOI31xp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_264), .A3(n_267), .B(n_269), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_263), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_251), .B(n_286), .Y(n_297) );
OR2x2_ASAP7_75t_L g321 ( .A(n_251), .B(n_291), .Y(n_321) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_252), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_334), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_252), .B(n_324), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_252), .B(n_360), .Y(n_359) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_252), .B(n_323), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_252), .B(n_378), .Y(n_388) );
AND2x2_ASAP7_75t_L g400 ( .A(n_252), .B(n_285), .Y(n_400) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g280 ( .A(n_253), .Y(n_280) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_263), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_265), .B(n_341), .Y(n_375) );
AND2x4_ASAP7_75t_L g286 ( .A(n_266), .B(n_287), .Y(n_286) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g365 ( .A(n_271), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_271), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g313 ( .A(n_272), .B(n_303), .Y(n_313) );
AND2x2_ASAP7_75t_L g407 ( .A(n_272), .B(n_277), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_272), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B1(n_281), .B2(n_282), .C(n_288), .Y(n_273) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_274), .Y(n_294) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_275), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_278), .B(n_329), .Y(n_348) );
INVx3_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g397 ( .A(n_279), .B(n_293), .Y(n_397) );
AND2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g341 ( .A(n_280), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_280), .B(n_324), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_280), .B(n_381), .C(n_412), .Y(n_411) );
AOI211xp5_ASAP7_75t_SL g344 ( .A1(n_281), .A2(n_345), .B(n_347), .C(n_355), .Y(n_344) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_283), .A2(n_334), .B1(n_335), .B2(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_284), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_284), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g426 ( .A(n_286), .B(n_400), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .B1(n_295), .B2(n_297), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_292), .B(n_341), .Y(n_372) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_295), .A2(n_387), .B1(n_418), .B2(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_306), .B1(n_308), .B2(n_313), .C(n_314), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_304), .A2(n_315), .B1(n_321), .B2(n_322), .C(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g357 ( .A(n_305), .Y(n_357) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g329 ( .A(n_310), .Y(n_329) );
OR2x2_ASAP7_75t_L g402 ( .A(n_310), .B(n_334), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_310), .B(n_312), .Y(n_404) );
INVx1_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_316), .A2(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g380 ( .A(n_316), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g354 ( .A(n_317), .B(n_338), .Y(n_354) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp33_ASAP7_75t_SL g371 ( .A(n_322), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_323), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_324), .B(n_360), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_327), .A2(n_340), .B(n_342), .C(n_343), .Y(n_339) );
NAND2x1_ASAP7_75t_SL g364 ( .A(n_327), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_328), .A2(n_377), .B1(n_379), .B2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_330), .B(n_420), .Y(n_419) );
NAND5xp2_ASAP7_75t_L g331 ( .A(n_332), .B(n_344), .C(n_362), .D(n_376), .E(n_385), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_339), .Y(n_332) );
INVx1_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_337), .A2(n_356), .B1(n_396), .B2(n_398), .C(n_401), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_338), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_341), .B(n_407), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_351), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g429 ( .A(n_358), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_370), .B2(n_371), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g413 ( .A(n_368), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g420 ( .A(n_378), .Y(n_420) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_393), .B(n_395), .C(n_408), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_418), .B(n_419), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_397), .B(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B(n_433), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g705 ( .A(n_435), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_437), .Y(n_706) );
OR3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_611), .C(n_658), .Y(n_437) );
NAND3xp33_ASAP7_75t_SL g438 ( .A(n_439), .B(n_557), .C(n_582), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_497), .B1(n_524), .B2(n_527), .C(n_535), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_465), .B(n_490), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_442), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_442), .B(n_540), .Y(n_655) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_456), .Y(n_442) );
AND2x2_ASAP7_75t_L g526 ( .A(n_443), .B(n_496), .Y(n_526) );
AND2x2_ASAP7_75t_L g575 ( .A(n_443), .B(n_495), .Y(n_575) );
AND2x2_ASAP7_75t_L g596 ( .A(n_443), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g601 ( .A(n_443), .B(n_568), .Y(n_601) );
OR2x2_ASAP7_75t_L g609 ( .A(n_443), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g681 ( .A(n_443), .B(n_478), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_443), .B(n_630), .Y(n_695) );
INVx3_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g541 ( .A(n_444), .B(n_456), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_444), .B(n_478), .Y(n_542) );
AND2x4_ASAP7_75t_L g563 ( .A(n_444), .B(n_496), .Y(n_563) );
AND2x2_ASAP7_75t_L g593 ( .A(n_444), .B(n_467), .Y(n_593) );
AND2x2_ASAP7_75t_L g602 ( .A(n_444), .B(n_592), .Y(n_602) );
AND2x2_ASAP7_75t_L g618 ( .A(n_444), .B(n_479), .Y(n_618) );
OR2x2_ASAP7_75t_L g627 ( .A(n_444), .B(n_610), .Y(n_627) );
AND2x2_ASAP7_75t_L g633 ( .A(n_444), .B(n_568), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_444), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g647 ( .A(n_444), .B(n_492), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_444), .B(n_537), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_444), .B(n_597), .Y(n_686) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_452), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g496 ( .A(n_456), .Y(n_496) );
AND2x2_ASAP7_75t_L g592 ( .A(n_456), .B(n_478), .Y(n_592) );
AND2x2_ASAP7_75t_L g597 ( .A(n_456), .B(n_479), .Y(n_597) );
INVx1_ASAP7_75t_L g653 ( .A(n_456), .Y(n_653) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_464), .Y(n_456) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_457), .A2(n_509), .B(n_515), .Y(n_508) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_457), .A2(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g562 ( .A(n_466), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_478), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_467), .B(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
OR2x2_ASAP7_75t_L g610 ( .A(n_467), .B(n_478), .Y(n_610) );
OR2x2_ASAP7_75t_L g671 ( .A(n_467), .B(n_578), .Y(n_671) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_476), .Y(n_467) );
INVx1_ASAP7_75t_L g493 ( .A(n_469), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_476), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_478), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g630 ( .A(n_478), .B(n_492), .Y(n_630) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_491), .A2(n_675), .B1(n_679), .B2(n_682), .C(n_683), .Y(n_674) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .Y(n_491) );
INVx1_ASAP7_75t_SL g538 ( .A(n_492), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_492), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g669 ( .A(n_492), .B(n_526), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_495), .B(n_540), .Y(n_661) );
AND2x2_ASAP7_75t_L g568 ( .A(n_496), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g572 ( .A(n_497), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_497), .B(n_578), .Y(n_608) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
AND2x2_ASAP7_75t_L g534 ( .A(n_498), .B(n_508), .Y(n_534) );
INVx4_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
BUFx3_ASAP7_75t_L g588 ( .A(n_498), .Y(n_588) );
AND3x2_ASAP7_75t_L g603 ( .A(n_498), .B(n_604), .C(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g685 ( .A(n_507), .B(n_599), .Y(n_685) );
AND2x2_ASAP7_75t_L g693 ( .A(n_507), .B(n_578), .Y(n_693) );
INVx1_ASAP7_75t_SL g698 ( .A(n_507), .Y(n_698) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
INVx1_ASAP7_75t_SL g556 ( .A(n_508), .Y(n_556) );
AND2x2_ASAP7_75t_L g579 ( .A(n_508), .B(n_546), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_508), .B(n_530), .Y(n_581) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_508), .Y(n_621) );
OR2x2_ASAP7_75t_L g626 ( .A(n_508), .B(n_546), .Y(n_626) );
INVx2_ASAP7_75t_L g532 ( .A(n_516), .Y(n_532) );
AND2x2_ASAP7_75t_L g566 ( .A(n_516), .B(n_547), .Y(n_566) );
OR2x2_ASAP7_75t_L g586 ( .A(n_516), .B(n_547), .Y(n_586) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_516), .Y(n_606) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
AOI21xp33_ASAP7_75t_L g656 ( .A1(n_525), .A2(n_565), .B(n_657), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_527), .A2(n_537), .A3(n_563), .B1(n_693), .B2(n_694), .C1(n_696), .C2(n_699), .Y(n_692) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_529), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_530), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g555 ( .A(n_531), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_546), .Y(n_623) );
AND2x2_ASAP7_75t_L g690 ( .A(n_532), .B(n_547), .Y(n_690) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g631 ( .A(n_534), .B(n_585), .Y(n_631) );
AOI31xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_539), .A3(n_542), .B(n_543), .Y(n_535) );
AND2x2_ASAP7_75t_L g590 ( .A(n_537), .B(n_568), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_537), .B(n_560), .Y(n_672) );
AND2x2_ASAP7_75t_L g691 ( .A(n_537), .B(n_596), .Y(n_691) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_540), .B(n_568), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g614 ( .A(n_540), .B(n_597), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_540), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_540), .B(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_541), .B(n_597), .Y(n_629) );
INVx1_ASAP7_75t_L g673 ( .A(n_541), .Y(n_673) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_555), .Y(n_544) );
INVxp67_ASAP7_75t_L g625 ( .A(n_545), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_546), .B(n_556), .Y(n_561) );
INVx1_ASAP7_75t_L g667 ( .A(n_546), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_546), .B(n_644), .Y(n_678) );
BUFx3_ASAP7_75t_L g578 ( .A(n_547), .Y(n_578) );
AND2x2_ASAP7_75t_L g604 ( .A(n_547), .B(n_556), .Y(n_604) );
INVx2_ASAP7_75t_L g644 ( .A(n_547), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_555), .B(n_677), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_562), .B(n_564), .C(n_573), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_559), .A2(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_560), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_560), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g640 ( .A(n_561), .B(n_586), .Y(n_640) );
INVx3_ASAP7_75t_L g571 ( .A(n_563), .Y(n_571) );
OAI22xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_567), .B1(n_570), .B2(n_572), .Y(n_564) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_566), .A2(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g615 ( .A(n_566), .B(n_579), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_566), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g570 ( .A(n_569), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g639 ( .A(n_569), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_570), .A2(n_584), .B(n_589), .Y(n_583) );
OAI22xp33_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_576), .B1(n_580), .B2(n_581), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_575), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g599 ( .A(n_578), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_578), .B(n_621), .Y(n_620) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_594), .C(n_607), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g649 ( .A1(n_584), .A2(n_650), .B1(n_654), .B2(n_655), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g654 ( .A(n_586), .B(n_587), .Y(n_654) );
AND2x2_ASAP7_75t_L g662 ( .A(n_587), .B(n_643), .Y(n_662) );
CKINVDCx16_ASAP7_75t_R g587 ( .A(n_588), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_SL g670 ( .A1(n_588), .A2(n_671), .B(n_672), .C(n_673), .Y(n_670) );
OR2x2_ASAP7_75t_L g697 ( .A(n_588), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_598), .B(n_600), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_596), .A2(n_633), .B(n_634), .C(n_637), .Y(n_632) );
OAI21xp33_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_602), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g665 ( .A(n_604), .B(n_623), .Y(n_665) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g643 ( .A(n_606), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g648 ( .A(n_608), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_632), .C(n_645), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_616), .C(n_624), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g682 ( .A(n_619), .Y(n_682) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g642 ( .A(n_621), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_621), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_627), .C(n_628), .Y(n_624) );
INVx2_ASAP7_75t_SL g636 ( .A(n_626), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_627), .A2(n_638), .B1(n_640), .B2(n_641), .Y(n_637) );
OAI21xp33_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_630), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B(n_649), .C(n_656), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVxp33_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g699 ( .A(n_653), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_674), .C(n_687), .D(n_692), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B(n_663), .C(n_670), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_668), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_664), .A2(n_684), .B(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_671), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g708 ( .A(n_700), .Y(n_708) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_704), .B1(n_706), .B2(n_707), .Y(n_702) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx3_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
endmodule