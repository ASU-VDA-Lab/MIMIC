module fake_netlist_5_1627_n_2962 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_2962);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2962;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_2771;
wire n_785;
wire n_549;
wire n_2617;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_556;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_659;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_579;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2959;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_436;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_475;
wire n_1070;
wire n_422;
wire n_1547;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1587;
wire n_1473;
wire n_680;
wire n_2682;
wire n_901;
wire n_553;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_2932;
wire n_2753;
wire n_464;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_477;
wire n_1585;
wire n_571;
wire n_461;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_1276;
wire n_702;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_1711;
wire n_599;
wire n_1891;
wire n_1662;
wire n_931;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_456;
wire n_959;
wire n_2459;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_457;
wire n_514;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_486;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_512;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2628;
wire n_2390;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_513;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_495;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_2953;
wire n_824;
wire n_1645;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_515;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_2475;
wire n_2733;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2533;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_398;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2282;
wire n_2002;
wire n_510;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_458;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_899;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_487;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_665;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_410;
wire n_2547;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_500;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_435;
wire n_2003;
wire n_1457;
wire n_766;
wire n_541;
wire n_2692;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2430;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_980;
wire n_1115;
wire n_698;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2284;
wire n_2187;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_2850;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_559;
wire n_825;
wire n_2819;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_2104;
wire n_2748;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_428;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_2957;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_2961;
wire n_413;
wire n_402;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_2940;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_2612;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_465;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_453;
wire n_403;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_412;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_2938;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_438;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g398 ( 
.A(n_40),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_87),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_85),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_98),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_52),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_155),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_155),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_97),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_157),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_154),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_212),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_333),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_80),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_200),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_8),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_19),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_214),
.Y(n_416)
);

INVxp33_ASAP7_75t_R g417 ( 
.A(n_6),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_180),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_104),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_296),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_170),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_260),
.Y(n_424)
);

BUFx2_ASAP7_75t_SL g425 ( 
.A(n_256),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_195),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_80),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_223),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_291),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_96),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_190),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_252),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_221),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_149),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_24),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_335),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_49),
.Y(n_437)
);

BUFx10_ASAP7_75t_L g438 ( 
.A(n_68),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_355),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_52),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_177),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_84),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_253),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_284),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_339),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_379),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_157),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_322),
.Y(n_448)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_64),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_391),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_77),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_24),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_189),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_108),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_249),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_345),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_313),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_174),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_241),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_109),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_47),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_139),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_21),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_385),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_377),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_264),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_277),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_162),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_280),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_344),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_83),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_394),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_294),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_47),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_169),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_281),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_12),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_39),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_82),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_378),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_321),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_102),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_149),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_367),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_210),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_60),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_195),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_92),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_338),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_246),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_220),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_183),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_205),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_224),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_51),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_334),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_167),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_208),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_44),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_389),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_134),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_370),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_167),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_371),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_134),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_369),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_125),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_109),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_199),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_50),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_272),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_327),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_324),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_245),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_273),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_59),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_82),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_91),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_61),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_171),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_54),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_196),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_119),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_165),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_206),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_343),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_10),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_384),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_178),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_74),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_262),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_84),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_143),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_85),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_320),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_98),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_328),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_96),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_395),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_316),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_4),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_43),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_5),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_307),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_125),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_75),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_363),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_337),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_143),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_78),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_68),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_210),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_347),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_44),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_141),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_10),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_28),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_269),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_312),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_16),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_164),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_268),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_188),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_380),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_61),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_200),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_89),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_382),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_53),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_213),
.Y(n_572)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_115),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_124),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_21),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_193),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_168),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_330),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_43),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_297),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_74),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_95),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_311),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_350),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_72),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_340),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_7),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_59),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_141),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_32),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_212),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_119),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_376),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_136),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_196),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_144),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_202),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_218),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_26),
.Y(n_599)
);

BUFx5_ASAP7_75t_L g600 ( 
.A(n_323),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_5),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_336),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_26),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_201),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_83),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_342),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_17),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_25),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_130),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_183),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_86),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_3),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_90),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_70),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_257),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_140),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_354),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_108),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_100),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_282),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_275),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_242),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_397),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_158),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_53),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_6),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_76),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_112),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_178),
.Y(n_629)
);

BUFx5_ASAP7_75t_L g630 ( 
.A(n_77),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_194),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_276),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_181),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_319),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_288),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_154),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_247),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_189),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_232),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_270),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_148),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_261),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_331),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_40),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_374),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_255),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_392),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_234),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_352),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_32),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_71),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_308),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_396),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_51),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_286),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_87),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_299),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_164),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_54),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_254),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_13),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_346),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_171),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_27),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_219),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_123),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_139),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_362),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_193),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_318),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_153),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_126),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_45),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_15),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_88),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_56),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_197),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_19),
.Y(n_678)
);

CKINVDCx14_ASAP7_75t_R g679 ( 
.A(n_393),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_227),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_165),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_390),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_15),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_172),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_63),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_208),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_274),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_387),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_176),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_386),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_263),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_368),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_206),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_38),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_215),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_300),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_381),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_226),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_22),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_180),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_388),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_188),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_170),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_293),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_630),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_472),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_630),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_630),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_630),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_630),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_630),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_424),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_400),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_630),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_457),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g716 ( 
.A(n_495),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_630),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_482),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_694),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_543),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_694),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_405),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_573),
.Y(n_723)
);

CKINVDCx16_ASAP7_75t_R g724 ( 
.A(n_534),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_694),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_694),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_694),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_543),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_543),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_449),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_441),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_656),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_441),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_655),
.Y(n_734)
);

CKINVDCx14_ASAP7_75t_R g735 ( 
.A(n_679),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_505),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_505),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_551),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_649),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_638),
.Y(n_740)
);

CKINVDCx16_ASAP7_75t_R g741 ( 
.A(n_438),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_542),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_551),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_574),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_477),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_574),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_595),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_595),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_442),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_442),
.Y(n_750)
);

INVxp33_ASAP7_75t_SL g751 ( 
.A(n_401),
.Y(n_751)
);

CKINVDCx14_ASAP7_75t_R g752 ( 
.A(n_664),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_454),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_481),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_484),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_685),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_486),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_465),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_438),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_486),
.Y(n_761)
);

INVxp67_ASAP7_75t_SL g762 ( 
.A(n_416),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_398),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_408),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_413),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_419),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_421),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_487),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_488),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_431),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_434),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_701),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_483),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_418),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_450),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_452),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_453),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_449),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_489),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_438),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_473),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_476),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_479),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_499),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_480),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_519),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_490),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_494),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_497),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_501),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_509),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_503),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_523),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_527),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_456),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_449),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_538),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_507),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_556),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_456),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_562),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_565),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_496),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_567),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_502),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_575),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_588),
.Y(n_807)
);

INVxp33_ASAP7_75t_SL g808 ( 
.A(n_401),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_449),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_592),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_420),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_510),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_596),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_597),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_599),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_610),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_612),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_519),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_402),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_614),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_519),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_504),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_449),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_506),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_618),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_624),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_429),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_511),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_627),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_629),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_651),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_654),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_674),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_676),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_433),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_678),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_568),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_686),
.Y(n_838)
);

INVxp33_ASAP7_75t_SL g839 ( 
.A(n_402),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_406),
.Y(n_841)
);

CKINVDCx16_ASAP7_75t_R g842 ( 
.A(n_568),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_512),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_518),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_406),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_436),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_719),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_758),
.B(n_496),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_732),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_722),
.Y(n_850)
);

OA21x2_ASAP7_75t_L g851 ( 
.A1(n_705),
.A2(n_634),
.B(n_513),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_719),
.Y(n_852)
);

CKINVDCx8_ASAP7_75t_R g853 ( 
.A(n_724),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_732),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_721),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_752),
.A2(n_521),
.B1(n_684),
.B2(n_399),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_721),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_725),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_722),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_723),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_SL g861 ( 
.A1(n_753),
.A2(n_544),
.B1(n_548),
.B2(n_485),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_761),
.B(n_513),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_725),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_722),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_705),
.A2(n_646),
.B(n_634),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_708),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_726),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_723),
.B(n_564),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_722),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_726),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_727),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_720),
.B(n_646),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_727),
.Y(n_873)
);

OAI22x1_ASAP7_75t_SL g874 ( 
.A1(n_759),
.A2(n_641),
.B1(n_663),
.B2(n_609),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_745),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_722),
.Y(n_876)
);

OA21x2_ASAP7_75t_L g877 ( 
.A1(n_707),
.A2(n_448),
.B(n_444),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_707),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_745),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_709),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_795),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_846),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_711),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_714),
.A2(n_469),
.B(n_463),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_773),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_709),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_735),
.B(n_478),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_749),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_749),
.B(n_440),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_491),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_710),
.Y(n_892)
);

AND2x6_ASAP7_75t_L g893 ( 
.A(n_730),
.B(n_405),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_730),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_712),
.A2(n_404),
.B1(n_409),
.B2(n_403),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_795),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_778),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_713),
.A2(n_404),
.B1(n_409),
.B2(n_403),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_795),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_717),
.Y(n_900)
);

OA21x2_ASAP7_75t_L g901 ( 
.A1(n_778),
.A2(n_493),
.B(n_492),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_706),
.A2(n_412),
.B1(n_415),
.B2(n_410),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_734),
.B(n_460),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_754),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_728),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_728),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_754),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_800),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_800),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_800),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_820),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_755),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_805),
.Y(n_913)
);

AND2x6_ASAP7_75t_L g914 ( 
.A(n_796),
.B(n_405),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_796),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_716),
.A2(n_412),
.B1(n_415),
.B2(n_410),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_SL g917 ( 
.A1(n_715),
.A2(n_423),
.B1(n_430),
.B2(n_426),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_762),
.B(n_498),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_820),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_742),
.A2(n_423),
.B1(n_430),
.B2(n_426),
.Y(n_920)
);

OAI22x1_ASAP7_75t_R g921 ( 
.A1(n_718),
.A2(n_417),
.B1(n_437),
.B2(n_435),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_741),
.B(n_460),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_809),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_774),
.B(n_530),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_811),
.B(n_537),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_822),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_803),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_827),
.B(n_541),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_825),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_809),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_823),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_835),
.B(n_550),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_823),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_803),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_803),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_729),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_729),
.Y(n_937)
);

AND2x2_ASAP7_75t_SL g938 ( 
.A(n_819),
.B(n_405),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_750),
.B(n_560),
.Y(n_939)
);

NOR2x1_ASAP7_75t_L g940 ( 
.A(n_824),
.B(n_425),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_825),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_826),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_731),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_731),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_826),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_755),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_733),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_750),
.A2(n_584),
.B(n_570),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_756),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_819),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_829),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_733),
.Y(n_952)
);

CKINVDCx6p67_ASAP7_75t_R g953 ( 
.A(n_786),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_829),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_736),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_736),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_756),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_831),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_751),
.A2(n_437),
.B1(n_447),
.B2(n_435),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_768),
.B(n_580),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_757),
.B(n_440),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_757),
.B(n_841),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_737),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_768),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_737),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_769),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_738),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_738),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_841),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_878),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_878),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_886),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_913),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_881),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_926),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_966),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_960),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_859),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_966),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_866),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_938),
.B(n_769),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_881),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_950),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_887),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_938),
.B(n_818),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_953),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_866),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_953),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_853),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_887),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_853),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_964),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_950),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_950),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_859),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_866),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_875),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_875),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_879),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_879),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_907),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_907),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_950),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_868),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_912),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_880),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_946),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_892),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_860),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_892),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_904),
.B(n_739),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_860),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_904),
.Y(n_1013)
);

XOR2xp5_ASAP7_75t_L g1014 ( 
.A(n_874),
.B(n_772),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_849),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_854),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_938),
.B(n_779),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_880),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_874),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_889),
.B(n_743),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_861),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_861),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_921),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_921),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_889),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_888),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_903),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_889),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_949),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_918),
.B(n_779),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_922),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_856),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_895),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_949),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_R g1035 ( 
.A(n_877),
.B(n_784),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_895),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_917),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_917),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_916),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_924),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_925),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_859),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_928),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_959),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_949),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_957),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_880),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_920),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_959),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_932),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_R g1051 ( 
.A(n_848),
.B(n_784),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_883),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_902),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_883),
.Y(n_1054)
);

BUFx10_ASAP7_75t_L g1055 ( 
.A(n_891),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_883),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_957),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_862),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_957),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_902),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_900),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_859),
.Y(n_1062)
);

XOR2xp5_ASAP7_75t_L g1063 ( 
.A(n_940),
.B(n_790),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_898),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_898),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_900),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_962),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_969),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_859),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_969),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_859),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_969),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_939),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_864),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_890),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_890),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_961),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_847),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_962),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_923),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_911),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_961),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_911),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_891),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_864),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_891),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_940),
.B(n_751),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_847),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_919),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_891),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_877),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_919),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_929),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_929),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_941),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_941),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_SL g1097 ( 
.A(n_872),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_872),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_942),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_872),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_942),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_855),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_877),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_945),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_872),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_877),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_901),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_945),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_SL g1109 ( 
.A(n_951),
.B(n_790),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_951),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_954),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_954),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_901),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_855),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_958),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_958),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_936),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_936),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_863),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_882),
.B(n_808),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_936),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_936),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_864),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_882),
.B(n_792),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_936),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_885),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_943),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_864),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_936),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_943),
.B(n_743),
.Y(n_1130)
);

NOR2xp67_ASAP7_75t_L g1131 ( 
.A(n_882),
.B(n_792),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_937),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_901),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_885),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_937),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_901),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_956),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_937),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_937),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_944),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1058),
.B(n_882),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1139),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1098),
.B(n_1067),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1079),
.B(n_905),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1055),
.Y(n_1145)
);

AO21x2_ASAP7_75t_L g1146 ( 
.A1(n_981),
.A2(n_948),
.B(n_598),
.Y(n_1146)
);

AND2x6_ASAP7_75t_L g1147 ( 
.A(n_1126),
.B(n_405),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1020),
.Y(n_1148)
);

INVxp33_ASAP7_75t_SL g1149 ( 
.A(n_1011),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_977),
.B(n_808),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1020),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1040),
.B(n_839),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1092),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1029),
.B(n_905),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1041),
.B(n_909),
.Y(n_1155)
);

INVx4_ASAP7_75t_SL g1156 ( 
.A(n_1097),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1025),
.B(n_906),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1043),
.B(n_798),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1028),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1068),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1126),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1070),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_1087),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1050),
.B(n_909),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1073),
.B(n_909),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1017),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_1134),
.B(n_475),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1134),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1107),
.A2(n_602),
.B1(n_668),
.B2(n_639),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1026),
.B(n_839),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_980),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1034),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1075),
.B(n_798),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1001),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_980),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1055),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1055),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1045),
.B(n_906),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1113),
.B(n_909),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_983),
.B(n_760),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_SL g1181 ( 
.A(n_1133),
.B(n_500),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1120),
.B(n_927),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1127),
.B(n_927),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1046),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1136),
.B(n_927),
.Y(n_1185)
);

NOR2x1p5_ASAP7_75t_L g1186 ( 
.A(n_993),
.B(n_812),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1093),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1108),
.B(n_927),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_SL g1189 ( 
.A(n_1004),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1057),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1111),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_987),
.Y(n_1192)
);

BUFx4f_ASAP7_75t_L g1193 ( 
.A(n_1008),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1082),
.B(n_812),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1081),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1076),
.B(n_828),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1083),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_987),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1109),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1108),
.B(n_475),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1100),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_996),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1089),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1137),
.B(n_586),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_996),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1096),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1077),
.B(n_828),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_970),
.B(n_923),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_971),
.B(n_923),
.Y(n_1209)
);

INVx4_ASAP7_75t_SL g1210 ( 
.A(n_1097),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1006),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_978),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1100),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_974),
.B(n_923),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_982),
.B(n_923),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_SL g1216 ( 
.A(n_993),
.B(n_994),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1101),
.Y(n_1217)
);

BUFx8_ASAP7_75t_SL g1218 ( 
.A(n_1023),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_978),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1006),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_984),
.B(n_923),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1013),
.B(n_843),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1105),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1018),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1105),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1104),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1094),
.Y(n_1227)
);

AND2x6_ASAP7_75t_L g1228 ( 
.A(n_1124),
.B(n_475),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1110),
.B(n_843),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1112),
.B(n_615),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1018),
.Y(n_1231)
);

AND2x2_ASAP7_75t_SL g1232 ( 
.A(n_1115),
.B(n_475),
.Y(n_1232)
);

AO22x2_ASAP7_75t_L g1233 ( 
.A1(n_985),
.A2(n_545),
.B1(n_500),
.B2(n_535),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1047),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1116),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_972),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1130),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1095),
.B(n_844),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1110),
.B(n_844),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1130),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1099),
.B(n_475),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1097),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_990),
.B(n_930),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1131),
.B(n_635),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1010),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1061),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1084),
.B(n_621),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1072),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1047),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_978),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_978),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1066),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1078),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1078),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1086),
.B(n_632),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_972),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1088),
.Y(n_1257)
);

AO22x2_ASAP7_75t_L g1258 ( 
.A1(n_1014),
.A2(n_1063),
.B1(n_545),
.B2(n_1060),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1090),
.B(n_637),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1039),
.B(n_740),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1035),
.B(n_821),
.C(n_780),
.Y(n_1261)
);

NOR2x1p5_ASAP7_75t_L g1262 ( 
.A(n_994),
.B(n_447),
.Y(n_1262)
);

NOR2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1003),
.B(n_455),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1059),
.B(n_842),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1088),
.Y(n_1265)
);

AND2x6_ASAP7_75t_L g1266 ( 
.A(n_995),
.B(n_635),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1102),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1052),
.B(n_642),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1102),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1091),
.B(n_1103),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1114),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_978),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1117),
.B(n_930),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1114),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1117),
.Y(n_1275)
);

NAND2xp33_ASAP7_75t_L g1276 ( 
.A(n_1106),
.B(n_449),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1080),
.B(n_851),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1054),
.B(n_645),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_L g1279 ( 
.A(n_1118),
.B(n_1121),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1119),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1064),
.A2(n_865),
.B1(n_851),
.B2(n_948),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1119),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_SL g1283 ( 
.A(n_992),
.B(n_460),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1118),
.B(n_930),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_995),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1030),
.B(n_635),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1121),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_997),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_995),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1122),
.B(n_930),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1056),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1065),
.B(n_837),
.C(n_522),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1004),
.B(n_830),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1122),
.B(n_635),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1042),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1042),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1042),
.Y(n_1297)
);

AND2x6_ASAP7_75t_L g1298 ( 
.A(n_1062),
.B(n_635),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1062),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_991),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1004),
.B(n_834),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1125),
.B(n_930),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1062),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1085),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1125),
.B(n_930),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1129),
.A2(n_691),
.B1(n_652),
.B2(n_657),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1085),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1048),
.B(n_414),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1085),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1021),
.A2(n_865),
.B1(n_851),
.B2(n_619),
.Y(n_1310)
);

AND2x6_ASAP7_75t_L g1311 ( 
.A(n_1123),
.B(n_648),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1069),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1123),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1129),
.B(n_933),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1132),
.Y(n_1315)
);

AND2x2_ASAP7_75t_SL g1316 ( 
.A(n_1080),
.B(n_662),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1132),
.B(n_933),
.Y(n_1317)
);

AND2x6_ASAP7_75t_L g1318 ( 
.A(n_1123),
.B(n_682),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1140),
.A2(n_865),
.B(n_851),
.Y(n_1319)
);

INVx5_ASAP7_75t_L g1320 ( 
.A(n_1069),
.Y(n_1320)
);

NAND2xp33_ASAP7_75t_L g1321 ( 
.A(n_1135),
.B(n_449),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1051),
.B(n_845),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1022),
.A2(n_865),
.B1(n_427),
.B2(n_600),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1128),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_998),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1135),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1015),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1128),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1069),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1128),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1138),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_999),
.B(n_845),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1048),
.A2(n_514),
.B1(n_515),
.B2(n_508),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1138),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1000),
.B(n_568),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1053),
.A2(n_600),
.B1(n_449),
.B2(n_687),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1160),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1327),
.B(n_973),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1253),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1177),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1270),
.A2(n_1031),
.B1(n_1027),
.B2(n_1032),
.Y(n_1341)
);

INVx8_ASAP7_75t_L g1342 ( 
.A(n_1143),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1193),
.B(n_1005),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1253),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1165),
.B(n_1080),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1155),
.B(n_1074),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1164),
.B(n_1074),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1193),
.B(n_1275),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1270),
.A2(n_1007),
.B1(n_1002),
.B2(n_1016),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1236),
.B(n_1256),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1150),
.B(n_1009),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_SL g1352 ( 
.A(n_1180),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1267),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1141),
.B(n_1074),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1174),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1150),
.B(n_1012),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_L g1357 ( 
.A1(n_1244),
.A2(n_688),
.B(n_695),
.C(n_967),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1275),
.B(n_989),
.Y(n_1358)
);

INVx4_ASAP7_75t_L g1359 ( 
.A(n_1177),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1267),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1308),
.A2(n_1049),
.B(n_1044),
.C(n_989),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1279),
.A2(n_1071),
.B(n_1069),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1152),
.B(n_992),
.C(n_1033),
.Y(n_1363)
);

AND2x2_ASAP7_75t_SL g1364 ( 
.A(n_1316),
.B(n_937),
.Y(n_1364)
);

OAI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1336),
.A2(n_1038),
.B1(n_1037),
.B2(n_1036),
.C(n_525),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1177),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1152),
.B(n_973),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1143),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1143),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1293),
.B(n_975),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1178),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1149),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1178),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1336),
.A2(n_600),
.B1(n_605),
.B2(n_459),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1301),
.B(n_975),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1308),
.B(n_986),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1269),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1170),
.B(n_1019),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1156),
.B(n_763),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1170),
.B(n_976),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1177),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1332),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1183),
.B(n_1074),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1323),
.A2(n_1316),
.B1(n_1233),
.B2(n_1276),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1331),
.B(n_1334),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_SL g1386 ( 
.A(n_1288),
.B(n_976),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1237),
.B(n_1069),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1269),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1310),
.A2(n_411),
.B1(n_422),
.B2(n_407),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1229),
.B(n_979),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1240),
.B(n_1074),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1287),
.B(n_986),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1276),
.A2(n_517),
.B1(n_528),
.B2(n_516),
.Y(n_1393)
);

BUFx8_ASAP7_75t_L g1394 ( 
.A(n_1189),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1287),
.B(n_979),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1158),
.B(n_988),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_L g1397 ( 
.A(n_1153),
.B(n_764),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1260),
.A2(n_967),
.B(n_411),
.C(n_422),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1323),
.A2(n_600),
.B1(n_605),
.B2(n_459),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1315),
.B(n_407),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1271),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1300),
.A2(n_1024),
.B1(n_461),
.B2(n_462),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1271),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1148),
.B(n_1071),
.Y(n_1404)
);

O2A1O1Ixp5_ASAP7_75t_L g1405 ( 
.A1(n_1244),
.A2(n_967),
.B(n_857),
.C(n_858),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1160),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1229),
.B(n_520),
.Y(n_1407)
);

NOR2xp67_ASAP7_75t_L g1408 ( 
.A(n_1187),
.B(n_1227),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1239),
.B(n_524),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1178),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1144),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1151),
.B(n_1071),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1310),
.B(n_1071),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1315),
.B(n_428),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1239),
.B(n_1260),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1261),
.B(n_526),
.Y(n_1416)
);

INVxp33_ASAP7_75t_L g1417 ( 
.A(n_1335),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1195),
.B(n_1071),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1144),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1169),
.A2(n_462),
.B1(n_464),
.B2(n_461),
.C(n_455),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1161),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1282),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1197),
.B(n_937),
.Y(n_1423)
);

AND2x4_ASAP7_75t_SL g1424 ( 
.A(n_1300),
.B(n_605),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1200),
.A2(n_1185),
.B(n_1179),
.C(n_1241),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1245),
.A2(n_967),
.B(n_432),
.C(n_439),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1203),
.B(n_884),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1196),
.B(n_765),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1206),
.B(n_1217),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1233),
.A2(n_600),
.B1(n_470),
.B2(n_554),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1179),
.A2(n_432),
.B1(n_439),
.B2(n_428),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1226),
.B(n_884),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1326),
.B(n_443),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1163),
.B(n_529),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1235),
.B(n_934),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1326),
.B(n_443),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1279),
.B(n_934),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_SL g1438 ( 
.A(n_1325),
.B(n_445),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1163),
.B(n_445),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1161),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1144),
.B(n_934),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1189),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1156),
.B(n_766),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1182),
.B(n_934),
.Y(n_1444)
);

NOR2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1201),
.B(n_464),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1162),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1207),
.B(n_1142),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1257),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1185),
.A2(n_539),
.B1(n_546),
.B2(n_533),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1248),
.B(n_446),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1238),
.B(n_531),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1274),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1188),
.A2(n_561),
.B1(n_566),
.B2(n_549),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1291),
.B(n_1201),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1159),
.B(n_915),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1172),
.B(n_915),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1213),
.B(n_1223),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1264),
.B(n_767),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1162),
.B(n_770),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1280),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1161),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1282),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1171),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1184),
.B(n_915),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1190),
.B(n_852),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1200),
.A2(n_857),
.B(n_858),
.C(n_852),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1322),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1213),
.B(n_446),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1154),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1154),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1154),
.B(n_870),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1223),
.B(n_451),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1233),
.A2(n_1232),
.B1(n_1321),
.B2(n_1161),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1191),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1246),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1173),
.B(n_532),
.Y(n_1476)
);

INVx8_ASAP7_75t_L g1477 ( 
.A(n_1247),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1168),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1252),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1254),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1194),
.B(n_536),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1254),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1199),
.B(n_540),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1204),
.B(n_870),
.Y(n_1484)
);

NAND3xp33_ASAP7_75t_L g1485 ( 
.A(n_1333),
.B(n_552),
.C(n_547),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1204),
.B(n_871),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1232),
.A2(n_600),
.B1(n_554),
.B2(n_557),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1204),
.B(n_871),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1415),
.B(n_1157),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1415),
.A2(n_1181),
.B1(n_1188),
.B2(n_1222),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1383),
.A2(n_1284),
.B(n_1273),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1463),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1351),
.B(n_1166),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1384),
.A2(n_1168),
.B1(n_1176),
.B2(n_1145),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1345),
.A2(n_1305),
.B(n_1290),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1421),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1407),
.B(n_1157),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1461),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1407),
.B(n_1157),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1409),
.A2(n_1241),
.B(n_1306),
.C(n_1286),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1462),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1339),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1364),
.B(n_1168),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1413),
.A2(n_1281),
.B(n_1321),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1346),
.A2(n_1314),
.B(n_1302),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1421),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_SL g1507 ( 
.A(n_1350),
.B(n_1218),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1364),
.B(n_1168),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1347),
.A2(n_1314),
.B(n_1302),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1382),
.B(n_1225),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1409),
.B(n_1268),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1382),
.B(n_1225),
.Y(n_1512)
);

AO21x1_ASAP7_75t_L g1513 ( 
.A1(n_1425),
.A2(n_1294),
.B(n_1286),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1354),
.A2(n_1317),
.B(n_1320),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1351),
.B(n_1264),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1384),
.A2(n_1176),
.B1(n_1145),
.B2(n_1281),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1344),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1355),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1405),
.A2(n_1294),
.B(n_1317),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1444),
.A2(n_1320),
.B(n_1277),
.Y(n_1520)
);

NOR2xp67_ASAP7_75t_L g1521 ( 
.A(n_1372),
.B(n_1292),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1353),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1421),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1467),
.B(n_1429),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1421),
.B(n_1242),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1362),
.A2(n_1320),
.B(n_1277),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_L g1527 ( 
.A(n_1356),
.B(n_1378),
.C(n_1367),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1370),
.B(n_1268),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1467),
.B(n_1268),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1375),
.B(n_1278),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1430),
.A2(n_1181),
.B(n_1283),
.C(n_1230),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1437),
.A2(n_1320),
.B(n_1219),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1342),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1430),
.A2(n_1230),
.B(n_1255),
.C(n_1247),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1441),
.A2(n_1219),
.B(n_1212),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1447),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1387),
.A2(n_1219),
.B(n_1212),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1484),
.B(n_1278),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1473),
.B(n_1242),
.Y(n_1539)
);

AND2x4_ASAP7_75t_SL g1540 ( 
.A(n_1340),
.B(n_1180),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1473),
.B(n_1411),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1356),
.B(n_1278),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1391),
.A2(n_1219),
.B(n_1212),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1404),
.A2(n_1250),
.B(n_1212),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1486),
.B(n_1230),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1340),
.B(n_1250),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1360),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1488),
.B(n_1247),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1461),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1405),
.A2(n_1209),
.B(n_1208),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1367),
.A2(n_1259),
.B1(n_1255),
.B2(n_1262),
.Y(n_1551)
);

INVx3_ASAP7_75t_SL g1552 ( 
.A(n_1442),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1412),
.A2(n_1398),
.B(n_1435),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1419),
.B(n_1471),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1469),
.B(n_1255),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1399),
.A2(n_1258),
.B1(n_1259),
.B2(n_1147),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1377),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1470),
.A2(n_1329),
.B1(n_1328),
.B2(n_1304),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1388),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1478),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1401),
.Y(n_1562)
);

NAND2x1p5_ASAP7_75t_L g1563 ( 
.A(n_1359),
.B(n_1250),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1451),
.B(n_1259),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1403),
.A2(n_1215),
.B(n_1214),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1418),
.A2(n_1251),
.B(n_1250),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1474),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1474),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1422),
.Y(n_1569)
);

BUFx8_ASAP7_75t_L g1570 ( 
.A(n_1446),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1451),
.B(n_1180),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_1363),
.B(n_1221),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1478),
.Y(n_1573)
);

NOR2xp67_ASAP7_75t_L g1574 ( 
.A(n_1338),
.B(n_1243),
.Y(n_1574)
);

INVx11_ASAP7_75t_L g1575 ( 
.A(n_1394),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1368),
.B(n_1156),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1511),
.B(n_1349),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1576),
.B(n_1410),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1576),
.B(n_1369),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1570),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1527),
.A2(n_1376),
.B(n_1390),
.C(n_1380),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1515),
.B(n_1493),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1489),
.B(n_1341),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1522),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1527),
.B(n_1390),
.C(n_1380),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1496),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1497),
.A2(n_1385),
.B1(n_1365),
.B2(n_1361),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1568),
.Y(n_1588)
);

OR2x4_ASAP7_75t_L g1589 ( 
.A(n_1515),
.B(n_1378),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_SL g1590 ( 
.A(n_1564),
.B(n_1420),
.C(n_1386),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1499),
.B(n_1476),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1495),
.A2(n_1348),
.B(n_1272),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1542),
.A2(n_1481),
.B1(n_1476),
.B2(n_1416),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1524),
.B(n_1538),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1545),
.B(n_1428),
.Y(n_1596)
);

CKINVDCx8_ASAP7_75t_R g1597 ( 
.A(n_1533),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1481),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1490),
.B(n_1408),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1493),
.B(n_1417),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1531),
.A2(n_1500),
.B(n_1534),
.C(n_1416),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1557),
.A2(n_1479),
.B1(n_1475),
.B2(n_1342),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1557),
.A2(n_1402),
.B1(n_1399),
.B2(n_1374),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1554),
.B(n_1483),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1491),
.A2(n_1272),
.B(n_1251),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1522),
.Y(n_1606)
);

INVx3_ASAP7_75t_SL g1607 ( 
.A(n_1552),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1504),
.A2(n_1272),
.B(n_1251),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1505),
.A2(n_1272),
.B(n_1251),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1536),
.B(n_1483),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1510),
.B(n_1458),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1534),
.B(n_1477),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1558),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1528),
.B(n_1448),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1503),
.A2(n_1342),
.B1(n_1366),
.B2(n_1359),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1530),
.B(n_1452),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1512),
.B(n_1434),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1558),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1529),
.B(n_1434),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_R g1621 ( 
.A(n_1507),
.B(n_1352),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1501),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1551),
.B(n_1438),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1526),
.A2(n_1319),
.B(n_1423),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1509),
.A2(n_1312),
.B(n_1366),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1520),
.A2(n_1357),
.B(n_1455),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1492),
.Y(n_1627)
);

NAND2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1503),
.B(n_1381),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1533),
.B(n_1381),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1622),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1601),
.A2(n_1516),
.B(n_1494),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1592),
.A2(n_1508),
.B(n_1553),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1607),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1585),
.A2(n_1594),
.B(n_1620),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1582),
.A2(n_1531),
.B(n_1487),
.C(n_1374),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1581),
.A2(n_1487),
.B(n_1541),
.C(n_1508),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1610),
.A2(n_1550),
.B(n_1514),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1597),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1605),
.A2(n_1532),
.B(n_1519),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1622),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1603),
.A2(n_1258),
.B1(n_1571),
.B2(n_1389),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1614),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1598),
.A2(n_1539),
.B(n_1541),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1594),
.B(n_1567),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1587),
.A2(n_1539),
.B(n_1572),
.C(n_1556),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1597),
.Y(n_1646)
);

NAND2x1p5_ASAP7_75t_L g1647 ( 
.A(n_1591),
.B(n_1533),
.Y(n_1647)
);

BUFx2_ASAP7_75t_R g1648 ( 
.A(n_1607),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1595),
.B(n_1518),
.Y(n_1649)
);

OAI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1604),
.A2(n_1485),
.B(n_1216),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1590),
.B(n_1343),
.C(n_1358),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1589),
.A2(n_1457),
.B1(n_1454),
.B2(n_1406),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1596),
.B(n_1396),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1596),
.B(n_1521),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1583),
.A2(n_1258),
.B1(n_1445),
.B2(n_1395),
.Y(n_1655)
);

AOI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1599),
.A2(n_1513),
.B(n_1525),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1577),
.A2(n_1477),
.B(n_1574),
.C(n_1426),
.Y(n_1657)
);

NAND3x1_ASAP7_75t_L g1658 ( 
.A(n_1618),
.B(n_1394),
.C(n_1575),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1603),
.A2(n_1623),
.B1(n_1600),
.B2(n_1611),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1614),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1626),
.A2(n_1565),
.B(n_1357),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1593),
.A2(n_1566),
.B(n_1543),
.Y(n_1662)
);

AOI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1625),
.A2(n_1525),
.B(n_1537),
.Y(n_1663)
);

AOI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1609),
.A2(n_1544),
.B(n_1559),
.Y(n_1664)
);

AO21x1_ASAP7_75t_L g1665 ( 
.A1(n_1602),
.A2(n_1555),
.B(n_1431),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1615),
.B(n_1397),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1459),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1591),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1588),
.Y(n_1669)
);

AO31x2_ASAP7_75t_L g1670 ( 
.A1(n_1584),
.A2(n_1535),
.A3(n_1517),
.B(n_1502),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1612),
.A2(n_1393),
.B(n_1449),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1624),
.A2(n_1626),
.B(n_1628),
.Y(n_1672)
);

AO32x2_ASAP7_75t_L g1673 ( 
.A1(n_1616),
.A2(n_1146),
.A3(n_1466),
.B1(n_1228),
.B2(n_1555),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1613),
.A2(n_1477),
.B(n_1546),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1627),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1624),
.A2(n_1464),
.B(n_1456),
.Y(n_1676)
);

O2A1O1Ixp33_ASAP7_75t_SL g1677 ( 
.A1(n_1584),
.A2(n_1400),
.B(n_1433),
.C(n_1414),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1613),
.A2(n_1563),
.B(n_1546),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1606),
.A2(n_1146),
.B(n_1465),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1659),
.B(n_1608),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1634),
.B(n_1588),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1641),
.A2(n_1439),
.B1(n_1459),
.B2(n_1613),
.Y(n_1682)
);

BUFx4f_ASAP7_75t_L g1683 ( 
.A(n_1646),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1635),
.A2(n_1617),
.B(n_1589),
.C(n_1540),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1630),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1637),
.A2(n_1619),
.B(n_1606),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1639),
.A2(n_1619),
.B(n_1432),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_SL g1688 ( 
.A1(n_1665),
.A2(n_1627),
.B(n_1591),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1641),
.A2(n_1659),
.B1(n_1635),
.B2(n_1631),
.C(n_1636),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1672),
.A2(n_1628),
.B(n_1586),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1642),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

CKINVDCx6p67_ASAP7_75t_R g1694 ( 
.A(n_1638),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1662),
.A2(n_1628),
.B(n_1586),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1675),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1649),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1617),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1670),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1645),
.A2(n_1436),
.B(n_1450),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

AOI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1664),
.A2(n_1613),
.B(n_1392),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1663),
.A2(n_1676),
.B(n_1656),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1644),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1632),
.A2(n_1427),
.B(n_1460),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1669),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1651),
.B(n_1453),
.C(n_1468),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1655),
.A2(n_1589),
.B1(n_1263),
.B2(n_1186),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1670),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1670),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1678),
.A2(n_1586),
.B(n_1440),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1674),
.B(n_1629),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1679),
.Y(n_1713)
);

OAI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1643),
.A2(n_1440),
.B(n_1563),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1661),
.A2(n_1175),
.B(n_1171),
.Y(n_1715)
);

OR2x6_ASAP7_75t_L g1716 ( 
.A(n_1645),
.B(n_1629),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1650),
.A2(n_1459),
.B1(n_1472),
.B2(n_1578),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1661),
.A2(n_1192),
.B(n_1175),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1644),
.B(n_1579),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1661),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1648),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1654),
.Y(n_1723)
);

OA21x2_ASAP7_75t_L g1724 ( 
.A1(n_1636),
.A2(n_1560),
.B(n_1547),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1657),
.A2(n_1569),
.B(n_1562),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1667),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1666),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1671),
.A2(n_1424),
.B1(n_1621),
.B2(n_1540),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1652),
.A2(n_1578),
.B1(n_1579),
.B2(n_1443),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1638),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1646),
.A2(n_1578),
.B1(n_1579),
.B2(n_1443),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1633),
.A2(n_1379),
.B1(n_1337),
.B2(n_1607),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1673),
.B(n_600),
.Y(n_1733)
);

BUFx12f_ASAP7_75t_L g1734 ( 
.A(n_1633),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1673),
.B(n_600),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1668),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1677),
.B(n_1218),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1668),
.A2(n_1198),
.B(n_1192),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1647),
.A2(n_1202),
.B(n_1198),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1673),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_SL g1741 ( 
.A1(n_1677),
.A2(n_1482),
.B(n_1480),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1658),
.A2(n_1580),
.B1(n_1552),
.B2(n_1379),
.Y(n_1742)
);

BUFx2_ASAP7_75t_SL g1743 ( 
.A(n_1658),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1657),
.A2(n_1580),
.B1(n_1570),
.B2(n_1629),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1647),
.B(n_1496),
.Y(n_1745)
);

CKINVDCx6p67_ASAP7_75t_R g1746 ( 
.A(n_1673),
.Y(n_1746)
);

AO21x2_ASAP7_75t_L g1747 ( 
.A1(n_1662),
.A2(n_1297),
.B(n_1296),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1672),
.A2(n_1205),
.B(n_1202),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1672),
.A2(n_1211),
.B(n_1205),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1659),
.B(n_553),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1630),
.Y(n_1751)
);

OAI21x1_ASAP7_75t_L g1752 ( 
.A1(n_1672),
.A2(n_1220),
.B(n_1211),
.Y(n_1752)
);

NAND2xp33_ASAP7_75t_R g1753 ( 
.A(n_1633),
.B(n_1498),
.Y(n_1753)
);

OAI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1655),
.A2(n_557),
.B1(n_558),
.B2(n_470),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1659),
.B(n_559),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1638),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1672),
.A2(n_1224),
.B(n_1220),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1672),
.A2(n_1231),
.B(n_1224),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1659),
.B(n_563),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_SL g1760 ( 
.A1(n_1665),
.A2(n_1289),
.B(n_1285),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1632),
.A2(n_1549),
.B(n_1498),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1672),
.A2(n_1234),
.B(n_1231),
.Y(n_1762)
);

OA21x2_ASAP7_75t_L g1763 ( 
.A1(n_1637),
.A2(n_873),
.B(n_746),
.Y(n_1763)
);

OAI21x1_ASAP7_75t_L g1764 ( 
.A1(n_1672),
.A2(n_1249),
.B(n_1234),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1642),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1704),
.B(n_831),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1693),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1692),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1689),
.B(n_1496),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1756),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1700),
.A2(n_1561),
.B(n_1549),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1703),
.A2(n_746),
.B(n_744),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1736),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1754),
.A2(n_631),
.B1(n_633),
.B2(n_628),
.C(n_558),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1707),
.A2(n_775),
.B(n_771),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1756),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1722),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1692),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1712),
.B(n_1765),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1684),
.A2(n_458),
.B(n_466),
.C(n_451),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1765),
.Y(n_1781)
);

BUFx12f_ASAP7_75t_L g1782 ( 
.A(n_1734),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1736),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1685),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1691),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1723),
.B(n_569),
.Y(n_1786)
);

AOI21x1_ASAP7_75t_L g1787 ( 
.A1(n_1702),
.A2(n_777),
.B(n_776),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1703),
.A2(n_747),
.B(n_744),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1694),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1681),
.B(n_832),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1701),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1750),
.A2(n_631),
.B1(n_633),
.B2(n_628),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1751),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1697),
.B(n_571),
.Y(n_1794)
);

OAI21x1_ASAP7_75t_L g1795 ( 
.A1(n_1702),
.A2(n_1561),
.B(n_1573),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1727),
.B(n_572),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1696),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1755),
.A2(n_644),
.B1(n_650),
.B2(n_636),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1737),
.A2(n_782),
.B1(n_783),
.B2(n_781),
.Y(n_1799)
);

AO21x2_ASAP7_75t_L g1800 ( 
.A1(n_1741),
.A2(n_833),
.B(n_832),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1681),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1759),
.A2(n_787),
.B(n_785),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1680),
.B(n_833),
.Y(n_1803)
);

A2O1A1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1684),
.A2(n_466),
.B(n_467),
.C(n_458),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1761),
.A2(n_1573),
.B(n_1506),
.Y(n_1805)
);

CKINVDCx11_ASAP7_75t_R g1806 ( 
.A(n_1734),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1716),
.A2(n_1506),
.B(n_1496),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1686),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1688),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1726),
.B(n_747),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1713),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1686),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1694),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1713),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1699),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1699),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1686),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1736),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1716),
.A2(n_1523),
.B(n_1506),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1698),
.B(n_576),
.Y(n_1820)
);

O2A1O1Ixp5_ASAP7_75t_L g1821 ( 
.A1(n_1733),
.A2(n_1735),
.B(n_1683),
.C(n_1740),
.Y(n_1821)
);

AO21x2_ASAP7_75t_L g1822 ( 
.A1(n_1741),
.A2(n_838),
.B(n_836),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1682),
.A2(n_468),
.B(n_471),
.C(n_467),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1712),
.B(n_1506),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1709),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1709),
.Y(n_1826)
);

BUFx8_ASAP7_75t_SL g1827 ( 
.A(n_1683),
.Y(n_1827)
);

NAND2x1p5_ASAP7_75t_L g1828 ( 
.A(n_1725),
.B(n_1523),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1720),
.B(n_748),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1716),
.A2(n_1725),
.B(n_1683),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1744),
.B(n_836),
.Y(n_1831)
);

OA21x2_ASAP7_75t_L g1832 ( 
.A1(n_1721),
.A2(n_748),
.B(n_838),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1710),
.Y(n_1833)
);

A2O1A1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1733),
.A2(n_471),
.B(n_474),
.C(n_468),
.Y(n_1834)
);

OA21x2_ASAP7_75t_L g1835 ( 
.A1(n_1721),
.A2(n_840),
.B(n_789),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_SL g1836 ( 
.A1(n_1688),
.A2(n_840),
.B(n_791),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1715),
.A2(n_1265),
.B(n_1304),
.Y(n_1837)
);

OA21x2_ASAP7_75t_L g1838 ( 
.A1(n_1717),
.A2(n_793),
.B(n_788),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1716),
.A2(n_1523),
.B(n_1312),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1706),
.B(n_956),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1701),
.Y(n_1841)
);

OR2x6_ASAP7_75t_L g1842 ( 
.A(n_1712),
.B(n_1523),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1730),
.B(n_794),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1735),
.B(n_577),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1736),
.B(n_579),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1736),
.B(n_581),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1745),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1745),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1710),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1717),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_L g1851 ( 
.A1(n_1715),
.A2(n_1265),
.B(n_1328),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1718),
.B(n_582),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1724),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1724),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1712),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1724),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1728),
.A2(n_799),
.B1(n_801),
.B2(n_797),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1745),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1719),
.A2(n_1289),
.B(n_1285),
.Y(n_1859)
);

AOI21x1_ASAP7_75t_L g1860 ( 
.A1(n_1760),
.A2(n_804),
.B(n_802),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1687),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1746),
.B(n_806),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1708),
.B(n_585),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1687),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1725),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1687),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1705),
.A2(n_1312),
.B(n_1249),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1729),
.A2(n_644),
.B1(n_650),
.B2(n_636),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1746),
.B(n_807),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1705),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1690),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1705),
.A2(n_1747),
.B(n_1695),
.Y(n_1872)
);

OAI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1719),
.A2(n_1299),
.B(n_1295),
.Y(n_1873)
);

AO31x2_ASAP7_75t_L g1874 ( 
.A1(n_1760),
.A2(n_873),
.A3(n_1309),
.B(n_1303),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1747),
.B(n_810),
.Y(n_1875)
);

AO21x2_ASAP7_75t_L g1876 ( 
.A1(n_1747),
.A2(n_814),
.B(n_813),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1743),
.B(n_1732),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1748),
.A2(n_816),
.B(n_815),
.Y(n_1878)
);

CKINVDCx16_ASAP7_75t_R g1879 ( 
.A(n_1753),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1711),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1690),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1711),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1743),
.A2(n_659),
.B1(n_661),
.B2(n_658),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1695),
.B(n_817),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1763),
.Y(n_1885)
);

OA21x2_ASAP7_75t_L g1886 ( 
.A1(n_1748),
.A2(n_965),
.B(n_963),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1714),
.A2(n_1312),
.B(n_1299),
.Y(n_1887)
);

OAI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1749),
.A2(n_1307),
.B(n_1295),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1731),
.A2(n_1228),
.B(n_1311),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1763),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1763),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1745),
.Y(n_1892)
);

INVx6_ASAP7_75t_L g1893 ( 
.A(n_1742),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1714),
.A2(n_659),
.B1(n_661),
.B2(n_658),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1749),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1752),
.B(n_587),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1739),
.A2(n_1330),
.B(n_1307),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1739),
.A2(n_1330),
.B(n_555),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1738),
.Y(n_1899)
);

AOI211xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1738),
.A2(n_965),
.B(n_968),
.C(n_963),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1752),
.A2(n_1228),
.B(n_1311),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1757),
.A2(n_965),
.B(n_963),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1757),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1758),
.A2(n_667),
.B1(n_669),
.B2(n_666),
.Y(n_1904)
);

OAI21x1_ASAP7_75t_L g1905 ( 
.A1(n_1758),
.A2(n_968),
.B(n_1313),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1762),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1762),
.B(n_968),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1764),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1764),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1726),
.B(n_0),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1700),
.A2(n_555),
.B(n_474),
.Y(n_1911)
);

A2O1A1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1689),
.A2(n_643),
.B(n_647),
.C(n_640),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1700),
.A2(n_643),
.B(n_640),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1689),
.A2(n_667),
.B1(n_669),
.B2(n_666),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1693),
.Y(n_1915)
);

INVx4_ASAP7_75t_L g1916 ( 
.A(n_1694),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1811),
.Y(n_1917)
);

INVxp67_ASAP7_75t_SL g1918 ( 
.A(n_1801),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1778),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1814),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1767),
.Y(n_1921)
);

BUFx3_ASAP7_75t_L g1922 ( 
.A(n_1789),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1915),
.Y(n_1923)
);

INVxp33_ASAP7_75t_L g1924 ( 
.A(n_1806),
.Y(n_1924)
);

INVx4_ASAP7_75t_SL g1925 ( 
.A(n_1893),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1768),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1784),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1791),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1791),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1779),
.B(n_0),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1785),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1781),
.Y(n_1932)
);

CKINVDCx12_ASAP7_75t_R g1933 ( 
.A(n_1829),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1779),
.B(n_1),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1790),
.B(n_589),
.Y(n_1935)
);

AO31x2_ASAP7_75t_L g1936 ( 
.A1(n_1865),
.A2(n_867),
.A3(n_863),
.B(n_908),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1793),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1808),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1797),
.Y(n_1939)
);

INVx2_ASAP7_75t_SL g1940 ( 
.A(n_1776),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1773),
.Y(n_1941)
);

INVx5_ASAP7_75t_L g1942 ( 
.A(n_1827),
.Y(n_1942)
);

INVx2_ASAP7_75t_SL g1943 ( 
.A(n_1776),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1841),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1841),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1808),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1821),
.B(n_1),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1817),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1850),
.Y(n_1949)
);

OR2x6_ASAP7_75t_L g1950 ( 
.A(n_1830),
.B(n_944),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1821),
.B(n_1855),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1809),
.B(n_2),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1776),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1809),
.B(n_2),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1813),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1817),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1815),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1812),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1872),
.A2(n_1324),
.B(n_867),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1842),
.B(n_3),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1787),
.A2(n_1867),
.B(n_1860),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1816),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1862),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1826),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1825),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1826),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1842),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1833),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1773),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1869),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1861),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1861),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1849),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1853),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1854),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1856),
.B(n_4),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1864),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1842),
.B(n_7),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1783),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1770),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1776),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1783),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1866),
.B(n_8),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1864),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1818),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1818),
.Y(n_1986)
);

AO21x2_ASAP7_75t_L g1987 ( 
.A1(n_1885),
.A2(n_910),
.B(n_908),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1835),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_SL g1989 ( 
.A1(n_1792),
.A2(n_9),
.B(n_11),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1835),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1858),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1858),
.B(n_9),
.Y(n_1992)
);

NAND2x1_ASAP7_75t_L g1993 ( 
.A(n_1838),
.B(n_1147),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1870),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1870),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1866),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1847),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1892),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1835),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_SL g2000 ( 
.A1(n_1879),
.A2(n_672),
.B1(n_673),
.B2(n_671),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1890),
.A2(n_935),
.B(n_910),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1832),
.Y(n_2002)
);

INVx4_ASAP7_75t_L g2003 ( 
.A(n_1916),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1832),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1838),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1838),
.Y(n_2006)
);

CKINVDCx14_ASAP7_75t_R g2007 ( 
.A(n_1806),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1810),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1790),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1832),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1871),
.B(n_11),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1881),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1828),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1828),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1884),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1891),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1892),
.B(n_12),
.Y(n_2017)
);

OA21x2_ASAP7_75t_L g2018 ( 
.A1(n_1891),
.A2(n_653),
.B(n_647),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1847),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1880),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1882),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1895),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1903),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1909),
.Y(n_2024)
);

AO21x2_ASAP7_75t_L g2025 ( 
.A1(n_1836),
.A2(n_935),
.B(n_1228),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1875),
.Y(n_2026)
);

OA21x2_ASAP7_75t_L g2027 ( 
.A1(n_1908),
.A2(n_660),
.B(n_653),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1908),
.Y(n_2028)
);

OR2x6_ASAP7_75t_L g2029 ( 
.A(n_1839),
.B(n_944),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1824),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1848),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1906),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_1800),
.A2(n_1822),
.B(n_1876),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1906),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1782),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1899),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1848),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1876),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1907),
.Y(n_2039)
);

AO21x2_ASAP7_75t_L g2040 ( 
.A1(n_1800),
.A2(n_1228),
.B(n_1167),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1766),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_SL g2042 ( 
.A1(n_1912),
.A2(n_672),
.B(n_671),
.Y(n_2042)
);

AOI21x1_ASAP7_75t_L g2043 ( 
.A1(n_1896),
.A2(n_1167),
.B(n_1147),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1874),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_1766),
.Y(n_2045)
);

OAI21x1_ASAP7_75t_L g2046 ( 
.A1(n_1837),
.A2(n_876),
.B(n_850),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1874),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1772),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1772),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_1824),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1844),
.B(n_13),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1916),
.B(n_14),
.Y(n_2052)
);

AO21x1_ASAP7_75t_SL g2053 ( 
.A1(n_1894),
.A2(n_1210),
.B(n_14),
.Y(n_2053)
);

NAND2x1_ASAP7_75t_L g2054 ( 
.A(n_1893),
.B(n_1147),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1874),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1803),
.B(n_590),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1777),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1874),
.Y(n_2058)
);

BUFx2_ASAP7_75t_L g2059 ( 
.A(n_1822),
.Y(n_2059)
);

AOI221xp5_ASAP7_75t_L g2060 ( 
.A1(n_1989),
.A2(n_1914),
.B1(n_1803),
.B2(n_1798),
.C(n_1792),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_1918),
.B(n_1840),
.Y(n_2061)
);

AOI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1947),
.A2(n_1843),
.B(n_1877),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_2053),
.A2(n_1914),
.B1(n_1893),
.B2(n_1913),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2042),
.A2(n_1912),
.B1(n_1823),
.B2(n_1780),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2009),
.B(n_1834),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2042),
.A2(n_1823),
.B1(n_1780),
.B2(n_1804),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1963),
.B(n_1834),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1970),
.B(n_1820),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_2053),
.A2(n_1911),
.B1(n_1831),
.B2(n_1798),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1947),
.A2(n_1831),
.B1(n_1863),
.B2(n_1889),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2026),
.A2(n_1894),
.B1(n_1883),
.B2(n_1774),
.Y(n_2071)
);

AOI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_2026),
.A2(n_1883),
.B1(n_1852),
.B2(n_1904),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1994),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2051),
.A2(n_1904),
.B1(n_1769),
.B2(n_1827),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_SL g2075 ( 
.A1(n_2007),
.A2(n_1786),
.B1(n_1796),
.B2(n_1799),
.Y(n_2075)
);

A2O1A1Ixp33_ASAP7_75t_L g2076 ( 
.A1(n_1935),
.A2(n_1804),
.B(n_1775),
.C(n_1802),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_2051),
.A2(n_1769),
.B1(n_1868),
.B2(n_1846),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2015),
.A2(n_1845),
.B1(n_1771),
.B2(n_1794),
.Y(n_2078)
);

OAI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2056),
.A2(n_2000),
.B1(n_1950),
.B2(n_1857),
.C(n_2008),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1917),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_2041),
.A2(n_1807),
.B1(n_1819),
.B2(n_1910),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1980),
.B(n_1772),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2050),
.B(n_1788),
.Y(n_2083)
);

AOI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_1960),
.A2(n_1978),
.B1(n_2052),
.B2(n_1950),
.Y(n_2084)
);

OAI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1942),
.A2(n_1900),
.B1(n_1805),
.B2(n_1898),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_1994),
.Y(n_2086)
);

OAI211xp5_ASAP7_75t_L g2087 ( 
.A1(n_2045),
.A2(n_675),
.B(n_677),
.C(n_673),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_2035),
.Y(n_2088)
);

BUFx4f_ASAP7_75t_SL g2089 ( 
.A(n_2035),
.Y(n_2089)
);

OAI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_2027),
.A2(n_1901),
.B(n_1795),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1995),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1917),
.Y(n_2092)
);

OAI221xp5_ASAP7_75t_L g2093 ( 
.A1(n_1950),
.A2(n_681),
.B1(n_683),
.B2(n_677),
.C(n_675),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1933),
.A2(n_1978),
.B1(n_1960),
.B2(n_2052),
.Y(n_2094)
);

AOI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_1952),
.A2(n_689),
.B1(n_693),
.B2(n_683),
.C(n_681),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2030),
.B(n_1788),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1920),
.Y(n_2097)
);

BUFx3_ASAP7_75t_L g2098 ( 
.A(n_1922),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1919),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1920),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1960),
.A2(n_693),
.B1(n_699),
.B2(n_689),
.Y(n_2101)
);

NAND3xp33_ASAP7_75t_L g2102 ( 
.A(n_2027),
.B(n_700),
.C(n_699),
.Y(n_2102)
);

OR2x6_ASAP7_75t_L g2103 ( 
.A(n_1950),
.B(n_1887),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_SL g2104 ( 
.A1(n_2027),
.A2(n_2018),
.B1(n_1942),
.B2(n_1978),
.Y(n_2104)
);

NAND4xp25_ASAP7_75t_L g2105 ( 
.A(n_1952),
.B(n_702),
.C(n_700),
.D(n_1897),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2030),
.B(n_1788),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2030),
.B(n_1878),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_1922),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_2057),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1942),
.A2(n_702),
.B1(n_594),
.B2(n_601),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1927),
.B(n_1878),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1921),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1919),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_SL g2114 ( 
.A1(n_2018),
.A2(n_1878),
.B(n_665),
.Y(n_2114)
);

CKINVDCx11_ASAP7_75t_R g2115 ( 
.A(n_1955),
.Y(n_2115)
);

OAI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1924),
.A2(n_603),
.B1(n_604),
.B2(n_591),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_SL g2117 ( 
.A1(n_2027),
.A2(n_608),
.B1(n_611),
.B2(n_607),
.Y(n_2117)
);

OAI22xp33_ASAP7_75t_L g2118 ( 
.A1(n_1942),
.A2(n_616),
.B1(n_625),
.B2(n_613),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1997),
.B(n_1851),
.Y(n_2119)
);

NAND3xp33_ASAP7_75t_L g2120 ( 
.A(n_2039),
.B(n_626),
.C(n_660),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1955),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1997),
.B(n_1886),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_2052),
.A2(n_1942),
.B1(n_1930),
.B2(n_1934),
.Y(n_2123)
);

OA21x2_ASAP7_75t_L g2124 ( 
.A1(n_1995),
.A2(n_1905),
.B(n_1873),
.Y(n_2124)
);

OAI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_2011),
.A2(n_1951),
.B1(n_2003),
.B2(n_1983),
.C(n_2039),
.Y(n_2125)
);

AO221x2_ASAP7_75t_L g2126 ( 
.A1(n_1944),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.C(n_20),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1932),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1932),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_1954),
.A2(n_680),
.B1(n_690),
.B2(n_670),
.C(n_665),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_1954),
.A2(n_690),
.B1(n_692),
.B2(n_680),
.C(n_670),
.Y(n_2130)
);

OAI211xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2011),
.A2(n_22),
.B(n_18),
.C(n_20),
.Y(n_2131)
);

AOI222xp33_ASAP7_75t_L g2132 ( 
.A1(n_1930),
.A2(n_704),
.B1(n_698),
.B2(n_697),
.C1(n_696),
.C2(n_692),
.Y(n_2132)
);

OAI211xp5_ASAP7_75t_SL g2133 ( 
.A1(n_1983),
.A2(n_27),
.B(n_23),
.C(n_25),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1921),
.B(n_1886),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_1953),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_1942),
.A2(n_1318),
.B1(n_1311),
.B2(n_947),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_2005),
.A2(n_1902),
.B(n_1886),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1934),
.A2(n_1318),
.B1(n_1311),
.B2(n_947),
.Y(n_2138)
);

INVx4_ASAP7_75t_L g2139 ( 
.A(n_2003),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2054),
.A2(n_697),
.B1(n_698),
.B2(n_696),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1923),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1923),
.B(n_1902),
.Y(n_2142)
);

OAI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_1951),
.A2(n_704),
.B1(n_593),
.B2(n_606),
.C(n_583),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_2057),
.Y(n_2144)
);

AOI221xp5_ASAP7_75t_L g2145 ( 
.A1(n_1992),
.A2(n_623),
.B1(n_617),
.B2(n_620),
.C(n_622),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1931),
.Y(n_2146)
);

A2O1A1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_1976),
.A2(n_578),
.B(n_29),
.C(n_23),
.Y(n_2147)
);

OAI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_2003),
.A2(n_2054),
.B1(n_2029),
.B2(n_2018),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1967),
.A2(n_1902),
.B1(n_947),
.B2(n_952),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1931),
.Y(n_2150)
);

AND2x4_ASAP7_75t_L g2151 ( 
.A(n_2019),
.B(n_1859),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1937),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1953),
.Y(n_2153)
);

AOI22xp33_ASAP7_75t_L g2154 ( 
.A1(n_1967),
.A2(n_2018),
.B1(n_1925),
.B2(n_2017),
.Y(n_2154)
);

OAI211xp5_ASAP7_75t_SL g2155 ( 
.A1(n_1976),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_2155)
);

AOI221xp5_ASAP7_75t_SL g2156 ( 
.A1(n_1944),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.C(n_34),
.Y(n_2156)
);

AOI221xp5_ASAP7_75t_L g2157 ( 
.A1(n_1992),
.A2(n_955),
.B1(n_952),
.B2(n_947),
.C(n_944),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1937),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1939),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1925),
.A2(n_1318),
.B1(n_1311),
.B2(n_944),
.Y(n_2160)
);

OAI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2029),
.A2(n_2031),
.B1(n_2019),
.B2(n_1981),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1939),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1941),
.Y(n_2163)
);

BUFx2_ASAP7_75t_L g2164 ( 
.A(n_1953),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2031),
.B(n_1888),
.Y(n_2165)
);

OAI21x1_ASAP7_75t_L g2166 ( 
.A1(n_2005),
.A2(n_876),
.B(n_850),
.Y(n_2166)
);

OAI211xp5_ASAP7_75t_SL g2167 ( 
.A1(n_2028),
.A2(n_34),
.B(n_31),
.C(n_33),
.Y(n_2167)
);

NAND3xp33_ASAP7_75t_L g2168 ( 
.A(n_2028),
.B(n_947),
.C(n_944),
.Y(n_2168)
);

OAI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2029),
.A2(n_952),
.B1(n_955),
.B2(n_947),
.Y(n_2169)
);

OAI211xp5_ASAP7_75t_SL g2170 ( 
.A1(n_2012),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_1933),
.A2(n_1318),
.B1(n_1210),
.B2(n_1167),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1953),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_1925),
.A2(n_1318),
.B1(n_952),
.B2(n_955),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1953),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1945),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2029),
.A2(n_955),
.B1(n_952),
.B2(n_37),
.Y(n_2176)
);

OAI221xp5_ASAP7_75t_L g2177 ( 
.A1(n_2037),
.A2(n_2013),
.B1(n_2014),
.B2(n_2017),
.C(n_1998),
.Y(n_2177)
);

OAI22xp33_ASAP7_75t_L g2178 ( 
.A1(n_2059),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_1981),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_1928),
.B(n_1929),
.Y(n_2180)
);

OAI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_2059),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1925),
.B(n_1981),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1981),
.A2(n_45),
.B1(n_41),
.B2(n_42),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1945),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_2037),
.A2(n_952),
.B1(n_955),
.B2(n_1147),
.Y(n_2185)
);

O2A1O1Ixp33_ASAP7_75t_SL g2186 ( 
.A1(n_1940),
.A2(n_49),
.B(n_46),
.C(n_48),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2025),
.A2(n_955),
.B1(n_1167),
.B2(n_1210),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_1991),
.B(n_46),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1926),
.B(n_48),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1993),
.A2(n_1167),
.B(n_50),
.Y(n_2190)
);

HB1xp67_ASAP7_75t_L g2191 ( 
.A(n_1996),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_1926),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_1981),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2193)
);

AOI222xp33_ASAP7_75t_L g2194 ( 
.A1(n_2038),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.C1(n_60),
.C2(n_62),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_SL g2195 ( 
.A1(n_2033),
.A2(n_63),
.B1(n_58),
.B2(n_62),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2025),
.A2(n_1266),
.B1(n_1298),
.B2(n_933),
.Y(n_2196)
);

OAI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2013),
.A2(n_64),
.B(n_65),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1982),
.B(n_65),
.Y(n_2198)
);

NAND3xp33_ASAP7_75t_L g2199 ( 
.A(n_2036),
.B(n_66),
.C(n_67),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1941),
.Y(n_2200)
);

AOI22xp33_ASAP7_75t_L g2201 ( 
.A1(n_2025),
.A2(n_1266),
.B1(n_1298),
.B2(n_933),
.Y(n_2201)
);

OAI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_1940),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2060),
.A2(n_2038),
.B1(n_2033),
.B2(n_1991),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2080),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_2180),
.B(n_1996),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2073),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2073),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2062),
.B(n_2061),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2086),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2068),
.B(n_1985),
.Y(n_2210)
);

INVx5_ASAP7_75t_L g2211 ( 
.A(n_2103),
.Y(n_2211)
);

INVx1_ASAP7_75t_SL g2212 ( 
.A(n_2115),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2092),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2108),
.B(n_1991),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2097),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2121),
.B(n_1998),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2086),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_2064),
.A2(n_2033),
.B1(n_1998),
.B2(n_2014),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_L g2219 ( 
.A(n_2117),
.B(n_2036),
.C(n_2012),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2164),
.B(n_1943),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_2091),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2089),
.B(n_1943),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2100),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2163),
.B(n_1986),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2200),
.B(n_1941),
.Y(n_2225)
);

NOR2x1_ASAP7_75t_L g2226 ( 
.A(n_2098),
.B(n_1969),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_2088),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2091),
.Y(n_2228)
);

AND2x6_ASAP7_75t_L g2229 ( 
.A(n_2094),
.B(n_2006),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2082),
.B(n_1974),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2191),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2191),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2192),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2192),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2175),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2179),
.B(n_1969),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2135),
.B(n_1969),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_2182),
.B(n_2032),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2184),
.Y(n_2239)
);

AND2x4_ASAP7_75t_L g2240 ( 
.A(n_2139),
.B(n_2032),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_2139),
.B(n_2034),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2158),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2112),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_2159),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_2075),
.B(n_1979),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_2066),
.A2(n_2040),
.B1(n_2047),
.B2(n_2044),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2141),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2083),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2065),
.B(n_1979),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2067),
.B(n_1979),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2125),
.B(n_1974),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2146),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2150),
.B(n_1949),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2117),
.A2(n_2040),
.B1(n_2047),
.B2(n_2044),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2152),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2162),
.B(n_1949),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2099),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2135),
.B(n_2034),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2111),
.B(n_1975),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2113),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2174),
.B(n_1938),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2078),
.B(n_1957),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2127),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2174),
.B(n_1938),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2172),
.B(n_2128),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2154),
.B(n_2198),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_2109),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2122),
.Y(n_2268)
);

AND2x4_ASAP7_75t_L g2269 ( 
.A(n_2119),
.B(n_1957),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_2107),
.B(n_1962),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_2144),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2081),
.B(n_1962),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_2188),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2153),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2070),
.B(n_1965),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2189),
.B(n_2104),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2153),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2096),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_L g2279 ( 
.A1(n_2102),
.A2(n_2040),
.B1(n_2058),
.B2(n_2055),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2104),
.B(n_2177),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2153),
.B(n_2161),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_2079),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2106),
.B(n_1946),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2165),
.B(n_2123),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2134),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2142),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2165),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2084),
.B(n_2151),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2151),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2137),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2148),
.B(n_1965),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2124),
.Y(n_2292)
);

BUFx2_ASAP7_75t_L g2293 ( 
.A(n_2103),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2103),
.B(n_1975),
.Y(n_2294)
);

OAI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2069),
.A2(n_1973),
.B1(n_1968),
.B2(n_2055),
.Y(n_2295)
);

OAI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_2063),
.A2(n_1973),
.B1(n_1968),
.B2(n_2058),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2090),
.B(n_1946),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2124),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2126),
.A2(n_2143),
.B1(n_2194),
.B2(n_2074),
.Y(n_2299)
);

OAI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2195),
.A2(n_1993),
.B1(n_2006),
.B2(n_1999),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2168),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_2116),
.B(n_69),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2166),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2077),
.B(n_2022),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2072),
.B(n_2022),
.Y(n_2305)
);

OR2x2_ASAP7_75t_L g2306 ( 
.A(n_2149),
.B(n_2023),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2126),
.B(n_2023),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2114),
.B(n_1948),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2199),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2197),
.B(n_1948),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2178),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2195),
.B(n_1956),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2101),
.B(n_1956),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2190),
.B(n_1971),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2176),
.Y(n_2315)
);

INVx2_ASAP7_75t_SL g2316 ( 
.A(n_2120),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_2093),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2156),
.B(n_2024),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2178),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2169),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2147),
.B(n_2024),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2167),
.A2(n_2133),
.B1(n_2131),
.B2(n_2118),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2202),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2255),
.Y(n_2324)
);

BUFx2_ASAP7_75t_L g2325 ( 
.A(n_2226),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_2211),
.B(n_1971),
.Y(n_2326)
);

INVxp67_ASAP7_75t_L g2327 ( 
.A(n_2307),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2299),
.A2(n_2076),
.B1(n_2071),
.B2(n_2181),
.Y(n_2328)
);

INVxp67_ASAP7_75t_L g2329 ( 
.A(n_2307),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2288),
.B(n_1972),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2288),
.B(n_1972),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2204),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2270),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2213),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2313),
.B(n_2181),
.Y(n_2335)
);

NAND2x1_ASAP7_75t_SL g2336 ( 
.A(n_2206),
.B(n_1977),
.Y(n_2336)
);

INVx4_ASAP7_75t_L g2337 ( 
.A(n_2267),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2313),
.B(n_2095),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2215),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2262),
.B(n_2087),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2255),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_2229),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2223),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2243),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2272),
.B(n_2087),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2284),
.B(n_1977),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2208),
.B(n_2251),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2227),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2284),
.B(n_1984),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2248),
.B(n_1984),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2247),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2293),
.B(n_1958),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_2203),
.B(n_2193),
.C(n_2133),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2252),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2209),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2270),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2293),
.B(n_1958),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2235),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2270),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2287),
.B(n_2020),
.Y(n_2360)
);

INVxp67_ASAP7_75t_L g2361 ( 
.A(n_2315),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2211),
.B(n_2020),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2287),
.B(n_2021),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2289),
.B(n_2021),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2235),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2239),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2309),
.B(n_2116),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2289),
.B(n_1964),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2269),
.B(n_1964),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2304),
.B(n_2085),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2269),
.B(n_1966),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2269),
.B(n_1966),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2292),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2239),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2214),
.B(n_2016),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2292),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2214),
.B(n_2016),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2233),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2249),
.B(n_2105),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2250),
.B(n_2157),
.Y(n_2380)
);

OR2x2_ASAP7_75t_L g2381 ( 
.A(n_2230),
.B(n_1936),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2211),
.B(n_2233),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2216),
.B(n_1999),
.Y(n_2383)
);

NAND3xp33_ASAP7_75t_L g2384 ( 
.A(n_2322),
.B(n_2131),
.C(n_2155),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2282),
.B(n_2118),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2234),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_SL g2387 ( 
.A(n_2211),
.B(n_2312),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2216),
.B(n_1988),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2298),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2220),
.B(n_1988),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2276),
.B(n_2183),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2275),
.B(n_2305),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2230),
.B(n_1936),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2220),
.B(n_1990),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2231),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2234),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2237),
.B(n_1990),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2237),
.B(n_1936),
.Y(n_2398)
);

HB1xp67_ASAP7_75t_L g2399 ( 
.A(n_2221),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_2267),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2273),
.B(n_2183),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2253),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2286),
.B(n_1936),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2236),
.B(n_1936),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2236),
.B(n_2002),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2274),
.B(n_2002),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2256),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2205),
.B(n_2004),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2274),
.B(n_2004),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2207),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2231),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2207),
.Y(n_2412)
);

AND2x2_ASAP7_75t_SL g2413 ( 
.A(n_2280),
.B(n_2129),
.Y(n_2413)
);

NAND2x1p5_ASAP7_75t_L g2414 ( 
.A(n_2211),
.B(n_1961),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2274),
.B(n_2238),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2238),
.B(n_2010),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2298),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2238),
.B(n_2010),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2261),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2312),
.B(n_2132),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2217),
.Y(n_2421)
);

AOI221xp5_ASAP7_75t_L g2422 ( 
.A1(n_2311),
.A2(n_2186),
.B1(n_2167),
.B2(n_2155),
.C(n_2170),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2217),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2261),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2228),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2264),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2265),
.B(n_1987),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2265),
.B(n_1987),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2228),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_2232),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2232),
.B(n_2190),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2308),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2264),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_2229),
.Y(n_2434)
);

OR2x2_ASAP7_75t_L g2435 ( 
.A(n_2205),
.B(n_1987),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2281),
.B(n_2001),
.Y(n_2436)
);

BUFx3_ASAP7_75t_L g2437 ( 
.A(n_2400),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2365),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2413),
.B(n_2323),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2413),
.B(n_2323),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2336),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2336),
.Y(n_2442)
);

OAI21x1_ASAP7_75t_L g2443 ( 
.A1(n_2414),
.A2(n_2376),
.B(n_2373),
.Y(n_2443)
);

OA21x2_ASAP7_75t_L g2444 ( 
.A1(n_2327),
.A2(n_2329),
.B(n_2342),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2333),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2365),
.Y(n_2446)
);

OAI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2328),
.A2(n_2384),
.B1(n_2353),
.B2(n_2391),
.C(n_2420),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2387),
.B(n_2278),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2337),
.Y(n_2449)
);

OAI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2392),
.A2(n_2317),
.B1(n_2316),
.B2(n_2218),
.C(n_2319),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2333),
.Y(n_2451)
);

BUFx2_ASAP7_75t_SL g2452 ( 
.A(n_2337),
.Y(n_2452)
);

INVx3_ASAP7_75t_L g2453 ( 
.A(n_2400),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2366),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2361),
.B(n_2291),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2387),
.B(n_2278),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2415),
.B(n_2229),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_2337),
.B(n_2212),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2356),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2415),
.B(n_2229),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2366),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2385),
.A2(n_2317),
.B1(n_2229),
.B2(n_2316),
.Y(n_2462)
);

OAI33xp33_ASAP7_75t_L g2463 ( 
.A1(n_2335),
.A2(n_2318),
.A3(n_2295),
.B1(n_2296),
.B2(n_2300),
.B3(n_2321),
.Y(n_2463)
);

OAI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2347),
.A2(n_2302),
.B1(n_2219),
.B2(n_2266),
.C(n_2245),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2374),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2400),
.B(n_2271),
.Y(n_2466)
);

OAI211xp5_ASAP7_75t_L g2467 ( 
.A1(n_2422),
.A2(n_2246),
.B(n_2254),
.C(n_2279),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2374),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2342),
.B(n_2229),
.Y(n_2469)
);

BUFx3_ASAP7_75t_L g2470 ( 
.A(n_2400),
.Y(n_2470)
);

AO22x1_ASAP7_75t_L g2471 ( 
.A1(n_2340),
.A2(n_2227),
.B1(n_2271),
.B2(n_2301),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2358),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_L g2473 ( 
.A(n_2370),
.B(n_2170),
.C(n_2290),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2356),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2434),
.A2(n_2320),
.B1(n_2210),
.B2(n_2277),
.Y(n_2475)
);

OAI33xp33_ASAP7_75t_L g2476 ( 
.A1(n_2345),
.A2(n_2259),
.A3(n_2306),
.B1(n_2294),
.B2(n_2110),
.B3(n_2263),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2400),
.B(n_2222),
.Y(n_2477)
);

AOI221xp5_ASAP7_75t_L g2478 ( 
.A1(n_2367),
.A2(n_2347),
.B1(n_2338),
.B2(n_2401),
.C(n_2432),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2395),
.Y(n_2479)
);

AOI33xp33_ASAP7_75t_L g2480 ( 
.A1(n_2436),
.A2(n_2310),
.A3(n_2308),
.B1(n_2297),
.B2(n_2130),
.B3(n_2320),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2380),
.B(n_2436),
.C(n_2386),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2395),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2348),
.B(n_2310),
.Y(n_2483)
);

OAI211xp5_ASAP7_75t_L g2484 ( 
.A1(n_2434),
.A2(n_2145),
.B(n_2285),
.C(n_2314),
.Y(n_2484)
);

OAI221xp5_ASAP7_75t_L g2485 ( 
.A1(n_2325),
.A2(n_2294),
.B1(n_2259),
.B2(n_2297),
.C(n_2268),
.Y(n_2485)
);

OAI221xp5_ASAP7_75t_L g2486 ( 
.A1(n_2325),
.A2(n_2268),
.B1(n_2303),
.B2(n_2171),
.C(n_2257),
.Y(n_2486)
);

INVx4_ASAP7_75t_L g2487 ( 
.A(n_2348),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2359),
.Y(n_2488)
);

OAI21xp5_ASAP7_75t_SL g2489 ( 
.A1(n_2379),
.A2(n_2314),
.B(n_2138),
.Y(n_2489)
);

AO21x2_ASAP7_75t_L g2490 ( 
.A1(n_2373),
.A2(n_2241),
.B(n_2240),
.Y(n_2490)
);

OAI33xp33_ASAP7_75t_L g2491 ( 
.A1(n_2378),
.A2(n_2306),
.A3(n_2263),
.B1(n_2242),
.B2(n_2260),
.B3(n_2140),
.Y(n_2491)
);

OR2x6_ASAP7_75t_L g2492 ( 
.A(n_2382),
.B(n_2240),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2359),
.B(n_2240),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_2355),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2376),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_2382),
.Y(n_2496)
);

OA21x2_ASAP7_75t_L g2497 ( 
.A1(n_2389),
.A2(n_2417),
.B(n_2382),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2411),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2330),
.B(n_2241),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2399),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2402),
.B(n_2244),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2389),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2326),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2425),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2417),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2330),
.B(n_2241),
.Y(n_2506)
);

OAI31xp33_ASAP7_75t_SL g2507 ( 
.A1(n_2431),
.A2(n_2224),
.A3(n_2225),
.B(n_2283),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2331),
.B(n_2225),
.Y(n_2508)
);

OAI221xp5_ASAP7_75t_L g2509 ( 
.A1(n_2407),
.A2(n_2260),
.B1(n_2242),
.B2(n_2224),
.C(n_2258),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2396),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2331),
.B(n_2258),
.Y(n_2511)
);

BUFx2_ASAP7_75t_L g2512 ( 
.A(n_2410),
.Y(n_2512)
);

OAI31xp33_ASAP7_75t_L g2513 ( 
.A1(n_2431),
.A2(n_2283),
.A3(n_2160),
.B(n_2173),
.Y(n_2513)
);

OAI31xp33_ASAP7_75t_SL g2514 ( 
.A1(n_2431),
.A2(n_1961),
.A3(n_1959),
.B(n_2046),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2425),
.Y(n_2515)
);

AOI221xp5_ASAP7_75t_SL g2516 ( 
.A1(n_2332),
.A2(n_2187),
.B1(n_2136),
.B2(n_2201),
.C(n_2196),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2412),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2369),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2346),
.B(n_2001),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2429),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2369),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2371),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2346),
.B(n_2001),
.Y(n_2523)
);

OAI33xp33_ASAP7_75t_L g2524 ( 
.A1(n_2421),
.A2(n_2048),
.A3(n_2049),
.B1(n_72),
.B2(n_73),
.B3(n_75),
.Y(n_2524)
);

INVx1_ASAP7_75t_SL g2525 ( 
.A(n_2500),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2458),
.B(n_2349),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2512),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2477),
.B(n_2349),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_2494),
.B(n_2419),
.Y(n_2529)
);

BUFx3_ASAP7_75t_L g2530 ( 
.A(n_2449),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2439),
.B(n_2334),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2462),
.B(n_2478),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_2455),
.B(n_2419),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2512),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2499),
.B(n_2424),
.Y(n_2535)
);

BUFx2_ASAP7_75t_SL g2536 ( 
.A(n_2500),
.Y(n_2536)
);

OR2x2_ASAP7_75t_L g2537 ( 
.A(n_2455),
.B(n_2424),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2499),
.B(n_2426),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2506),
.B(n_2426),
.Y(n_2539)
);

INVx1_ASAP7_75t_SL g2540 ( 
.A(n_2452),
.Y(n_2540)
);

AOI211x1_ASAP7_75t_L g2541 ( 
.A1(n_2467),
.A2(n_2343),
.B(n_2344),
.C(n_2339),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2452),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2506),
.B(n_2433),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2447),
.B(n_2463),
.Y(n_2544)
);

HB1xp67_ASAP7_75t_L g2545 ( 
.A(n_2517),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2440),
.B(n_2351),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_2517),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2520),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2496),
.Y(n_2549)
);

INVx6_ASAP7_75t_L g2550 ( 
.A(n_2487),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2457),
.B(n_2460),
.Y(n_2551)
);

INVx2_ASAP7_75t_SL g2552 ( 
.A(n_2496),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2497),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2520),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2449),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2457),
.B(n_2433),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2460),
.B(n_2493),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2483),
.B(n_2354),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2497),
.Y(n_2559)
);

INVx1_ASAP7_75t_SL g2560 ( 
.A(n_2437),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2487),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2480),
.B(n_2352),
.Y(n_2562)
);

NOR2xp67_ASAP7_75t_L g2563 ( 
.A(n_2496),
.B(n_2430),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_2444),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2471),
.B(n_2487),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2473),
.B(n_2484),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2503),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2471),
.B(n_2352),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2437),
.B(n_2362),
.Y(n_2569)
);

INVx1_ASAP7_75t_SL g2570 ( 
.A(n_2470),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2446),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2470),
.B(n_2357),
.Y(n_2572)
);

OR2x2_ASAP7_75t_L g2573 ( 
.A(n_2501),
.B(n_2423),
.Y(n_2573)
);

OR2x2_ASAP7_75t_L g2574 ( 
.A(n_2481),
.B(n_2444),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2464),
.A2(n_2414),
.B1(n_2326),
.B2(n_2362),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2446),
.Y(n_2576)
);

AOI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2450),
.A2(n_2362),
.B1(n_2357),
.B2(n_2326),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2493),
.B(n_2375),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2461),
.Y(n_2579)
);

OR2x2_ASAP7_75t_L g2580 ( 
.A(n_2444),
.B(n_2489),
.Y(n_2580)
);

INVx4_ASAP7_75t_L g2581 ( 
.A(n_2453),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2475),
.B(n_2324),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2466),
.B(n_2375),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2497),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2453),
.B(n_2513),
.Y(n_2585)
);

NAND5xp2_ASAP7_75t_L g2586 ( 
.A(n_2507),
.B(n_2414),
.C(n_2341),
.D(n_2324),
.E(n_2427),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2453),
.B(n_2427),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2461),
.Y(n_2588)
);

OR2x2_ASAP7_75t_L g2589 ( 
.A(n_2518),
.B(n_2341),
.Y(n_2589)
);

AND2x4_ASAP7_75t_L g2590 ( 
.A(n_2492),
.B(n_2383),
.Y(n_2590)
);

OR2x6_ASAP7_75t_L g2591 ( 
.A(n_2492),
.B(n_2428),
.Y(n_2591)
);

AOI33xp33_ASAP7_75t_L g2592 ( 
.A1(n_2510),
.A2(n_2428),
.A3(n_2404),
.B1(n_2398),
.B2(n_2383),
.B3(n_2406),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2445),
.B(n_2368),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2476),
.B(n_2368),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2465),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2465),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2503),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2479),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2508),
.B(n_2377),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2445),
.B(n_2371),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2503),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2490),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2451),
.B(n_2372),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2508),
.B(n_2511),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2479),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2469),
.B(n_2416),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2527),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2527),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2536),
.B(n_2492),
.Y(n_2609)
);

NOR2x1_ASAP7_75t_SL g2610 ( 
.A(n_2530),
.B(n_2492),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2525),
.B(n_2469),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2545),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2551),
.B(n_2448),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2560),
.B(n_2451),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2570),
.B(n_2459),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2557),
.B(n_2606),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2544),
.B(n_2459),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2584),
.Y(n_2618)
);

INVx1_ASAP7_75t_SL g2619 ( 
.A(n_2540),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2529),
.B(n_2518),
.Y(n_2620)
);

OR2x2_ASAP7_75t_L g2621 ( 
.A(n_2533),
.B(n_2537),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2544),
.B(n_2474),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2606),
.B(n_2448),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2545),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2526),
.B(n_2456),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2584),
.Y(n_2626)
);

NAND2x1p5_ASAP7_75t_L g2627 ( 
.A(n_2542),
.B(n_2530),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2547),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2547),
.Y(n_2629)
);

INVx1_ASAP7_75t_SL g2630 ( 
.A(n_2550),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2604),
.B(n_2456),
.Y(n_2631)
);

OR2x2_ASAP7_75t_L g2632 ( 
.A(n_2562),
.B(n_2521),
.Y(n_2632)
);

OR2x2_ASAP7_75t_L g2633 ( 
.A(n_2580),
.B(n_2521),
.Y(n_2633)
);

NAND2x1p5_ASAP7_75t_L g2634 ( 
.A(n_2555),
.B(n_2443),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2564),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2594),
.B(n_2474),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2594),
.B(n_2488),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2566),
.B(n_2488),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2564),
.Y(n_2639)
);

HB1xp67_ASAP7_75t_L g2640 ( 
.A(n_2563),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2555),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2531),
.B(n_2522),
.Y(n_2642)
);

NAND2x1p5_ASAP7_75t_L g2643 ( 
.A(n_2561),
.B(n_2443),
.Y(n_2643)
);

OR2x2_ASAP7_75t_L g2644 ( 
.A(n_2546),
.B(n_2522),
.Y(n_2644)
);

AND2x2_ASAP7_75t_SL g2645 ( 
.A(n_2574),
.B(n_2441),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2566),
.B(n_2472),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2528),
.B(n_2511),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2583),
.B(n_2441),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2534),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2548),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2554),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2541),
.B(n_2532),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2571),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2532),
.A2(n_2491),
.B1(n_2524),
.B2(n_2486),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2597),
.B(n_2495),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2585),
.B(n_2498),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2561),
.B(n_2498),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2576),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2561),
.B(n_2438),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2550),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2579),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2569),
.B(n_2442),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2569),
.B(n_2442),
.Y(n_2663)
);

OR2x2_ASAP7_75t_L g2664 ( 
.A(n_2568),
.B(n_2509),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2569),
.B(n_2495),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2556),
.B(n_2502),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2572),
.B(n_2485),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2578),
.B(n_2502),
.Y(n_2668)
);

OAI32xp33_ASAP7_75t_L g2669 ( 
.A1(n_2652),
.A2(n_2565),
.A3(n_2582),
.B1(n_2575),
.B2(n_2553),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_L g2670 ( 
.A(n_2619),
.B(n_2550),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2616),
.B(n_2613),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2616),
.B(n_2535),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2641),
.Y(n_2673)
);

INVxp67_ASAP7_75t_SL g2674 ( 
.A(n_2627),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_SL g2675 ( 
.A1(n_2645),
.A2(n_2586),
.B1(n_2590),
.B2(n_2552),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2641),
.Y(n_2676)
);

NAND3xp33_ASAP7_75t_SL g2677 ( 
.A(n_2654),
.B(n_2577),
.C(n_2575),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2607),
.B(n_2549),
.Y(n_2678)
);

OR2x2_ASAP7_75t_L g2679 ( 
.A(n_2614),
.B(n_2558),
.Y(n_2679)
);

OAI32xp33_ASAP7_75t_L g2680 ( 
.A1(n_2636),
.A2(n_2553),
.A3(n_2559),
.B1(n_2581),
.B2(n_2573),
.Y(n_2680)
);

AOI21xp33_ASAP7_75t_SL g2681 ( 
.A1(n_2627),
.A2(n_2552),
.B(n_2549),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2618),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2618),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2626),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2626),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2608),
.B(n_2588),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2612),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2624),
.B(n_2595),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2613),
.B(n_2538),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2628),
.Y(n_2690)
);

OR2x2_ASAP7_75t_L g2691 ( 
.A(n_2615),
.B(n_2621),
.Y(n_2691)
);

OAI21xp33_ASAP7_75t_SL g2692 ( 
.A1(n_2645),
.A2(n_2592),
.B(n_2567),
.Y(n_2692)
);

AOI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2637),
.A2(n_2567),
.B(n_2559),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2629),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2635),
.Y(n_2695)
);

OR2x2_ASAP7_75t_L g2696 ( 
.A(n_2633),
.B(n_2600),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2611),
.B(n_2539),
.Y(n_2697)
);

OAI33xp33_ASAP7_75t_L g2698 ( 
.A1(n_2617),
.A2(n_2605),
.A3(n_2596),
.B1(n_2598),
.B2(n_2601),
.B3(n_2597),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2611),
.B(n_2601),
.Y(n_2699)
);

NAND4xp25_ASAP7_75t_L g2700 ( 
.A(n_2609),
.B(n_2581),
.C(n_2592),
.D(n_2587),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2639),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2640),
.Y(n_2702)
);

INVxp67_ASAP7_75t_SL g2703 ( 
.A(n_2640),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2622),
.B(n_2581),
.Y(n_2704)
);

NAND3xp33_ASAP7_75t_L g2705 ( 
.A(n_2646),
.B(n_2603),
.C(n_2602),
.Y(n_2705)
);

HB1xp67_ASAP7_75t_L g2706 ( 
.A(n_2623),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2655),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2649),
.B(n_2454),
.Y(n_2708)
);

OAI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2664),
.A2(n_2656),
.B(n_2609),
.Y(n_2709)
);

NAND2x1p5_ASAP7_75t_L g2710 ( 
.A(n_2630),
.B(n_2590),
.Y(n_2710)
);

O2A1O1Ixp5_ASAP7_75t_L g2711 ( 
.A1(n_2638),
.A2(n_2590),
.B(n_2602),
.C(n_2593),
.Y(n_2711)
);

INVx2_ASAP7_75t_SL g2712 ( 
.A(n_2665),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2610),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2650),
.B(n_2468),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2665),
.Y(n_2715)
);

OAI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2675),
.A2(n_2667),
.B1(n_2632),
.B2(n_2631),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2710),
.Y(n_2717)
);

O2A1O1Ixp5_ASAP7_75t_L g2718 ( 
.A1(n_2669),
.A2(n_2660),
.B(n_2651),
.C(n_2659),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2706),
.Y(n_2719)
);

OAI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2692),
.A2(n_2634),
.B(n_2648),
.Y(n_2720)
);

NAND4xp25_ASAP7_75t_L g2721 ( 
.A(n_2709),
.B(n_2660),
.C(n_2657),
.D(n_2658),
.Y(n_2721)
);

AOI22xp5_ASAP7_75t_L g2722 ( 
.A1(n_2677),
.A2(n_2631),
.B1(n_2625),
.B2(n_2623),
.Y(n_2722)
);

OAI32xp33_ASAP7_75t_L g2723 ( 
.A1(n_2710),
.A2(n_2634),
.A3(n_2643),
.B1(n_2620),
.B2(n_2642),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2671),
.B(n_2648),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2713),
.B(n_2625),
.Y(n_2725)
);

NAND2x1_ASAP7_75t_L g2726 ( 
.A(n_2715),
.B(n_2662),
.Y(n_2726)
);

AOI221xp5_ASAP7_75t_L g2727 ( 
.A1(n_2680),
.A2(n_2681),
.B1(n_2693),
.B2(n_2711),
.C(n_2674),
.Y(n_2727)
);

OR2x2_ASAP7_75t_L g2728 ( 
.A(n_2699),
.B(n_2644),
.Y(n_2728)
);

CKINVDCx14_ASAP7_75t_R g2729 ( 
.A(n_2670),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2702),
.Y(n_2730)
);

INVxp67_ASAP7_75t_L g2731 ( 
.A(n_2703),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_R g2732 ( 
.A(n_2673),
.B(n_2653),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2704),
.A2(n_2666),
.B(n_2663),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2697),
.A2(n_2647),
.B1(n_2543),
.B2(n_2668),
.Y(n_2734)
);

OAI321xp33_ASAP7_75t_L g2735 ( 
.A1(n_2700),
.A2(n_2643),
.A3(n_2663),
.B1(n_2662),
.B2(n_2666),
.C(n_2591),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2676),
.Y(n_2736)
);

OAI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2691),
.A2(n_2591),
.B1(n_2655),
.B2(n_2589),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2699),
.Y(n_2738)
);

AOI22xp33_ASAP7_75t_L g2739 ( 
.A1(n_2672),
.A2(n_2647),
.B1(n_2668),
.B2(n_2591),
.Y(n_2739)
);

NAND4xp25_ASAP7_75t_SL g2740 ( 
.A(n_2704),
.B(n_2689),
.C(n_2705),
.D(n_2678),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2715),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2712),
.B(n_2599),
.Y(n_2742)
);

OAI221xp5_ASAP7_75t_L g2743 ( 
.A1(n_2696),
.A2(n_2661),
.B1(n_2514),
.B2(n_2482),
.C(n_2515),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2687),
.B(n_2482),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_2682),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2683),
.Y(n_2746)
);

OAI32xp33_ASAP7_75t_L g2747 ( 
.A1(n_2679),
.A2(n_2515),
.A3(n_2504),
.B1(n_2505),
.B2(n_2393),
.Y(n_2747)
);

OAI211xp5_ASAP7_75t_SL g2748 ( 
.A1(n_2678),
.A2(n_2505),
.B(n_2504),
.C(n_2381),
.Y(n_2748)
);

AOI221xp5_ASAP7_75t_L g2749 ( 
.A1(n_2698),
.A2(n_2490),
.B1(n_2516),
.B2(n_2519),
.C(n_2523),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2684),
.Y(n_2750)
);

INVxp67_ASAP7_75t_SL g2751 ( 
.A(n_2707),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_SL g2752 ( 
.A1(n_2685),
.A2(n_2523),
.B(n_2519),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2695),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2726),
.Y(n_2754)
);

AOI32xp33_ASAP7_75t_L g2755 ( 
.A1(n_2727),
.A2(n_2735),
.A3(n_2716),
.B1(n_2748),
.B2(n_2742),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2745),
.Y(n_2756)
);

AOI222xp33_ASAP7_75t_L g2757 ( 
.A1(n_2731),
.A2(n_2694),
.B1(n_2690),
.B2(n_2701),
.C1(n_2686),
.C2(n_2688),
.Y(n_2757)
);

OAI322xp33_ASAP7_75t_L g2758 ( 
.A1(n_2722),
.A2(n_2688),
.A3(n_2686),
.B1(n_2714),
.B2(n_2708),
.C1(n_2381),
.C2(n_2393),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2729),
.B(n_2708),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2734),
.B(n_2714),
.Y(n_2760)
);

AOI32xp33_ASAP7_75t_L g2761 ( 
.A1(n_2737),
.A2(n_2416),
.A3(n_2418),
.B1(n_2404),
.B2(n_2398),
.Y(n_2761)
);

INVxp67_ASAP7_75t_L g2762 ( 
.A(n_2724),
.Y(n_2762)
);

NAND3xp33_ASAP7_75t_L g2763 ( 
.A(n_2720),
.B(n_2403),
.C(n_2406),
.Y(n_2763)
);

AOI21xp33_ASAP7_75t_SL g2764 ( 
.A1(n_2717),
.A2(n_2490),
.B(n_70),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2745),
.Y(n_2765)
);

AOI322xp5_ASAP7_75t_L g2766 ( 
.A1(n_2751),
.A2(n_2418),
.A3(n_2388),
.B1(n_2409),
.B2(n_2390),
.C1(n_2394),
.C2(n_2405),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2721),
.B(n_2408),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2745),
.Y(n_2768)
);

OAI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2721),
.A2(n_2403),
.B1(n_2435),
.B2(n_2408),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2741),
.Y(n_2770)
);

OAI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2743),
.A2(n_2435),
.B1(n_2409),
.B2(n_2388),
.Y(n_2771)
);

INVxp67_ASAP7_75t_L g2772 ( 
.A(n_2725),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2730),
.Y(n_2773)
);

OAI32xp33_ASAP7_75t_L g2774 ( 
.A1(n_2719),
.A2(n_2394),
.A3(n_2390),
.B1(n_2405),
.B2(n_2397),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2733),
.B(n_2372),
.Y(n_2775)
);

AO21x1_ASAP7_75t_L g2776 ( 
.A1(n_2746),
.A2(n_2363),
.B(n_2360),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2736),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2728),
.Y(n_2778)
);

OAI221xp5_ASAP7_75t_SL g2779 ( 
.A1(n_2749),
.A2(n_2397),
.B1(n_2350),
.B2(n_2377),
.C(n_2363),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2750),
.Y(n_2780)
);

OAI222xp33_ASAP7_75t_L g2781 ( 
.A1(n_2739),
.A2(n_2350),
.B1(n_2360),
.B2(n_2364),
.C1(n_2043),
.C2(n_2185),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2740),
.B(n_2364),
.Y(n_2782)
);

OAI322xp33_ASAP7_75t_L g2783 ( 
.A1(n_2738),
.A2(n_71),
.A3(n_73),
.B1(n_76),
.B2(n_78),
.C1(n_79),
.C2(n_81),
.Y(n_2783)
);

AOI21xp33_ASAP7_75t_L g2784 ( 
.A1(n_2723),
.A2(n_79),
.B(n_81),
.Y(n_2784)
);

OAI22xp33_ASAP7_75t_SL g2785 ( 
.A1(n_2753),
.A2(n_2043),
.B1(n_89),
.B2(n_86),
.Y(n_2785)
);

OAI221xp5_ASAP7_75t_SL g2786 ( 
.A1(n_2755),
.A2(n_2744),
.B1(n_2752),
.B2(n_2718),
.C(n_2732),
.Y(n_2786)
);

AOI221xp5_ASAP7_75t_L g2787 ( 
.A1(n_2784),
.A2(n_2747),
.B1(n_2752),
.B2(n_91),
.C(n_92),
.Y(n_2787)
);

NOR2x1_ASAP7_75t_L g2788 ( 
.A(n_2759),
.B(n_2756),
.Y(n_2788)
);

NOR2xp67_ASAP7_75t_L g2789 ( 
.A(n_2754),
.B(n_88),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2784),
.A2(n_1959),
.B(n_90),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2765),
.Y(n_2791)
);

AOI222xp33_ASAP7_75t_L g2792 ( 
.A1(n_2772),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.C1(n_97),
.C2(n_99),
.Y(n_2792)
);

AOI221xp5_ASAP7_75t_L g2793 ( 
.A1(n_2758),
.A2(n_2779),
.B1(n_2764),
.B2(n_2782),
.C(n_2771),
.Y(n_2793)
);

AOI222xp33_ASAP7_75t_L g2794 ( 
.A1(n_2760),
.A2(n_93),
.B1(n_94),
.B2(n_99),
.C1(n_100),
.C2(n_101),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2768),
.B(n_101),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2757),
.B(n_102),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2778),
.A2(n_103),
.B(n_104),
.Y(n_2797)
);

OAI221xp5_ASAP7_75t_L g2798 ( 
.A1(n_2761),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.C(n_107),
.Y(n_2798)
);

AOI211xp5_ASAP7_75t_L g2799 ( 
.A1(n_2770),
.A2(n_2773),
.B(n_2762),
.C(n_2783),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_L g2800 ( 
.A(n_2767),
.B(n_105),
.Y(n_2800)
);

AOI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2775),
.A2(n_2049),
.B1(n_2048),
.B2(n_2046),
.Y(n_2801)
);

OAI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2763),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2757),
.B(n_110),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_SL g2804 ( 
.A1(n_2785),
.A2(n_111),
.B(n_112),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2777),
.B(n_111),
.Y(n_2805)
);

AND3x1_ASAP7_75t_L g2806 ( 
.A(n_2780),
.B(n_2781),
.C(n_2776),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2769),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_2807)
);

OAI322xp33_ASAP7_75t_L g2808 ( 
.A1(n_2774),
.A2(n_113),
.A3(n_114),
.B1(n_116),
.B2(n_117),
.C1(n_118),
.C2(n_120),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2766),
.B(n_116),
.Y(n_2809)
);

A2O1A1Ixp33_ASAP7_75t_L g2810 ( 
.A1(n_2755),
.A2(n_117),
.B(n_118),
.C(n_120),
.Y(n_2810)
);

AOI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2786),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.C(n_124),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2789),
.Y(n_2812)
);

O2A1O1Ixp5_ASAP7_75t_L g2813 ( 
.A1(n_2796),
.A2(n_121),
.B(n_122),
.C(n_126),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_SL g2814 ( 
.A1(n_2803),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_2814)
);

AOI221xp5_ASAP7_75t_L g2815 ( 
.A1(n_2810),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_2815)
);

AOI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2793),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_2816)
);

AOI221xp5_ASAP7_75t_L g2817 ( 
.A1(n_2806),
.A2(n_2787),
.B1(n_2802),
.B2(n_2807),
.C(n_2800),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2788),
.Y(n_2818)
);

OAI21xp5_ASAP7_75t_SL g2819 ( 
.A1(n_2798),
.A2(n_131),
.B(n_132),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2809),
.A2(n_2791),
.B1(n_2799),
.B2(n_2805),
.Y(n_2820)
);

AOI221x1_ASAP7_75t_L g2821 ( 
.A1(n_2797),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.C(n_137),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2795),
.Y(n_2822)
);

OAI211xp5_ASAP7_75t_SL g2823 ( 
.A1(n_2804),
.A2(n_135),
.B(n_137),
.C(n_138),
.Y(n_2823)
);

AOI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2794),
.A2(n_2792),
.B1(n_2790),
.B2(n_2801),
.Y(n_2824)
);

INVxp67_ASAP7_75t_L g2825 ( 
.A(n_2808),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2789),
.Y(n_2826)
);

BUFx6f_ASAP7_75t_L g2827 ( 
.A(n_2791),
.Y(n_2827)
);

AOI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2796),
.A2(n_138),
.B(n_140),
.Y(n_2828)
);

AOI221x1_ASAP7_75t_L g2829 ( 
.A1(n_2810),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.C(n_146),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2812),
.Y(n_2830)
);

OAI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2816),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2826),
.Y(n_2832)
);

OAI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2825),
.A2(n_147),
.B(n_148),
.Y(n_2833)
);

AOI21xp33_ASAP7_75t_L g2834 ( 
.A1(n_2818),
.A2(n_2820),
.B(n_2822),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2814),
.B(n_147),
.Y(n_2835)
);

OAI21xp33_ASAP7_75t_L g2836 ( 
.A1(n_2811),
.A2(n_150),
.B(n_151),
.Y(n_2836)
);

OAI32xp33_ASAP7_75t_L g2837 ( 
.A1(n_2823),
.A2(n_150),
.A3(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_2837)
);

OAI21x1_ASAP7_75t_L g2838 ( 
.A1(n_2813),
.A2(n_152),
.B(n_156),
.Y(n_2838)
);

OAI321xp33_ASAP7_75t_L g2839 ( 
.A1(n_2817),
.A2(n_156),
.A3(n_158),
.B1(n_159),
.B2(n_160),
.C(n_161),
.Y(n_2839)
);

AOI22x1_ASAP7_75t_L g2840 ( 
.A1(n_2827),
.A2(n_2828),
.B1(n_2829),
.B2(n_2821),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2827),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2827),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_2842)
);

AOI31xp33_ASAP7_75t_L g2843 ( 
.A1(n_2834),
.A2(n_2841),
.A3(n_2830),
.B(n_2832),
.Y(n_2843)
);

INVxp67_ASAP7_75t_L g2844 ( 
.A(n_2840),
.Y(n_2844)
);

NOR4xp25_ASAP7_75t_L g2845 ( 
.A(n_2836),
.B(n_2819),
.C(n_2815),
.D(n_2824),
.Y(n_2845)
);

AOI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2839),
.A2(n_162),
.B(n_163),
.Y(n_2846)
);

XNOR2x1_ASAP7_75t_L g2847 ( 
.A(n_2833),
.B(n_163),
.Y(n_2847)
);

OAI21xp33_ASAP7_75t_SL g2848 ( 
.A1(n_2838),
.A2(n_166),
.B(n_168),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2835),
.Y(n_2849)
);

AOI321xp33_ASAP7_75t_L g2850 ( 
.A1(n_2837),
.A2(n_166),
.A3(n_169),
.B1(n_172),
.B2(n_173),
.C(n_174),
.Y(n_2850)
);

NAND2x1p5_ASAP7_75t_L g2851 ( 
.A(n_2839),
.B(n_173),
.Y(n_2851)
);

NAND5xp2_ASAP7_75t_L g2852 ( 
.A(n_2842),
.B(n_175),
.C(n_176),
.D(n_177),
.E(n_179),
.Y(n_2852)
);

XOR2xp5_ASAP7_75t_L g2853 ( 
.A(n_2831),
.B(n_175),
.Y(n_2853)
);

A2O1A1Ixp33_ASAP7_75t_L g2854 ( 
.A1(n_2839),
.A2(n_179),
.B(n_181),
.C(n_182),
.Y(n_2854)
);

XNOR2xp5_ASAP7_75t_L g2855 ( 
.A(n_2840),
.B(n_182),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2855),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2851),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2844),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2853),
.Y(n_2859)
);

NOR2xp67_ASAP7_75t_L g2860 ( 
.A(n_2848),
.B(n_184),
.Y(n_2860)
);

AOI221xp5_ASAP7_75t_L g2861 ( 
.A1(n_2843),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.C(n_190),
.Y(n_2861)
);

NOR2x1_ASAP7_75t_L g2862 ( 
.A(n_2846),
.B(n_187),
.Y(n_2862)
);

NOR2x1_ASAP7_75t_L g2863 ( 
.A(n_2854),
.B(n_2847),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2850),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2845),
.B(n_191),
.Y(n_2865)
);

NOR2x1_ASAP7_75t_L g2866 ( 
.A(n_2852),
.B(n_191),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2849),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2844),
.A2(n_192),
.B1(n_194),
.B2(n_197),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2855),
.Y(n_2869)
);

NOR2x1_ASAP7_75t_L g2870 ( 
.A(n_2855),
.B(n_192),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2851),
.Y(n_2871)
);

OR2x2_ASAP7_75t_L g2872 ( 
.A(n_2851),
.B(n_198),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2872),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_SL g2874 ( 
.A(n_2857),
.B(n_198),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2871),
.Y(n_2875)
);

OR2x2_ASAP7_75t_L g2876 ( 
.A(n_2865),
.B(n_199),
.Y(n_2876)
);

AOI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2864),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_2877)
);

AO22x2_ASAP7_75t_L g2878 ( 
.A1(n_2856),
.A2(n_2869),
.B1(n_2867),
.B2(n_2859),
.Y(n_2878)
);

NOR2x1_ASAP7_75t_L g2879 ( 
.A(n_2870),
.B(n_203),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2866),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_2880)
);

AOI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2863),
.A2(n_204),
.B1(n_207),
.B2(n_209),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2860),
.B(n_2858),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2862),
.Y(n_2883)
);

NOR2x1p5_ASAP7_75t_L g2884 ( 
.A(n_2861),
.B(n_209),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2868),
.Y(n_2885)
);

NAND4xp75_ASAP7_75t_L g2886 ( 
.A(n_2870),
.B(n_211),
.C(n_213),
.D(n_216),
.Y(n_2886)
);

INVxp33_ASAP7_75t_L g2887 ( 
.A(n_2866),
.Y(n_2887)
);

OAI21xp5_ASAP7_75t_SL g2888 ( 
.A1(n_2880),
.A2(n_211),
.B(n_217),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2879),
.Y(n_2889)
);

AOI22xp5_ASAP7_75t_L g2890 ( 
.A1(n_2875),
.A2(n_1298),
.B1(n_1266),
.B2(n_893),
.Y(n_2890)
);

NAND3xp33_ASAP7_75t_SL g2891 ( 
.A(n_2874),
.B(n_222),
.C(n_225),
.Y(n_2891)
);

AOI221xp5_ASAP7_75t_L g2892 ( 
.A1(n_2887),
.A2(n_876),
.B1(n_850),
.B2(n_230),
.C(n_231),
.Y(n_2892)
);

AOI211xp5_ASAP7_75t_L g2893 ( 
.A1(n_2883),
.A2(n_228),
.B(n_229),
.C(n_233),
.Y(n_2893)
);

AOI221xp5_ASAP7_75t_L g2894 ( 
.A1(n_2878),
.A2(n_876),
.B1(n_850),
.B2(n_237),
.C(n_238),
.Y(n_2894)
);

OAI211xp5_ASAP7_75t_L g2895 ( 
.A1(n_2882),
.A2(n_235),
.B(n_236),
.C(n_239),
.Y(n_2895)
);

OAI211xp5_ASAP7_75t_L g2896 ( 
.A1(n_2881),
.A2(n_240),
.B(n_243),
.C(n_244),
.Y(n_2896)
);

OAI22x1_ASAP7_75t_L g2897 ( 
.A1(n_2877),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_2897)
);

AOI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_2878),
.A2(n_899),
.B(n_896),
.Y(n_2898)
);

AOI221xp5_ASAP7_75t_L g2899 ( 
.A1(n_2873),
.A2(n_258),
.B1(n_259),
.B2(n_265),
.C(n_266),
.Y(n_2899)
);

XNOR2xp5_ASAP7_75t_L g2900 ( 
.A(n_2889),
.B(n_2884),
.Y(n_2900)
);

INVx3_ASAP7_75t_L g2901 ( 
.A(n_2891),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2888),
.B(n_2886),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2898),
.B(n_2885),
.Y(n_2903)
);

AOI21xp5_ASAP7_75t_L g2904 ( 
.A1(n_2897),
.A2(n_2876),
.B(n_896),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2895),
.Y(n_2905)
);

XNOR2xp5_ASAP7_75t_L g2906 ( 
.A(n_2896),
.B(n_267),
.Y(n_2906)
);

BUFx3_ASAP7_75t_L g2907 ( 
.A(n_2893),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2894),
.B(n_271),
.Y(n_2908)
);

AND2x4_ASAP7_75t_L g2909 ( 
.A(n_2890),
.B(n_278),
.Y(n_2909)
);

XNOR2x1_ASAP7_75t_L g2910 ( 
.A(n_2892),
.B(n_279),
.Y(n_2910)
);

NAND2x1p5_ASAP7_75t_L g2911 ( 
.A(n_2901),
.B(n_2899),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2900),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2904),
.B(n_283),
.Y(n_2913)
);

XNOR2xp5_ASAP7_75t_L g2914 ( 
.A(n_2900),
.B(n_285),
.Y(n_2914)
);

AOI22xp33_ASAP7_75t_L g2915 ( 
.A1(n_2907),
.A2(n_1298),
.B1(n_1266),
.B2(n_893),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2902),
.A2(n_896),
.B(n_899),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2906),
.Y(n_2917)
);

XOR2xp5_ASAP7_75t_L g2918 ( 
.A(n_2910),
.B(n_287),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2905),
.B(n_289),
.Y(n_2919)
);

AOI31xp33_ASAP7_75t_L g2920 ( 
.A1(n_2903),
.A2(n_290),
.A3(n_292),
.B(n_295),
.Y(n_2920)
);

XNOR2xp5_ASAP7_75t_L g2921 ( 
.A(n_2909),
.B(n_298),
.Y(n_2921)
);

NOR2x1_ASAP7_75t_L g2922 ( 
.A(n_2908),
.B(n_301),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2914),
.Y(n_2923)
);

AOI22xp33_ASAP7_75t_L g2924 ( 
.A1(n_2912),
.A2(n_1298),
.B1(n_1266),
.B2(n_893),
.Y(n_2924)
);

NAND2x1p5_ASAP7_75t_L g2925 ( 
.A(n_2922),
.B(n_899),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2921),
.Y(n_2926)
);

BUFx2_ASAP7_75t_L g2927 ( 
.A(n_2911),
.Y(n_2927)
);

XOR2xp5_ASAP7_75t_L g2928 ( 
.A(n_2918),
.B(n_302),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2920),
.B(n_303),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2928),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2927),
.Y(n_2931)
);

NOR2xp67_ASAP7_75t_L g2932 ( 
.A(n_2929),
.B(n_2919),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2925),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2923),
.Y(n_2934)
);

INVxp33_ASAP7_75t_SL g2935 ( 
.A(n_2926),
.Y(n_2935)
);

OAI22xp5_ASAP7_75t_SL g2936 ( 
.A1(n_2924),
.A2(n_2917),
.B1(n_2913),
.B2(n_2916),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2927),
.A2(n_2915),
.B1(n_893),
.B2(n_914),
.Y(n_2937)
);

XNOR2xp5_ASAP7_75t_L g2938 ( 
.A(n_2928),
.B(n_304),
.Y(n_2938)
);

XOR2xp5_ASAP7_75t_L g2939 ( 
.A(n_2928),
.B(n_305),
.Y(n_2939)
);

AOI22x1_ASAP7_75t_L g2940 ( 
.A1(n_2927),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_SL g2941 ( 
.A1(n_2931),
.A2(n_314),
.B1(n_315),
.B2(n_317),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_SL g2942 ( 
.A1(n_2939),
.A2(n_326),
.B1(n_341),
.B2(n_348),
.Y(n_2942)
);

AOI22x1_ASAP7_75t_L g2943 ( 
.A1(n_2938),
.A2(n_351),
.B1(n_353),
.B2(n_356),
.Y(n_2943)
);

HB1xp67_ASAP7_75t_L g2944 ( 
.A(n_2932),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2940),
.Y(n_2945)
);

OAI22xp5_ASAP7_75t_L g2946 ( 
.A1(n_2935),
.A2(n_899),
.B1(n_896),
.B2(n_359),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2945),
.A2(n_2934),
.B1(n_2930),
.B2(n_2936),
.Y(n_2947)
);

OAI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2944),
.A2(n_2937),
.B(n_2933),
.Y(n_2948)
);

AOI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2942),
.A2(n_914),
.B1(n_893),
.B2(n_869),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2943),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2946),
.A2(n_899),
.B(n_896),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2941),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2947),
.A2(n_899),
.B(n_896),
.Y(n_2953)
);

AOI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2952),
.A2(n_931),
.B(n_897),
.Y(n_2954)
);

AOI21xp33_ASAP7_75t_SL g2955 ( 
.A1(n_2950),
.A2(n_357),
.B(n_358),
.Y(n_2955)
);

INVxp67_ASAP7_75t_SL g2956 ( 
.A(n_2949),
.Y(n_2956)
);

AOI222xp33_ASAP7_75t_L g2957 ( 
.A1(n_2956),
.A2(n_2948),
.B1(n_2951),
.B2(n_914),
.C1(n_893),
.C2(n_366),
.Y(n_2957)
);

OAI221xp5_ASAP7_75t_L g2958 ( 
.A1(n_2955),
.A2(n_360),
.B1(n_361),
.B2(n_364),
.C(n_365),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2958),
.A2(n_2954),
.B1(n_2953),
.B2(n_914),
.Y(n_2959)
);

OA21x2_ASAP7_75t_L g2960 ( 
.A1(n_2959),
.A2(n_2957),
.B(n_372),
.Y(n_2960)
);

AOI221xp5_ASAP7_75t_L g2961 ( 
.A1(n_2960),
.A2(n_869),
.B1(n_864),
.B2(n_894),
.C(n_931),
.Y(n_2961)
);

AOI211xp5_ASAP7_75t_L g2962 ( 
.A1(n_2961),
.A2(n_869),
.B(n_864),
.C(n_375),
.Y(n_2962)
);


endmodule