module fake_ariane_1955_n_2095 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2095);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2095;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_209),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_48),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_40),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx6p67_ASAP7_75t_R g222 ( 
.A(n_50),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_25),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_0),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_11),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_183),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_39),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_190),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_78),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_148),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_98),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_156),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_105),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_114),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_200),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_45),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_7),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_120),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_37),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_169),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_119),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_199),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_59),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_94),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_37),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_159),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_24),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_113),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_54),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_152),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_57),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_49),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_103),
.Y(n_269)
);

BUFx8_ASAP7_75t_SL g270 ( 
.A(n_93),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_116),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_86),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_67),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_147),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_28),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_206),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_33),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_17),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_100),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_110),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_160),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_212),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_163),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_81),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_158),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_91),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_43),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_168),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_41),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_15),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_185),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_19),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_144),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_9),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_96),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_155),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_28),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_22),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_194),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_22),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_71),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_64),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_112),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_157),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_64),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_79),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_65),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_31),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_138),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_24),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_77),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_49),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_27),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_83),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_67),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_65),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_63),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_26),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_184),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_117),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_56),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_181),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_23),
.Y(n_333)
);

BUFx8_ASAP7_75t_SL g334 ( 
.A(n_76),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_45),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_201),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_101),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_124),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_189),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_31),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_85),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_123),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_48),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_125),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_12),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_205),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_102),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_18),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_3),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_80),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_75),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_211),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_130),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_44),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_18),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_139),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_207),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_38),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_29),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_26),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_131),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_59),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_29),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_38),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_115),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_63),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_191),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_127),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_137),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_87),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_97),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_145),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_13),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_70),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_171),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_134),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_53),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_23),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_2),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_172),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_198),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_58),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_25),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_55),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_151),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_153),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_99),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_142),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_1),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_33),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_75),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_58),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_17),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_140),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_11),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_30),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_36),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_44),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_121),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_68),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_135),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_106),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_162),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_71),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_32),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_54),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_2),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_72),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_35),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_88),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_90),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_40),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_69),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_72),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_141),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_173),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_208),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_133),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_334),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_219),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_270),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_321),
.Y(n_425)
);

BUFx6f_ASAP7_75t_SL g426 ( 
.A(n_363),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_222),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_219),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_219),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_219),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_222),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_243),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_220),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_219),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_353),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_220),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_391),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_224),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_343),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_R g442 ( 
.A(n_257),
.B(n_82),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_226),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_224),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_309),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_224),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_224),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_256),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_262),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_224),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_266),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_247),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_268),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_249),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_317),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_247),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_343),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_275),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_247),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_R g460 ( 
.A(n_338),
.B(n_84),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_293),
.Y(n_461)
);

BUFx2_ASAP7_75t_SL g462 ( 
.A(n_363),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_294),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_285),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_247),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_322),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_285),
.B(n_1),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_346),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_247),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_295),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_R g472 ( 
.A(n_213),
.B(n_136),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_377),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_420),
.B(n_4),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_215),
.B(n_4),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_223),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_297),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_299),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_230),
.B(n_5),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_362),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_259),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_377),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_306),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_235),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_392),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_307),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_235),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_291),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_259),
.B(n_5),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_291),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_221),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_363),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_221),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_378),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_378),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_378),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_310),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_227),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_272),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_271),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_271),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_248),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_311),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_264),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_267),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_272),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_259),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_276),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_251),
.B(n_6),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_278),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_280),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_281),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_314),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_409),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_409),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_409),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_411),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_302),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_411),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_304),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_316),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_226),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_323),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_325),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_411),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_326),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_320),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_327),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_454),
.B(n_213),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_379),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_445),
.B(n_233),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_448),
.B(n_449),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_341),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_462),
.B(n_426),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_430),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_431),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_491),
.B(n_381),
.C(n_355),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_451),
.B(n_214),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_441),
.B(n_417),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_501),
.B(n_341),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_440),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_444),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_501),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_446),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_457),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_480),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_459),
.B(n_274),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_493),
.B(n_288),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_296),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_447),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_447),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_455),
.B(n_233),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_435),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_474),
.A2(n_395),
.B1(n_399),
.B2(n_416),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_495),
.B(n_301),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_458),
.B(n_461),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_463),
.B(n_214),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_452),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_437),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_462),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_424),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_456),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_491),
.B(n_495),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_456),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_465),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_465),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_469),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_426),
.B(n_417),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_471),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_471),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_473),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_476),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_476),
.Y(n_595)
);

BUFx8_ASAP7_75t_L g596 ( 
.A(n_517),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_484),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_484),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_504),
.B(n_386),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_502),
.B(n_387),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_502),
.B(n_305),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_500),
.B(n_417),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_503),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_434),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_486),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_486),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_489),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_489),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_490),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_308),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_490),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_504),
.B(n_318),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_477),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_512),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_492),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_580),
.B(n_470),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_583),
.B(n_517),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_583),
.B(n_478),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_580),
.B(n_479),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_583),
.B(n_485),
.Y(n_622)
);

AOI21x1_ASAP7_75t_L g623 ( 
.A1(n_563),
.A2(n_475),
.B(n_329),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_535),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_535),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_539),
.B(n_488),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_537),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_612),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_545),
.B(n_499),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_537),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_540),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_583),
.B(n_505),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_549),
.B(n_460),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_612),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_572),
.B(n_511),
.C(n_481),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_589),
.B(n_515),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_555),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_579),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_555),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_525),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_532),
.B(n_526),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_538),
.B(n_528),
.Y(n_642)
);

OAI21xp33_ASAP7_75t_SL g643 ( 
.A1(n_611),
.A2(n_467),
.B(n_507),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_602),
.B(n_290),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_579),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_615),
.B(n_616),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_579),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_540),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_579),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_572),
.A2(n_442),
.B1(n_443),
.B2(n_438),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_587),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_555),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_589),
.B(n_530),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_541),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_538),
.B(n_508),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_587),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_604),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_602),
.A2(n_472),
.B1(n_433),
.B2(n_428),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_596),
.B(n_483),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_538),
.B(n_546),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_596),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_587),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_587),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_596),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_612),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_541),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_596),
.B(n_524),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_549),
.B(n_538),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_568),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_568),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_546),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_568),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_534),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_581),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_615),
.B(n_507),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_550),
.B(n_510),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_577),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_550),
.B(n_510),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_534),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_611),
.B(n_513),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_615),
.B(n_616),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_612),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_550),
.A2(n_398),
.B1(n_400),
.B2(n_393),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_577),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_542),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_616),
.B(n_513),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_542),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_612),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_577),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_585),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_550),
.Y(n_693)
);

BUFx4f_ASAP7_75t_L g694 ( 
.A(n_612),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_600),
.A2(n_403),
.B1(n_401),
.B2(n_494),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_543),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_578),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_543),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_SL g699 ( 
.A1(n_566),
.A2(n_497),
.B1(n_498),
.B2(n_496),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_570),
.B(n_422),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_600),
.B(n_514),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_531),
.B(n_425),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_548),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_561),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_612),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_600),
.A2(n_560),
.B1(n_599),
.B2(n_607),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_562),
.B(n_560),
.Y(n_707)
);

BUFx4f_ASAP7_75t_L g708 ( 
.A(n_567),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_562),
.B(n_514),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_574),
.B(n_464),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_599),
.B(n_566),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_605),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_585),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_567),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_560),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_603),
.B(n_520),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_585),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_614),
.B(n_258),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_551),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_570),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_533),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_603),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_566),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_598),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_553),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_600),
.B(n_599),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_533),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_569),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_553),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_536),
.B(n_520),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_569),
.B(n_529),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_557),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_557),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_606),
.B(n_522),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_607),
.A2(n_229),
.B1(n_333),
.B2(n_366),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_558),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_544),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_558),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_559),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_559),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_567),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_571),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_571),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_608),
.A2(n_529),
.B1(n_522),
.B2(n_523),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_575),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_575),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_614),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_606),
.B(n_523),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_561),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_582),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_598),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_606),
.B(n_245),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_566),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_SL g757 ( 
.A(n_544),
.B(n_509),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_608),
.Y(n_758)
);

BUFx4f_ASAP7_75t_L g759 ( 
.A(n_567),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_260),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_610),
.B(n_245),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_563),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_582),
.Y(n_763)
);

BUFx8_ASAP7_75t_SL g764 ( 
.A(n_610),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_598),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_586),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_586),
.B(n_290),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_547),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_567),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_565),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_768),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_L g772 ( 
.A(n_663),
.B(n_216),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_624),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_733),
.B(n_216),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_750),
.B(n_762),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_762),
.B(n_610),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_770),
.B(n_610),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_768),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_723),
.B(n_516),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_770),
.B(n_217),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_626),
.B(n_609),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_641),
.B(n_250),
.C(n_246),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_662),
.B(n_565),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_625),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_726),
.B(n_439),
.Y(n_785)
);

AO22x2_ASAP7_75t_L g786 ( 
.A1(n_635),
.A2(n_734),
.B1(n_730),
.B2(n_731),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_625),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_723),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_L g790 ( 
.A(n_711),
.B(n_250),
.C(n_246),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_673),
.B(n_217),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_675),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_707),
.A2(n_601),
.B(n_573),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_673),
.B(n_573),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_642),
.B(n_601),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_682),
.B(n_609),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_675),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_682),
.B(n_613),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_682),
.B(n_613),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_657),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_682),
.B(n_617),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_710),
.B(n_617),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_620),
.B(n_328),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_646),
.B(n_617),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_663),
.B(n_218),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_622),
.B(n_331),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_646),
.B(n_588),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_683),
.B(n_588),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_683),
.B(n_590),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_666),
.B(n_394),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_632),
.B(n_335),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_627),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_726),
.B(n_466),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_650),
.B(n_640),
.C(n_629),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_751),
.B(n_590),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_756),
.B(n_518),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_671),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_751),
.B(n_592),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_630),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_630),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_755),
.B(n_592),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_666),
.B(n_218),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_681),
.B(n_734),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_670),
.B(n_349),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_681),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_671),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_672),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_729),
.A2(n_597),
.B1(n_594),
.B2(n_552),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_628),
.B(n_225),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_755),
.B(n_594),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_693),
.B(n_350),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_672),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_628),
.B(n_225),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_693),
.B(n_352),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_694),
.A2(n_597),
.B(n_332),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_628),
.B(n_228),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_761),
.B(n_303),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_729),
.A2(n_547),
.B1(n_552),
.B2(n_554),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_706),
.A2(n_394),
.B1(n_395),
.B2(n_399),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_655),
.B(n_519),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_674),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_761),
.B(n_374),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_674),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_725),
.A2(n_554),
.B1(n_547),
.B2(n_552),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_657),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_631),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_644),
.A2(n_228),
.B1(n_252),
.B2(n_244),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_756),
.B(n_521),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_619),
.A2(n_407),
.B1(n_408),
.B2(n_410),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_700),
.B(n_714),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_657),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_660),
.B(n_527),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_677),
.B(n_384),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_633),
.B(n_408),
.C(n_407),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_677),
.B(n_688),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_628),
.B(n_231),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_679),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_758),
.A2(n_554),
.B1(n_556),
.B2(n_564),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_688),
.B(n_231),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_676),
.B(n_468),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_679),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_644),
.B(n_232),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_628),
.B(n_232),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_644),
.B(n_234),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_644),
.B(n_234),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_644),
.B(n_236),
.Y(n_866)
);

AND2x4_ASAP7_75t_SL g867 ( 
.A(n_676),
.B(n_740),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_631),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_644),
.B(n_236),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_644),
.B(n_237),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_697),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_648),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_693),
.A2(n_619),
.B1(n_701),
.B2(n_643),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_700),
.B(n_412),
.C(n_410),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_701),
.B(n_237),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_760),
.B(n_238),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_718),
.B(n_238),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_694),
.A2(n_336),
.B(n_319),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_648),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_676),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_697),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_636),
.B(n_239),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_654),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_618),
.B(n_356),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_686),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_695),
.B(n_482),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_712),
.B(n_239),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_654),
.Y(n_888)
);

NOR2x1p5_ASAP7_75t_L g889 ( 
.A(n_678),
.B(n_412),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_712),
.B(n_240),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_757),
.Y(n_891)
);

OAI221xp5_ASAP7_75t_L g892 ( 
.A1(n_685),
.A2(n_415),
.B1(n_416),
.B2(n_365),
.C(n_369),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_668),
.A2(n_556),
.B1(n_564),
.B2(n_561),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_712),
.B(n_240),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_619),
.A2(n_712),
.B1(n_653),
.B2(n_669),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_L g896 ( 
.A(n_634),
.B(n_241),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_668),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_687),
.A2(n_556),
.B1(n_564),
.B2(n_561),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_687),
.A2(n_561),
.B1(n_593),
.B2(n_591),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_621),
.B(n_357),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_712),
.B(n_487),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_619),
.B(n_360),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_712),
.B(n_241),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_661),
.B(n_345),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_712),
.B(n_242),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_652),
.B(n_638),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_689),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_658),
.B(n_361),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_702),
.B(n_242),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_638),
.B(n_244),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_638),
.B(n_252),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_689),
.Y(n_912)
);

BUFx6f_ASAP7_75t_SL g913 ( 
.A(n_740),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_696),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_737),
.B(n_389),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_634),
.B(n_389),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_658),
.B(n_397),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_680),
.B(n_397),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_740),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_696),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_634),
.B(n_402),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_698),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_658),
.B(n_402),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_686),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_659),
.B(n_415),
.C(n_380),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_659),
.B(n_413),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_659),
.B(n_413),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_691),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_691),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_634),
.B(n_414),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_637),
.A2(n_414),
.B1(n_418),
.B2(n_419),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_698),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_637),
.B(n_364),
.Y(n_933)
);

NAND2x1_ASAP7_75t_L g934 ( 
.A(n_637),
.B(n_561),
.Y(n_934)
);

NAND2x1_ASAP7_75t_L g935 ( 
.A(n_639),
.B(n_567),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_719),
.B(n_724),
.C(n_699),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_639),
.B(n_418),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_703),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_SL g939 ( 
.A(n_703),
.B(n_367),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_764),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_738),
.B(n_376),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_639),
.A2(n_347),
.B1(n_351),
.B2(n_368),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_773),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_906),
.A2(n_694),
.B(n_708),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_867),
.B(n_747),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_935),
.Y(n_946)
);

CKINVDCx10_ASAP7_75t_R g947 ( 
.A(n_913),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_793),
.A2(n_759),
.B(n_708),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_867),
.B(n_709),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_783),
.A2(n_647),
.B(n_645),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_814),
.B(n_645),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_792),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_781),
.A2(n_777),
.B(n_776),
.Y(n_953)
);

AOI33xp33_ASAP7_75t_L g954 ( 
.A1(n_797),
.A2(n_722),
.A3(n_763),
.B1(n_753),
.B2(n_749),
.B3(n_748),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_783),
.A2(n_649),
.B(n_647),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_795),
.B(n_794),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_795),
.B(n_709),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_794),
.B(n_713),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_775),
.B(n_649),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_802),
.A2(n_759),
.B(n_708),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_855),
.A2(n_665),
.B(n_664),
.C(n_651),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_771),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_771),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_871),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_919),
.B(n_713),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_788),
.Y(n_966)
);

O2A1O1Ixp5_ASAP7_75t_L g967 ( 
.A1(n_821),
.A2(n_623),
.B(n_742),
.C(n_766),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_784),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_780),
.B(n_651),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_873),
.B(n_634),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_782),
.B(n_385),
.C(n_382),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_804),
.A2(n_664),
.B(n_656),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_823),
.B(n_722),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_815),
.A2(n_759),
.B(n_721),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_837),
.B(n_728),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_779),
.B(n_728),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_818),
.A2(n_721),
.B(n_665),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_780),
.B(n_803),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_850),
.B(n_735),
.C(n_732),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_842),
.B(n_803),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_806),
.B(n_732),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_806),
.B(n_656),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_811),
.B(n_735),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_825),
.B(n_736),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_881),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_811),
.A2(n_749),
.B(n_766),
.C(n_742),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_909),
.B(n_690),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_830),
.A2(n_684),
.B(n_667),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_787),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_789),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_831),
.A2(n_739),
.B(n_736),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_853),
.B(n_831),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_812),
.A2(n_745),
.B1(n_741),
.B2(n_763),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_807),
.A2(n_741),
.B(n_739),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_790),
.B(n_667),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_808),
.A2(n_684),
.B(n_667),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_880),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_774),
.B(n_684),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_880),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_824),
.B(n_705),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_834),
.A2(n_748),
.B1(n_745),
.B2(n_746),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_809),
.A2(n_746),
.B(n_743),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_934),
.A2(n_705),
.B(n_743),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_913),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_796),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_923),
.A2(n_705),
.B(n_753),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_800),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_824),
.B(n_623),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_875),
.B(n_717),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_834),
.B(n_692),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_819),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_926),
.A2(n_769),
.B(n_717),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_798),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_895),
.B(n_690),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_927),
.A2(n_769),
.B(n_717),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_859),
.B(n_692),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_910),
.A2(n_911),
.B(n_846),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_800),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_908),
.B(n_715),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_845),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_778),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_820),
.A2(n_769),
.B(n_744),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_908),
.B(n_933),
.C(n_900),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_933),
.B(n_799),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_839),
.A2(n_744),
.B(n_765),
.C(n_720),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_840),
.B(n_852),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_868),
.B(n_715),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_845),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_872),
.B(n_720),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_879),
.B(n_727),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_860),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_918),
.A2(n_744),
.B(n_754),
.C(n_765),
.Y(n_1032)
);

AOI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_884),
.A2(n_754),
.B(n_727),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_883),
.A2(n_690),
.B(n_752),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_888),
.B(n_690),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_897),
.B(n_690),
.Y(n_1036)
);

AND2x2_ASAP7_75t_SL g1037 ( 
.A(n_772),
.B(n_375),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_907),
.B(n_912),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_914),
.A2(n_752),
.B(n_704),
.Y(n_1039)
);

NOR2x2_ASAP7_75t_L g1040 ( 
.A(n_813),
.B(n_7),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_785),
.Y(n_1041)
);

OAI321xp33_ASAP7_75t_L g1042 ( 
.A1(n_892),
.A2(n_941),
.A3(n_849),
.B1(n_884),
.B2(n_900),
.C(n_942),
.Y(n_1042)
);

OAI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_920),
.A2(n_406),
.B1(n_390),
.B2(n_404),
.Y(n_1043)
);

OAI321xp33_ASAP7_75t_L g1044 ( 
.A1(n_902),
.A2(n_405),
.A3(n_595),
.B1(n_584),
.B2(n_567),
.C(n_593),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_886),
.B(n_584),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_922),
.Y(n_1046)
);

NOR2x2_ASAP7_75t_L g1047 ( 
.A(n_813),
.B(n_9),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_932),
.B(n_752),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_938),
.A2(n_752),
.B(n_704),
.C(n_716),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_835),
.A2(n_704),
.B(n_716),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_851),
.A2(n_752),
.B(n_704),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_887),
.A2(n_716),
.B(n_704),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_876),
.B(n_716),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_801),
.A2(n_716),
.B(n_767),
.Y(n_1054)
);

AOI33xp33_ASAP7_75t_L g1055 ( 
.A1(n_828),
.A2(n_931),
.A3(n_816),
.B1(n_848),
.B2(n_874),
.B3(n_785),
.Y(n_1055)
);

NAND2x1p5_ASAP7_75t_L g1056 ( 
.A(n_851),
.B(n_584),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_917),
.A2(n_313),
.B(n_254),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_902),
.A2(n_584),
.B(n_591),
.C(n_593),
.Y(n_1058)
);

OAI21xp33_ASAP7_75t_L g1059 ( 
.A1(n_915),
.A2(n_877),
.B(n_791),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_854),
.B(n_388),
.C(n_282),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_828),
.A2(n_584),
.B1(n_591),
.B2(n_593),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_817),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_937),
.A2(n_921),
.B(n_833),
.C(n_856),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_833),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_826),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_826),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_827),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_822),
.A2(n_584),
.B1(n_591),
.B2(n_593),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_891),
.B(n_253),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_836),
.A2(n_863),
.B(n_930),
.C(n_856),
.Y(n_1070)
);

OAI321xp33_ASAP7_75t_L g1071 ( 
.A1(n_904),
.A2(n_847),
.A3(n_822),
.B1(n_925),
.B2(n_930),
.C(n_836),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_939),
.B(n_255),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_940),
.B(n_261),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_827),
.B(n_263),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_863),
.A2(n_584),
.B1(n_593),
.B2(n_595),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_832),
.A2(n_767),
.B(n_330),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_916),
.A2(n_324),
.B(n_269),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_832),
.B(n_265),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_816),
.B(n_848),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_878),
.A2(n_595),
.B(n_591),
.C(n_593),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_904),
.B(n_10),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_841),
.A2(n_767),
.B(n_337),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_810),
.A2(n_595),
.B(n_591),
.C(n_284),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_843),
.B(n_273),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_786),
.B(n_591),
.Y(n_1085)
);

BUFx12f_ASAP7_75t_L g1086 ( 
.A(n_813),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_843),
.A2(n_595),
.B(n_277),
.C(n_283),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_857),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_857),
.B(n_279),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_901),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_916),
.A2(n_344),
.B(n_287),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_904),
.B(n_14),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_786),
.B(n_595),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_921),
.A2(n_861),
.B(n_929),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_901),
.B(n_286),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_889),
.B(n_767),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_805),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_885),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_885),
.B(n_595),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_924),
.B(n_289),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_890),
.A2(n_767),
.B(n_258),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_882),
.Y(n_1102)
);

CKINVDCx6p67_ASAP7_75t_R g1103 ( 
.A(n_862),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_936),
.B(n_298),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_928),
.A2(n_929),
.B(n_905),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_894),
.Y(n_1106)
);

AO21x1_ASAP7_75t_L g1107 ( 
.A1(n_903),
.A2(n_258),
.B(n_767),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_838),
.B(n_300),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_864),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_829),
.A2(n_258),
.B(n_767),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_896),
.A2(n_421),
.B(n_383),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_865),
.A2(n_869),
.B(n_866),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_870),
.A2(n_373),
.B(n_372),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_838),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_786),
.A2(n_371),
.B(n_370),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_899),
.A2(n_359),
.B(n_358),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_893),
.B(n_16),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_893),
.B(n_354),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_844),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_844),
.B(n_858),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_898),
.B(n_348),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_898),
.B(n_342),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_899),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_858),
.A2(n_339),
.B(n_315),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_795),
.B(n_312),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_814),
.A2(n_292),
.B(n_290),
.C(n_21),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_814),
.A2(n_292),
.B(n_290),
.C(n_21),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_800),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_871),
.B(n_292),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_999),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_956),
.A2(n_1023),
.B1(n_957),
.B2(n_978),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_978),
.A2(n_292),
.B(n_290),
.C(n_258),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_973),
.B(n_19),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_958),
.A2(n_292),
.B(n_89),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_SL g1135 ( 
.A(n_964),
.B(n_20),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1086),
.B(n_20),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_980),
.B(n_32),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_981),
.A2(n_92),
.B(n_210),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1052),
.A2(n_258),
.B(n_202),
.Y(n_1139)
);

CKINVDCx11_ASAP7_75t_R g1140 ( 
.A(n_1004),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_985),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_943),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_979),
.B(n_34),
.Y(n_1143)
);

OAI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1042),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_985),
.B(n_39),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_992),
.A2(n_41),
.B1(n_42),
.B2(n_46),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1026),
.B(n_42),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_952),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_976),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1037),
.B(n_258),
.Y(n_1150)
);

AND2x2_ASAP7_75t_SL g1151 ( 
.A(n_1037),
.B(n_46),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_979),
.B(n_47),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_962),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_983),
.A2(n_109),
.B(n_188),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_963),
.Y(n_1155)
);

AND2x2_ASAP7_75t_SL g1156 ( 
.A(n_1081),
.B(n_1092),
.Y(n_1156)
);

BUFx2_ASAP7_75t_SL g1157 ( 
.A(n_1004),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1125),
.A2(n_47),
.B(n_50),
.C(n_51),
.Y(n_1158)
);

NAND2x1_ASAP7_75t_L g1159 ( 
.A(n_1007),
.B(n_111),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_947),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1105),
.A2(n_258),
.B(n_118),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_968),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1123),
.B(n_52),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1005),
.B(n_52),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_945),
.B(n_1079),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_984),
.B(n_53),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1031),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_953),
.A2(n_122),
.B(n_180),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1010),
.A2(n_104),
.B(n_175),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_989),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_990),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1005),
.B(n_55),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1024),
.A2(n_95),
.B(n_167),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1008),
.A2(n_982),
.B(n_1000),
.C(n_951),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1013),
.B(n_57),
.Y(n_1175)
);

CKINVDCx8_ASAP7_75t_R g1176 ( 
.A(n_1090),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1065),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1041),
.B(n_60),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1013),
.B(n_60),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_986),
.A2(n_61),
.B(n_62),
.C(n_66),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_966),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_949),
.B(n_61),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_949),
.B(n_62),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_945),
.B(n_965),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1019),
.A2(n_128),
.B(n_166),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_965),
.B(n_66),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_997),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_997),
.Y(n_1188)
);

NAND2x1_ASAP7_75t_L g1189 ( 
.A(n_1007),
.B(n_132),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_991),
.A2(n_126),
.B(n_154),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1129),
.B(n_68),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_975),
.B(n_69),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_959),
.B(n_73),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1001),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1073),
.B(n_143),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_982),
.A2(n_146),
.B1(n_149),
.B2(n_182),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1038),
.A2(n_1000),
.B1(n_1046),
.B2(n_1011),
.Y(n_1197)
);

BUFx4f_ASAP7_75t_L g1198 ( 
.A(n_1103),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1104),
.B(n_1069),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1021),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1123),
.A2(n_993),
.B1(n_994),
.B2(n_1002),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_967),
.A2(n_951),
.B(n_969),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_959),
.B(n_1045),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_954),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_971),
.A2(n_1081),
.B(n_1092),
.C(n_1059),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1040),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1085),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1093),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1065),
.Y(n_1209)
);

NAND2x1p5_ASAP7_75t_L g1210 ( 
.A(n_1018),
.B(n_1020),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1066),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1018),
.B(n_1020),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1093),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1071),
.B(n_971),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_R g1215 ( 
.A(n_1102),
.B(n_1008),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1096),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1115),
.B(n_1043),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_1035),
.A2(n_1036),
.B(n_950),
.C(n_955),
.Y(n_1219)
);

BUFx8_ASAP7_75t_SL g1220 ( 
.A(n_946),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1067),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1018),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1043),
.B(n_995),
.Y(n_1223)
);

OR2x6_ASAP7_75t_L g1224 ( 
.A(n_1120),
.B(n_1114),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1095),
.Y(n_1225)
);

AND2x2_ASAP7_75t_SL g1226 ( 
.A(n_1117),
.B(n_1055),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_R g1227 ( 
.A(n_1117),
.B(n_995),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1016),
.B(n_1009),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_969),
.B(n_998),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1063),
.A2(n_1009),
.B(n_1127),
.C(n_1126),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1119),
.B(n_1062),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_970),
.A2(n_1014),
.B(n_1101),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1064),
.B(n_1097),
.Y(n_1233)
);

NOR2xp67_ASAP7_75t_L g1234 ( 
.A(n_1072),
.B(n_998),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1022),
.A2(n_1017),
.B(n_1060),
.C(n_948),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1060),
.A2(n_961),
.B(n_1058),
.C(n_1070),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1088),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1070),
.A2(n_967),
.B(n_1032),
.C(n_1083),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_970),
.A2(n_1044),
.B(n_1025),
.C(n_1033),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1047),
.A2(n_1108),
.B1(n_1121),
.B2(n_1122),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1065),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1098),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_960),
.A2(n_944),
.B(n_1053),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1048),
.A2(n_1030),
.B1(n_1027),
.B2(n_1029),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1062),
.B(n_1128),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1049),
.B(n_1054),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1018),
.B(n_1028),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_974),
.A2(n_977),
.B(n_1015),
.Y(n_1248)
);

OAI22x1_ASAP7_75t_L g1249 ( 
.A1(n_1109),
.A2(n_987),
.B1(n_1099),
.B2(n_1128),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1012),
.A2(n_1034),
.B(n_1006),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_988),
.A2(n_996),
.B(n_1039),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1065),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1074),
.B(n_1084),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1020),
.B(n_1028),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1078),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1020),
.B(n_1028),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_972),
.A2(n_1094),
.B(n_1003),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1028),
.B(n_1089),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1080),
.A2(n_1112),
.B(n_1087),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1099),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1051),
.A2(n_1050),
.B(n_1056),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_946),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1100),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1106),
.B(n_946),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1106),
.B(n_946),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1106),
.B(n_1124),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1076),
.A2(n_1082),
.B(n_1091),
.C(n_1077),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1106),
.B(n_1118),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1061),
.C(n_1057),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1056),
.Y(n_1270)
);

AO32x1_ASAP7_75t_L g1271 ( 
.A1(n_1075),
.A2(n_1068),
.A3(n_1107),
.B1(n_1110),
.B2(n_1111),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_964),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1004),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1052),
.A2(n_970),
.B(n_1014),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_956),
.A2(n_957),
.B(n_958),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_956),
.A2(n_957),
.B(n_958),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_964),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_956),
.B(n_750),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_956),
.B(n_750),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_956),
.B(n_788),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_967),
.A2(n_1070),
.B(n_1094),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_L g1282 ( 
.A(n_1004),
.B(n_880),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1023),
.B(n_978),
.C(n_814),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1026),
.B(n_823),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_943),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_964),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_978),
.A2(n_697),
.B1(n_814),
.B2(n_641),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_999),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1165),
.B(n_1216),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1174),
.A2(n_1283),
.B(n_1201),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1131),
.Y(n_1291)
);

AOI221x1_ASAP7_75t_L g1292 ( 
.A1(n_1223),
.A2(n_1217),
.B1(n_1283),
.B2(n_1194),
.C(n_1146),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1220),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1149),
.B(n_1287),
.Y(n_1296)
);

NOR4xp25_ASAP7_75t_L g1297 ( 
.A(n_1144),
.B(n_1205),
.C(n_1214),
.D(n_1158),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1198),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1251),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1261),
.A2(n_1197),
.B(n_1228),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1250),
.A2(n_1161),
.B(n_1257),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1219),
.A2(n_1244),
.B(n_1202),
.Y(n_1302)
);

AO32x2_ASAP7_75t_L g1303 ( 
.A1(n_1240),
.A2(n_1196),
.A3(n_1225),
.B1(n_1224),
.B2(n_1163),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1246),
.A2(n_1235),
.B(n_1257),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1199),
.A2(n_1229),
.B(n_1137),
.C(n_1147),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1151),
.A2(n_1164),
.B(n_1193),
.C(n_1152),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1232),
.A2(n_1274),
.B(n_1139),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1156),
.B(n_1284),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1262),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1163),
.B(n_1227),
.C(n_1215),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1268),
.A2(n_1239),
.A3(n_1249),
.B(n_1132),
.Y(n_1311)
);

BUFx8_ASAP7_75t_SL g1312 ( 
.A(n_1160),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1141),
.B(n_1184),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1162),
.Y(n_1314)
);

NOR2xp67_ASAP7_75t_L g1315 ( 
.A(n_1187),
.B(n_1254),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1143),
.A2(n_1192),
.B(n_1253),
.C(n_1263),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1259),
.A2(n_1238),
.B(n_1266),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1259),
.A2(n_1168),
.B(n_1236),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1246),
.A2(n_1230),
.B(n_1267),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1281),
.A2(n_1134),
.B(n_1190),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1269),
.A2(n_1231),
.A3(n_1203),
.B(n_1260),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1170),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1167),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1281),
.A2(n_1185),
.B(n_1169),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1240),
.B(n_1255),
.Y(n_1325)
);

BUFx2_ASAP7_75t_R g1326 ( 
.A(n_1277),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1171),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1148),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1181),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_R g1330 ( 
.A(n_1145),
.B(n_1166),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1138),
.A2(n_1154),
.B(n_1159),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1173),
.A2(n_1247),
.B(n_1271),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1271),
.A2(n_1256),
.B(n_1258),
.Y(n_1333)
);

BUFx4f_ASAP7_75t_SL g1334 ( 
.A(n_1272),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1204),
.B(n_1226),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1130),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1271),
.A2(n_1245),
.B(n_1280),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1189),
.A2(n_1195),
.B(n_1133),
.C(n_1175),
.Y(n_1338)
);

NOR2x1_ASAP7_75t_R g1339 ( 
.A(n_1140),
.B(n_1286),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1176),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1233),
.A2(n_1234),
.B(n_1270),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1187),
.B(n_1198),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1273),
.Y(n_1343)
);

O2A1O1Ixp5_ASAP7_75t_L g1344 ( 
.A1(n_1150),
.A2(n_1172),
.B(n_1191),
.C(n_1265),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1186),
.A2(n_1179),
.B1(n_1183),
.B2(n_1224),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1285),
.Y(n_1346)
);

AND2x6_ASAP7_75t_L g1347 ( 
.A(n_1208),
.B(n_1213),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1233),
.A2(n_1212),
.B(n_1210),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1222),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1210),
.A2(n_1212),
.B(n_1264),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1180),
.A2(n_1177),
.B(n_1241),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1237),
.A2(n_1242),
.B(n_1182),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1208),
.A2(n_1213),
.B(n_1178),
.C(n_1207),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1177),
.A2(n_1241),
.B(n_1209),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1136),
.A2(n_1206),
.B(n_1165),
.C(n_1282),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1224),
.B(n_1288),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1286),
.B(n_1130),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1155),
.A2(n_1200),
.B(n_1221),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1209),
.A2(n_1252),
.B(n_1187),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1218),
.A2(n_1188),
.B(n_1211),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1218),
.A2(n_1188),
.B(n_1273),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1273),
.A2(n_1157),
.B(n_1181),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1136),
.A2(n_1288),
.B1(n_1130),
.B2(n_1135),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1288),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1136),
.A2(n_978),
.B(n_1223),
.C(n_814),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1287),
.B(n_1223),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1141),
.Y(n_1369)
);

AOI221x1_ASAP7_75t_L g1370 ( 
.A1(n_1223),
.A2(n_1217),
.B1(n_1283),
.B2(n_1131),
.C(n_1023),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1174),
.A2(n_1283),
.B(n_1201),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1375)
);

CKINVDCx8_ASAP7_75t_R g1376 ( 
.A(n_1160),
.Y(n_1376)
);

BUFx2_ASAP7_75t_R g1377 ( 
.A(n_1160),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1220),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1243),
.A2(n_1259),
.B(n_1202),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1153),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1287),
.B(n_871),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1156),
.B(n_823),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1130),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1142),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1251),
.Y(n_1388)
);

AND2x6_ASAP7_75t_L g1389 ( 
.A(n_1208),
.B(n_1213),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1160),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1287),
.B(n_1023),
.C(n_1223),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1251),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1223),
.A2(n_978),
.B(n_814),
.C(n_1023),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1153),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1243),
.A2(n_1174),
.A3(n_1008),
.B(n_1201),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1130),
.Y(n_1400)
);

AO21x1_ASAP7_75t_L g1401 ( 
.A1(n_1223),
.A2(n_1214),
.B(n_1163),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1243),
.A2(n_1259),
.B(n_1202),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1205),
.A2(n_1197),
.B(n_1201),
.Y(n_1403)
);

OAI22x1_ASAP7_75t_L g1404 ( 
.A1(n_1287),
.A2(n_1223),
.B1(n_1214),
.B2(n_1081),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_SL g1405 ( 
.A1(n_1131),
.A2(n_956),
.B(n_1023),
.C(n_957),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1160),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1223),
.A2(n_956),
.B1(n_1287),
.B2(n_1131),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1287),
.B(n_1223),
.Y(n_1408)
);

NOR2xp67_ASAP7_75t_L g1409 ( 
.A(n_1283),
.B(n_1023),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1174),
.A2(n_1283),
.B(n_1201),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1262),
.Y(n_1412)
);

NAND4xp25_ASAP7_75t_L g1413 ( 
.A(n_1287),
.B(n_635),
.C(n_782),
.D(n_641),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1414)
);

INVx3_ASAP7_75t_SL g1415 ( 
.A(n_1160),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1223),
.A2(n_1151),
.B1(n_1156),
.B2(n_1163),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1153),
.Y(n_1417)
);

AOI221x1_ASAP7_75t_L g1418 ( 
.A1(n_1223),
.A2(n_1217),
.B1(n_1283),
.B2(n_1131),
.C(n_1023),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1287),
.A2(n_956),
.B1(n_1223),
.B2(n_1023),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1250),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1220),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1174),
.A2(n_957),
.B(n_1223),
.Y(n_1423)
);

AO31x2_ASAP7_75t_L g1424 ( 
.A1(n_1243),
.A2(n_1174),
.A3(n_1008),
.B(n_1201),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1223),
.A2(n_978),
.B(n_814),
.C(n_1023),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1262),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1223),
.A2(n_978),
.B(n_814),
.C(n_1023),
.Y(n_1429)
);

AO31x2_ASAP7_75t_L g1430 ( 
.A1(n_1243),
.A2(n_1174),
.A3(n_1008),
.B(n_1201),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1287),
.B(n_871),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1251),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1220),
.Y(n_1435)
);

AO32x2_ASAP7_75t_L g1436 ( 
.A1(n_1201),
.A2(n_1131),
.A3(n_1240),
.B1(n_1197),
.B2(n_1194),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1262),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1187),
.B(n_1198),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1156),
.B(n_823),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1287),
.A2(n_956),
.B1(n_1223),
.B2(n_1023),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1243),
.A2(n_1174),
.A3(n_1008),
.B(n_1201),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_SL g1442 ( 
.A1(n_1131),
.A2(n_956),
.B(n_1023),
.C(n_957),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1223),
.A2(n_956),
.B1(n_1287),
.B2(n_1131),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1130),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1287),
.B(n_1223),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1243),
.A2(n_1174),
.A3(n_1008),
.B(n_1201),
.Y(n_1448)
);

NOR4xp25_ASAP7_75t_L g1449 ( 
.A(n_1144),
.B(n_1205),
.C(n_1283),
.D(n_1223),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1243),
.A2(n_1248),
.B(n_1251),
.Y(n_1450)
);

INVx3_ASAP7_75t_SL g1451 ( 
.A(n_1160),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1156),
.B(n_823),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1174),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1272),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1243),
.A2(n_1259),
.B(n_1202),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1294),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1416),
.A2(n_1408),
.B1(n_1368),
.B2(n_1446),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1349),
.Y(n_1458)
);

INVx3_ASAP7_75t_SL g1459 ( 
.A(n_1340),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1314),
.Y(n_1460)
);

INVx3_ASAP7_75t_SL g1461 ( 
.A(n_1415),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1308),
.B(n_1356),
.Y(n_1462)
);

BUFx10_ASAP7_75t_L g1463 ( 
.A(n_1349),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1323),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1369),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1336),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1385),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1416),
.A2(n_1401),
.B1(n_1404),
.B2(n_1325),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1454),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1395),
.A2(n_1407),
.B1(n_1444),
.B2(n_1310),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1322),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1395),
.A2(n_1407),
.B1(n_1444),
.B2(n_1419),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1423),
.A2(n_1440),
.B1(n_1306),
.B2(n_1429),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1346),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1412),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1386),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1345),
.A2(n_1403),
.B1(n_1431),
.B2(n_1383),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1413),
.A2(n_1452),
.B1(n_1384),
.B2(n_1439),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1413),
.A2(n_1290),
.B1(n_1411),
.B2(n_1372),
.Y(n_1480)
);

CKINVDCx11_ASAP7_75t_R g1481 ( 
.A(n_1376),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1406),
.Y(n_1482)
);

INVx8_ASAP7_75t_L g1483 ( 
.A(n_1312),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1397),
.A2(n_1425),
.B1(n_1365),
.B2(n_1305),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1290),
.A2(n_1411),
.B1(n_1372),
.B2(n_1409),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1451),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1393),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1303),
.A2(n_1363),
.B1(n_1335),
.B2(n_1296),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1400),
.Y(n_1489)
);

CKINVDCx6p67_ASAP7_75t_R g1490 ( 
.A(n_1393),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1409),
.A2(n_1382),
.B1(n_1398),
.B2(n_1417),
.Y(n_1491)
);

BUFx10_ASAP7_75t_L g1492 ( 
.A(n_1349),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_1357),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1316),
.A2(n_1319),
.B1(n_1392),
.B2(n_1414),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1370),
.B(n_1418),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1352),
.A2(n_1391),
.B1(n_1390),
.B2(n_1447),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1449),
.B(n_1291),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1445),
.Y(n_1498)
);

INVx3_ASAP7_75t_SL g1499 ( 
.A(n_1427),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1334),
.Y(n_1500)
);

CKINVDCx6p67_ASAP7_75t_R g1501 ( 
.A(n_1295),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1363),
.A2(n_1449),
.B1(n_1380),
.B2(n_1435),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1303),
.A2(n_1436),
.B1(n_1352),
.B2(n_1289),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1303),
.A2(n_1436),
.B1(n_1293),
.B2(n_1428),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1436),
.A2(n_1373),
.B1(n_1426),
.B2(n_1367),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1422),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1427),
.Y(n_1507)
);

CKINVDCx11_ASAP7_75t_R g1508 ( 
.A(n_1329),
.Y(n_1508)
);

INVx6_ASAP7_75t_L g1509 ( 
.A(n_1427),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1437),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1358),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1405),
.B(n_1442),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1377),
.Y(n_1513)
);

BUFx10_ASAP7_75t_L g1514 ( 
.A(n_1437),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1292),
.A2(n_1313),
.B1(n_1328),
.B2(n_1341),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1366),
.B(n_1371),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1374),
.B(n_1375),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1311),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1353),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1347),
.A2(n_1389),
.B1(n_1360),
.B2(n_1337),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1378),
.B(n_1387),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1321),
.Y(n_1522)
);

BUFx10_ASAP7_75t_L g1523 ( 
.A(n_1298),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1297),
.A2(n_1389),
.B1(n_1347),
.B2(n_1364),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1379),
.B(n_1432),
.Y(n_1525)
);

INVx8_ASAP7_75t_L g1526 ( 
.A(n_1389),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1389),
.Y(n_1527)
);

CKINVDCx16_ASAP7_75t_R g1528 ( 
.A(n_1326),
.Y(n_1528)
);

BUFx8_ASAP7_75t_SL g1529 ( 
.A(n_1339),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1311),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1438),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1394),
.A2(n_1434),
.B1(n_1453),
.B2(n_1443),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_1302),
.B2(n_1300),
.Y(n_1533)
);

CKINVDCx11_ASAP7_75t_R g1534 ( 
.A(n_1339),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1362),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1317),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1304),
.A2(n_1348),
.B1(n_1355),
.B2(n_1330),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1315),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1315),
.Y(n_1539)
);

INVx6_ASAP7_75t_L g1540 ( 
.A(n_1343),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1350),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1344),
.Y(n_1542)
);

BUFx8_ASAP7_75t_L g1543 ( 
.A(n_1297),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1381),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1351),
.Y(n_1545)
);

BUFx4f_ASAP7_75t_SL g1546 ( 
.A(n_1361),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1420),
.A2(n_1318),
.B(n_1455),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1402),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1455),
.A2(n_1332),
.B1(n_1333),
.B2(n_1320),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1359),
.A2(n_1354),
.B1(n_1331),
.B2(n_1307),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1420),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1338),
.Y(n_1552)
);

INVx3_ASAP7_75t_SL g1553 ( 
.A(n_1399),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1301),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1399),
.Y(n_1555)
);

INVx5_ASAP7_75t_L g1556 ( 
.A(n_1424),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1424),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1424),
.A2(n_1430),
.B(n_1448),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1299),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1430),
.A2(n_1441),
.B1(n_1448),
.B2(n_1324),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1430),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1441),
.A2(n_1448),
.B1(n_1396),
.B2(n_1433),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1441),
.A2(n_1416),
.B1(n_1444),
.B2(n_1407),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1388),
.A2(n_1151),
.B1(n_1217),
.B2(n_1156),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1450),
.A2(n_1217),
.B1(n_1151),
.B2(n_1223),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1323),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1336),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1294),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1342),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1356),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1416),
.A2(n_1444),
.B1(n_1407),
.B2(n_1408),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1336),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1336),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1294),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1294),
.Y(n_1575)
);

BUFx12f_ASAP7_75t_L g1576 ( 
.A(n_1454),
.Y(n_1576)
);

OAI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1416),
.A2(n_1163),
.B1(n_1287),
.B2(n_1042),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1416),
.A2(n_1163),
.B1(n_1287),
.B2(n_1042),
.Y(n_1578)
);

BUFx10_ASAP7_75t_L g1579 ( 
.A(n_1340),
.Y(n_1579)
);

INVx6_ASAP7_75t_L g1580 ( 
.A(n_1309),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1416),
.A2(n_1444),
.B(n_1407),
.Y(n_1581)
);

AOI21xp33_ASAP7_75t_L g1582 ( 
.A1(n_1404),
.A2(n_1223),
.B(n_1217),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1294),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1454),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1309),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1325),
.A2(n_1151),
.B1(n_1217),
.B2(n_1156),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1289),
.B(n_1252),
.Y(n_1587)
);

CKINVDCx11_ASAP7_75t_R g1588 ( 
.A(n_1376),
.Y(n_1588)
);

CKINVDCx11_ASAP7_75t_R g1589 ( 
.A(n_1376),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1416),
.A2(n_1163),
.B1(n_1287),
.B2(n_1042),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1407),
.B(n_1444),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1416),
.A2(n_1217),
.B1(n_1151),
.B2(n_1223),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1416),
.A2(n_1217),
.B1(n_1151),
.B2(n_1223),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1416),
.A2(n_1444),
.B1(n_1407),
.B2(n_1408),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1416),
.A2(n_1444),
.B1(n_1407),
.B2(n_1408),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1454),
.Y(n_1596)
);

INVx5_ASAP7_75t_L g1597 ( 
.A(n_1347),
.Y(n_1597)
);

BUFx4_ASAP7_75t_SL g1598 ( 
.A(n_1406),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1356),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1416),
.A2(n_1151),
.B1(n_1223),
.B2(n_1156),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1416),
.A2(n_1444),
.B1(n_1407),
.B2(n_1408),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1416),
.A2(n_1151),
.B1(n_1223),
.B2(n_1156),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1349),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1465),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1530),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1466),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1456),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1541),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1464),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1511),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1489),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1582),
.A2(n_1495),
.B(n_1547),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1563),
.B(n_1561),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1591),
.B(n_1563),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_SL g1615 ( 
.A1(n_1581),
.A2(n_1594),
.B(n_1571),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1522),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1591),
.B(n_1581),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1547),
.A2(n_1533),
.B(n_1532),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1464),
.Y(n_1619)
);

AO31x2_ASAP7_75t_L g1620 ( 
.A1(n_1532),
.A2(n_1557),
.A3(n_1555),
.B(n_1533),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1497),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1473),
.A2(n_1472),
.B(n_1571),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1536),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1513),
.B(n_1528),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1516),
.A2(n_1521),
.B(n_1517),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1518),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1460),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1553),
.B(n_1471),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1505),
.B(n_1480),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1474),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1567),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1566),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1475),
.B(n_1477),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1542),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1572),
.Y(n_1636)
);

AOI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1495),
.A2(n_1537),
.B(n_1517),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1598),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1568),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1516),
.A2(n_1525),
.B(n_1521),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1574),
.B(n_1575),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1583),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1525),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1545),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1535),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1595),
.B(n_1601),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1544),
.Y(n_1648)
);

AO31x2_ASAP7_75t_L g1649 ( 
.A1(n_1557),
.A2(n_1548),
.A3(n_1473),
.B(n_1601),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1481),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1544),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1485),
.B(n_1558),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1548),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1462),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1543),
.A2(n_1484),
.B1(n_1494),
.B2(n_1502),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1556),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1558),
.B(n_1470),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1582),
.A2(n_1578),
.B(n_1590),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1565),
.B(n_1556),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1543),
.A2(n_1586),
.B1(n_1592),
.B2(n_1593),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1556),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1526),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1527),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1494),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1562),
.A2(n_1550),
.B(n_1559),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1551),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1551),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1570),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1496),
.B(n_1504),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1526),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1588),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1512),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1554),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1560),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1573),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1484),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1554),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1493),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1457),
.B(n_1600),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1570),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1577),
.A2(n_1519),
.B(n_1515),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1549),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1524),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1520),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1537),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1599),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1599),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1602),
.A2(n_1564),
.B(n_1478),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1538),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1467),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1468),
.B(n_1488),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1493),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1479),
.B(n_1498),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1552),
.B(n_1539),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1491),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1546),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1587),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1540),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1458),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1499),
.B(n_1501),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1531),
.A2(n_1569),
.B(n_1523),
.Y(n_1702)
);

BUFx4f_ASAP7_75t_L g1703 ( 
.A(n_1507),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1507),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1603),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1523),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1469),
.A2(n_1596),
.B(n_1584),
.Y(n_1707)
);

BUFx4f_ASAP7_75t_SL g1708 ( 
.A(n_1500),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1463),
.A2(n_1514),
.B(n_1492),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1459),
.B(n_1461),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1463),
.B(n_1514),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1589),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1476),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1508),
.B(n_1482),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1604),
.B(n_1579),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1606),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1635),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1689),
.A2(n_1534),
.B(n_1483),
.C(n_1529),
.Y(n_1718)
);

OAI211xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1622),
.A2(n_1686),
.B(n_1706),
.C(n_1617),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1654),
.B(n_1490),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1652),
.B(n_1585),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1652),
.B(n_1509),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1627),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1627),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1646),
.A2(n_1506),
.B(n_1580),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1609),
.B(n_1619),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1630),
.B(n_1510),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1646),
.A2(n_1510),
.B(n_1576),
.C(n_1579),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1613),
.B(n_1486),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1629),
.A2(n_1483),
.B1(n_1487),
.B2(n_1670),
.C(n_1621),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1677),
.B(n_1633),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1647),
.A2(n_1483),
.B(n_1655),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1614),
.B(n_1697),
.Y(n_1733)
);

AO21x2_ASAP7_75t_L g1734 ( 
.A1(n_1683),
.A2(n_1637),
.B(n_1612),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1618),
.A2(n_1640),
.B(n_1625),
.Y(n_1735)
);

AND2x2_ASAP7_75t_SL g1736 ( 
.A(n_1657),
.B(n_1665),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1657),
.A2(n_1665),
.B(n_1686),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1669),
.B(n_1681),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1691),
.B(n_1634),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1697),
.B(n_1679),
.Y(n_1740)
);

AO21x2_ASAP7_75t_L g1741 ( 
.A1(n_1683),
.A2(n_1637),
.B(n_1612),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1660),
.A2(n_1692),
.B1(n_1680),
.B2(n_1684),
.C(n_1685),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1666),
.A2(n_1653),
.B(n_1667),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1673),
.B(n_1641),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1666),
.A2(n_1675),
.B(n_1668),
.Y(n_1745)
);

NOR2xp67_ASAP7_75t_L g1746 ( 
.A(n_1693),
.B(n_1695),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1688),
.B(n_1631),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1641),
.B(n_1631),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1620),
.B(n_1639),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1620),
.B(n_1642),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1680),
.A2(n_1692),
.B(n_1684),
.C(n_1685),
.Y(n_1751)
);

BUFx2_ASAP7_75t_SL g1752 ( 
.A(n_1606),
.Y(n_1752)
);

INVx3_ASAP7_75t_SL g1753 ( 
.A(n_1638),
.Y(n_1753)
);

OAI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1615),
.A2(n_1675),
.B(n_1643),
.C(n_1706),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1615),
.A2(n_1658),
.B1(n_1682),
.B2(n_1690),
.C(n_1607),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1659),
.A2(n_1694),
.B(n_1661),
.C(n_1696),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1611),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1687),
.B(n_1690),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1620),
.B(n_1612),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1620),
.B(n_1628),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1659),
.A2(n_1694),
.B(n_1661),
.C(n_1696),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1620),
.B(n_1628),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1610),
.B(n_1649),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_1708),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1610),
.B(n_1649),
.Y(n_1765)
);

OAI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1643),
.A2(n_1693),
.B(n_1668),
.C(n_1664),
.Y(n_1766)
);

OA21x2_ASAP7_75t_L g1767 ( 
.A1(n_1648),
.A2(n_1678),
.B(n_1651),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1649),
.B(n_1674),
.Y(n_1768)
);

AO21x2_ASAP7_75t_L g1769 ( 
.A1(n_1678),
.A2(n_1658),
.B(n_1682),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1701),
.A2(n_1710),
.B(n_1623),
.C(n_1700),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1649),
.B(n_1626),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1658),
.A2(n_1682),
.B(n_1699),
.C(n_1713),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1644),
.Y(n_1773)
);

AND2x2_ASAP7_75t_SL g1774 ( 
.A(n_1630),
.B(n_1702),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1630),
.A2(n_1663),
.B(n_1702),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1701),
.A2(n_1703),
.B1(n_1636),
.B2(n_1676),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1632),
.B(n_1636),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1648),
.B(n_1608),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1605),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1653),
.A2(n_1667),
.B(n_1656),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1623),
.B(n_1645),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1632),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1704),
.B(n_1705),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1616),
.B(n_1698),
.Y(n_1784)
);

INVx4_ASAP7_75t_SL g1785 ( 
.A(n_1727),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1773),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1749),
.B(n_1750),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1767),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1717),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1773),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1750),
.B(n_1760),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1717),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1763),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1780),
.Y(n_1794)
);

OR2x6_ASAP7_75t_SL g1795 ( 
.A(n_1765),
.B(n_1738),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1779),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1716),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1778),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1723),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1724),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1762),
.B(n_1656),
.Y(n_1801)
);

INVx4_ASAP7_75t_R g1802 ( 
.A(n_1716),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1781),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_SL g1804 ( 
.A1(n_1736),
.A2(n_1624),
.B1(n_1663),
.B2(n_1671),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1745),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1727),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1759),
.B(n_1739),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1764),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1768),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1755),
.B(n_1705),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1758),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1748),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1731),
.B(n_1747),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1781),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1784),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1745),
.B(n_1662),
.Y(n_1816)
);

NOR2xp67_ASAP7_75t_L g1817 ( 
.A(n_1766),
.B(n_1771),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1745),
.B(n_1733),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1818),
.B(n_1744),
.Y(n_1819)
);

AND2x2_ASAP7_75t_SL g1820 ( 
.A(n_1791),
.B(n_1736),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1807),
.B(n_1735),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1786),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1806),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1797),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1788),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1786),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1818),
.B(n_1790),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1817),
.A2(n_1742),
.B1(n_1719),
.B2(n_1769),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1785),
.B(n_1743),
.Y(n_1829)
);

OAI31xp33_ASAP7_75t_L g1830 ( 
.A1(n_1818),
.A2(n_1751),
.A3(n_1754),
.B(n_1718),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1789),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1807),
.B(n_1735),
.Y(n_1832)
);

INVxp67_ASAP7_75t_SL g1833 ( 
.A(n_1805),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1817),
.A2(n_1769),
.B1(n_1730),
.B2(n_1737),
.Y(n_1834)
);

OAI31xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1804),
.A2(n_1732),
.A3(n_1729),
.B(n_1770),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1791),
.A2(n_1729),
.B1(n_1741),
.B2(n_1734),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_L g1837 ( 
.A(n_1810),
.B(n_1772),
.C(n_1718),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1807),
.B(n_1735),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1811),
.B(n_1734),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1806),
.B(n_1774),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1787),
.B(n_1741),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1789),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1787),
.B(n_1726),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1791),
.B(n_1798),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1796),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1792),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1804),
.B(n_1746),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1794),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1811),
.B(n_1783),
.Y(n_1849)
);

INVx5_ASAP7_75t_L g1850 ( 
.A(n_1794),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1805),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1810),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1809),
.B(n_1756),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1844),
.B(n_1795),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1837),
.A2(n_1793),
.B1(n_1751),
.B2(n_1756),
.C(n_1761),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1852),
.B(n_1792),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1844),
.B(n_1795),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1844),
.B(n_1795),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1825),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1829),
.B(n_1816),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1830),
.A2(n_1721),
.B1(n_1722),
.B2(n_1793),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1852),
.B(n_1815),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1822),
.B(n_1815),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1821),
.B(n_1803),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1822),
.B(n_1812),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1850),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1821),
.B(n_1803),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1845),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1821),
.B(n_1801),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1821),
.B(n_1801),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1819),
.B(n_1813),
.Y(n_1871)
);

NAND4xp25_ASAP7_75t_SL g1872 ( 
.A(n_1830),
.B(n_1728),
.C(n_1725),
.D(n_1764),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1837),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1845),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1825),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1847),
.B(n_1808),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1822),
.B(n_1812),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1819),
.B(n_1813),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1829),
.B(n_1816),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1825),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1826),
.B(n_1799),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1832),
.B(n_1814),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1819),
.B(n_1827),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1842),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1838),
.B(n_1797),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1825),
.Y(n_1886)
);

INVx4_ASAP7_75t_L g1887 ( 
.A(n_1823),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1826),
.B(n_1800),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1864),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1854),
.B(n_1824),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1868),
.Y(n_1891)
);

NAND2x1_ASAP7_75t_SL g1892 ( 
.A(n_1887),
.B(n_1829),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1854),
.B(n_1824),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1864),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1868),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1873),
.B(n_1835),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1887),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1874),
.Y(n_1898)
);

NAND2x1_ASAP7_75t_L g1899 ( 
.A(n_1887),
.B(n_1802),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1874),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1871),
.B(n_1827),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1854),
.B(n_1820),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1873),
.B(n_1835),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1864),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1861),
.A2(n_1820),
.B1(n_1828),
.B2(n_1834),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1871),
.B(n_1843),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1856),
.B(n_1846),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1856),
.B(n_1846),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1857),
.B(n_1820),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1881),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1862),
.B(n_1849),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1881),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1862),
.B(n_1849),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1867),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1857),
.B(n_1820),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1888),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1888),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1884),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1871),
.B(n_1843),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1876),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1884),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1861),
.B(n_1843),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1878),
.B(n_1831),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1863),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1887),
.B(n_1829),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1887),
.B(n_1775),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1867),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1863),
.Y(n_1928)
);

AOI211xp5_ASAP7_75t_L g1929 ( 
.A1(n_1872),
.A2(n_1847),
.B(n_1833),
.C(n_1851),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1857),
.B(n_1823),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1865),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1858),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1865),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1877),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1877),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1902),
.B(n_1858),
.Y(n_1936)
);

INVxp33_ASAP7_75t_SL g1937 ( 
.A(n_1896),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1903),
.B(n_1878),
.Y(n_1938)
);

NOR2xp67_ASAP7_75t_L g1939 ( 
.A(n_1932),
.B(n_1872),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1906),
.B(n_1878),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1891),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1906),
.B(n_1883),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1891),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1902),
.B(n_1858),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1909),
.B(n_1869),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1919),
.B(n_1883),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1898),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1909),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1898),
.Y(n_1949)
);

OA211x2_ASAP7_75t_L g1950 ( 
.A1(n_1899),
.A2(n_1876),
.B(n_1714),
.C(n_1740),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1919),
.B(n_1885),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1929),
.B(n_1836),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1920),
.B(n_1753),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1915),
.B(n_1869),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1923),
.B(n_1883),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1918),
.B(n_1885),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1932),
.B(n_1860),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1900),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1889),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1900),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1915),
.B(n_1869),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1930),
.B(n_1870),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1895),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1911),
.B(n_1885),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1921),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1930),
.B(n_1870),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1889),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1913),
.B(n_1855),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1897),
.B(n_1753),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1910),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1890),
.Y(n_1971)
);

A2O1A1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1905),
.A2(n_1855),
.B(n_1836),
.C(n_1828),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1894),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1928),
.B(n_1882),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1941),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1937),
.Y(n_1976)
);

XNOR2xp5_ASAP7_75t_L g1977 ( 
.A(n_1939),
.B(n_1650),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1948),
.Y(n_1978)
);

AOI31xp33_ASAP7_75t_L g1979 ( 
.A1(n_1952),
.A2(n_1638),
.A3(n_1672),
.B(n_1650),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1968),
.B(n_1938),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1972),
.A2(n_1834),
.B1(n_1922),
.B2(n_1893),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1971),
.B(n_1890),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1941),
.Y(n_1983)
);

AOI222xp33_ASAP7_75t_L g1984 ( 
.A1(n_1939),
.A2(n_1853),
.B1(n_1851),
.B2(n_1833),
.C1(n_1893),
.C2(n_1924),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1948),
.A2(n_1892),
.B(n_1907),
.Y(n_1985)
);

AO22x1_ASAP7_75t_L g1986 ( 
.A1(n_1948),
.A2(n_1953),
.B1(n_1971),
.B2(n_1969),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1943),
.Y(n_1987)
);

O2A1O1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1965),
.A2(n_1908),
.B(n_1897),
.C(n_1926),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1948),
.A2(n_1853),
.B1(n_1840),
.B2(n_1841),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1965),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1943),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1940),
.B(n_1933),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1947),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1947),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1942),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1942),
.B(n_1935),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1946),
.B(n_1955),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1949),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1946),
.B(n_1917),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1936),
.B(n_1944),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1970),
.B(n_1934),
.C(n_1931),
.Y(n_2001)
);

AOI211xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1936),
.A2(n_1925),
.B(n_1866),
.C(n_1934),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1944),
.B(n_1925),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1949),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1975),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1976),
.B(n_2000),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1976),
.B(n_1672),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1977),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1984),
.A2(n_1977),
.B(n_1981),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1978),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1980),
.A2(n_1950),
.B1(n_1957),
.B2(n_1954),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_2000),
.B(n_1962),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_SL g2013 ( 
.A1(n_1985),
.A2(n_1945),
.B1(n_1961),
.B2(n_1954),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1979),
.A2(n_1899),
.B(n_1970),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1983),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1995),
.B(n_1712),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1978),
.Y(n_2017)
);

NAND3xp33_ASAP7_75t_SL g2018 ( 
.A(n_2002),
.B(n_1951),
.C(n_1962),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1997),
.B(n_1955),
.Y(n_2019)
);

OAI21xp33_ASAP7_75t_L g2020 ( 
.A1(n_1982),
.A2(n_2003),
.B(n_1992),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1987),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_2003),
.B(n_1966),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1996),
.B(n_1964),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1991),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1986),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1993),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2010),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2010),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_2009),
.A2(n_2001),
.B(n_1990),
.Y(n_2029)
);

AOI21xp33_ASAP7_75t_L g2030 ( 
.A1(n_2025),
.A2(n_2008),
.B(n_2006),
.Y(n_2030)
);

INVxp67_ASAP7_75t_SL g2031 ( 
.A(n_2007),
.Y(n_2031)
);

NOR3xp33_ASAP7_75t_L g2032 ( 
.A(n_2007),
.B(n_2025),
.C(n_2016),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2017),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_2016),
.B(n_1712),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2017),
.Y(n_2035)
);

NAND3xp33_ASAP7_75t_L g2036 ( 
.A(n_2013),
.B(n_1988),
.C(n_1994),
.Y(n_2036)
);

OAI32xp33_ASAP7_75t_L g2037 ( 
.A1(n_2019),
.A2(n_1998),
.A3(n_2004),
.B1(n_1999),
.B2(n_1960),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2022),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2022),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2012),
.B(n_1945),
.Y(n_2040)
);

NAND3xp33_ASAP7_75t_SL g2041 ( 
.A(n_2029),
.B(n_2011),
.C(n_2014),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2031),
.B(n_2020),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2038),
.B(n_2023),
.Y(n_2043)
);

OAI21xp33_ASAP7_75t_L g2044 ( 
.A1(n_2032),
.A2(n_2018),
.B(n_2015),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_2034),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2039),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2040),
.Y(n_2047)
);

NOR3xp33_ASAP7_75t_L g2048 ( 
.A(n_2030),
.B(n_2021),
.C(n_2005),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2027),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_2028),
.Y(n_2050)
);

OAI321xp33_ASAP7_75t_L g2051 ( 
.A1(n_2036),
.A2(n_2026),
.A3(n_2024),
.B1(n_1989),
.B2(n_1973),
.C(n_1967),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2033),
.B(n_1966),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_2034),
.B(n_2037),
.Y(n_2053)
);

O2A1O1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_2037),
.A2(n_2035),
.B(n_1960),
.C(n_1958),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2050),
.B(n_1961),
.Y(n_2055)
);

O2A1O1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_2051),
.A2(n_1958),
.B(n_1973),
.C(n_1967),
.Y(n_2056)
);

NAND4xp25_ASAP7_75t_L g2057 ( 
.A(n_2044),
.B(n_1950),
.C(n_1957),
.D(n_1967),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2041),
.A2(n_1973),
.B1(n_1959),
.B2(n_1957),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2052),
.Y(n_2059)
);

NOR4xp75_ASAP7_75t_SL g2060 ( 
.A(n_2043),
.B(n_1956),
.C(n_1974),
.D(n_1892),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2042),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2053),
.A2(n_1963),
.B(n_1959),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2045),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2063),
.A2(n_2045),
.B1(n_2048),
.B2(n_2049),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_L g2065 ( 
.A(n_2061),
.B(n_2046),
.C(n_2054),
.Y(n_2065)
);

AOI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2056),
.A2(n_2062),
.B1(n_2058),
.B2(n_2057),
.C(n_2055),
.Y(n_2066)
);

AOI321xp33_ASAP7_75t_L g2067 ( 
.A1(n_2059),
.A2(n_2047),
.A3(n_1959),
.B1(n_1963),
.B2(n_1957),
.C(n_1925),
.Y(n_2067)
);

AOI21xp33_ASAP7_75t_L g2068 ( 
.A1(n_2060),
.A2(n_1926),
.B(n_1875),
.Y(n_2068)
);

AOI21xp33_ASAP7_75t_SL g2069 ( 
.A1(n_2063),
.A2(n_1707),
.B(n_1926),
.Y(n_2069)
);

AOI221xp5_ASAP7_75t_L g2070 ( 
.A1(n_2056),
.A2(n_1931),
.B1(n_1924),
.B2(n_1916),
.C(n_1912),
.Y(n_2070)
);

NAND4xp25_ASAP7_75t_L g2071 ( 
.A(n_2055),
.B(n_1740),
.C(n_1866),
.D(n_1927),
.Y(n_2071)
);

NOR2xp67_ASAP7_75t_L g2072 ( 
.A(n_2064),
.B(n_2071),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_2067),
.Y(n_2073)
);

AND2x2_ASAP7_75t_SL g2074 ( 
.A(n_2065),
.B(n_1707),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2066),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2069),
.B(n_1707),
.Y(n_2076)
);

NOR4xp75_ASAP7_75t_L g2077 ( 
.A(n_2068),
.B(n_1866),
.C(n_1715),
.D(n_1776),
.Y(n_2077)
);

AOI221xp5_ASAP7_75t_L g2078 ( 
.A1(n_2073),
.A2(n_2075),
.B1(n_2076),
.B2(n_2070),
.C(n_2074),
.Y(n_2078)
);

OAI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2073),
.A2(n_1926),
.B1(n_1707),
.B2(n_1866),
.C(n_1916),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2072),
.B(n_1901),
.Y(n_2080)
);

NAND3xp33_ASAP7_75t_L g2081 ( 
.A(n_2077),
.B(n_1912),
.C(n_1904),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2080),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_2078),
.B(n_1894),
.Y(n_2083)
);

NAND4xp25_ASAP7_75t_L g2084 ( 
.A(n_2082),
.B(n_2079),
.C(n_2081),
.D(n_1676),
.Y(n_2084)
);

OAI22x1_ASAP7_75t_L g2085 ( 
.A1(n_2084),
.A2(n_2083),
.B1(n_1927),
.B2(n_1914),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2084),
.A2(n_1880),
.B1(n_1875),
.B2(n_1859),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2086),
.A2(n_1901),
.B1(n_1914),
.B2(n_1904),
.Y(n_2087)
);

OAI321xp33_ASAP7_75t_L g2088 ( 
.A1(n_2085),
.A2(n_1840),
.A3(n_1839),
.B1(n_1841),
.B2(n_1720),
.C(n_1875),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2087),
.B(n_1859),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2088),
.A2(n_1875),
.B1(n_1880),
.B2(n_1886),
.Y(n_2090)
);

OAI22x1_ASAP7_75t_L g2091 ( 
.A1(n_2089),
.A2(n_1757),
.B1(n_1782),
.B2(n_1879),
.Y(n_2091)
);

AOI22x1_ASAP7_75t_L g2092 ( 
.A1(n_2091),
.A2(n_2090),
.B1(n_1848),
.B2(n_1752),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_2092),
.A2(n_1880),
.B(n_1859),
.Y(n_2093)
);

OAI221xp5_ASAP7_75t_R g2094 ( 
.A1(n_2093),
.A2(n_1848),
.B1(n_1866),
.B2(n_1831),
.C(n_1860),
.Y(n_2094)
);

AOI211xp5_ASAP7_75t_L g2095 ( 
.A1(n_2094),
.A2(n_1711),
.B(n_1777),
.C(n_1709),
.Y(n_2095)
);


endmodule