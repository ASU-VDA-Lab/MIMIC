module real_jpeg_1112_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_286;
wire n_215;
wire n_249;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_238;
wire n_76;
wire n_79;
wire n_67;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_202;
wire n_244;
wire n_128;
wire n_295;
wire n_179;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_0),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_0),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_0),
.A2(n_29),
.B1(n_46),
.B2(n_50),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_2),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_2),
.A2(n_36),
.B1(n_38),
.B2(n_132),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_132),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_2),
.A2(n_46),
.B1(n_50),
.B2(n_132),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_3),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_3),
.A2(n_36),
.B1(n_38),
.B2(n_177),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_46),
.B1(n_50),
.B2(n_177),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_5),
.A2(n_36),
.B1(n_38),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_5),
.A2(n_46),
.B1(n_50),
.B2(n_61),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_7),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_7),
.A2(n_36),
.B1(n_38),
.B2(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_157),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_7),
.A2(n_46),
.B1(n_50),
.B2(n_157),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_9),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_9),
.A2(n_36),
.B1(n_38),
.B2(n_95),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_95),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_9),
.A2(n_46),
.B1(n_50),
.B2(n_95),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_26),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_10),
.A2(n_26),
.B(n_167),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_10),
.B(n_64),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_38),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_10),
.B(n_46),
.C(n_49),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_10),
.B(n_86),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_10),
.B(n_44),
.Y(n_258)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_13),
.A2(n_46),
.B1(n_50),
.B2(n_57),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_57),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_36),
.B1(n_38),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_14),
.A2(n_46),
.B1(n_50),
.B2(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_16),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_16),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_16),
.A2(n_40),
.B1(n_46),
.B2(n_50),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_21),
.B(n_96),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_79),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_22),
.A2(n_72),
.B1(n_73),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_22),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_23),
.A2(n_24),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_43),
.C(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_35),
.B2(n_39),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_25),
.A2(n_30),
.B1(n_35),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_27),
.A2(n_34),
.A3(n_38),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_30),
.A2(n_35),
.B1(n_39),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_30),
.A2(n_35),
.B1(n_94),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_30),
.A2(n_35),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_30),
.A2(n_35),
.B1(n_176),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_31),
.A2(n_131),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_33),
.B(n_36),
.Y(n_168)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_35),
.Y(n_158)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_38),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_36),
.B(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_38),
.A2(n_54),
.A3(n_65),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_58),
.B1(n_59),
.B2(n_71),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_71),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_51),
.B1(n_56),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_44),
.A2(n_51),
.B1(n_78),
.B2(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_44),
.A2(n_51),
.B1(n_91),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_44),
.A2(n_51),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_44),
.A2(n_51),
.B1(n_199),
.B2(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_44),
.A2(n_51),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_44),
.A2(n_51),
.B1(n_226),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_45),
.A2(n_125),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_45),
.A2(n_150),
.B1(n_198),
.B2(n_238),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_46),
.B(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_51),
.Y(n_150)
);

AO22x2_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_53),
.B(n_66),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_54),
.B(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_68),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_62),
.A2(n_64),
.B1(n_128),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_69),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_63),
.A2(n_76),
.B1(n_103),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_63),
.A2(n_103),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_63),
.A2(n_103),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_63),
.A2(n_103),
.B1(n_173),
.B2(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_63),
.A2(n_103),
.B1(n_188),
.B2(n_235),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_79),
.B(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_92),
.B(n_93),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_81),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_92),
.B1(n_93),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_83),
.A2(n_85),
.B1(n_121),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_83),
.A2(n_85),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_83),
.A2(n_85),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_84),
.A2(n_86),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_84),
.A2(n_86),
.B1(n_170),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_84),
.A2(n_86),
.B1(n_207),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_84),
.A2(n_86),
.B1(n_203),
.B2(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_84),
.A2(n_86),
.B1(n_256),
.B2(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_293),
.B(n_298),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_159),
.B(n_292),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_141),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_114),
.B(n_141),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_133),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_115),
.B(n_135),
.C(n_140),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_126),
.C(n_129),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_117),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_129),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.C(n_155),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_148),
.B(n_151),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_155),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_182),
.B(n_291),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_180),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_161),
.B(n_180),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_179),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_162),
.B(n_179),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_164),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_172),
.C(n_175),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_165),
.B(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_169),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_172),
.B(n_175),
.Y(n_282)
);

AOI31xp33_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_276),
.A3(n_285),
.B(n_288),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_221),
.B(n_275),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_209),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_185),
.B(n_209),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.C(n_200),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_186),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_191),
.C(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_196),
.B(n_200),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_209),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_209),
.B(n_286),
.Y(n_289)
);

FAx1_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.CI(n_212),
.CON(n_209),
.SN(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_213),
.B(n_216),
.C(n_220),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_270),
.B(n_274),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_239),
.B(n_269),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_231),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_228),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_234),
.C(n_237),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_250),
.B(n_268),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_262),
.B(n_267),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_257),
.B(n_261),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_259),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_266),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_273),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);


endmodule