module fake_jpeg_21540_n_84 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_32),
.B1(n_38),
.B2(n_31),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_49),
.B1(n_51),
.B2(n_4),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_33),
.B1(n_37),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_38),
.B1(n_17),
.B2(n_18),
.Y(n_51)
);

OR2x4_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_60),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_50),
.A3(n_49),
.B1(n_48),
.B2(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_27),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_58),
.B1(n_60),
.B2(n_5),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_68),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_72),
.B1(n_75),
.B2(n_68),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_76),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_71),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_9),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_14),
.B(n_15),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_19),
.B(n_22),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_24),
.Y(n_84)
);


endmodule