module fake_jpeg_31214_n_446 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_446);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_27),
.A2(n_18),
.B1(n_16),
.B2(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_72),
.Y(n_136)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_91),
.Y(n_94)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_89),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_18),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_99),
.A2(n_34),
.B1(n_38),
.B2(n_52),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_25),
.C(n_28),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_33),
.C(n_28),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_53),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_54),
.A2(n_23),
.B(n_25),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_40),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_34),
.Y(n_171)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_140),
.B(n_168),
.Y(n_192)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_24),
.B1(n_62),
.B2(n_56),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_145),
.B(n_165),
.Y(n_202)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_151),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_161),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_155),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_55),
.B1(n_63),
.B2(n_49),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_153),
.A2(n_156),
.B1(n_98),
.B2(n_96),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_24),
.B1(n_56),
.B2(n_61),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_163),
.B1(n_170),
.B2(n_172),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g155 ( 
.A(n_104),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_51),
.B1(n_64),
.B2(n_68),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_24),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_71),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_166),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_61),
.B1(n_72),
.B2(n_66),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_104),
.A2(n_59),
.B1(n_34),
.B2(n_38),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_91),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_94),
.B(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_93),
.A2(n_34),
.B1(n_38),
.B2(n_52),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_175),
.B1(n_114),
.B2(n_102),
.Y(n_193)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_191),
.B1(n_197),
.B2(n_198),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_16),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_140),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_136),
.B(n_124),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_165),
.B(n_171),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_96),
.B1(n_102),
.B2(n_114),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_85),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_107),
.B1(n_134),
.B2(n_118),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_144),
.A2(n_107),
.B1(n_76),
.B2(n_77),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g199 ( 
.A1(n_144),
.A2(n_98),
.B1(n_87),
.B2(n_80),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_50),
.B1(n_113),
.B2(n_132),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_180),
.B1(n_179),
.B2(n_197),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_211),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_199),
.B1(n_188),
.B2(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_218),
.B1(n_189),
.B2(n_193),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_222),
.B1(n_177),
.B2(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_150),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_182),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_182),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_166),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_176),
.B1(n_178),
.B2(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_178),
.A2(n_188),
.B1(n_183),
.B2(n_199),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_140),
.B(n_159),
.C(n_145),
.Y(n_220)
);

INVx3_ASAP7_75t_SL g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_155),
.B1(n_160),
.B2(n_113),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_230),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_147),
.C(n_149),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_226),
.C(n_195),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_152),
.C(n_158),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_139),
.B1(n_141),
.B2(n_146),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_199),
.A2(n_164),
.B1(n_175),
.B2(n_174),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_236),
.B1(n_245),
.B2(n_246),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_234),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_202),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_237),
.C(n_234),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_220),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_207),
.A2(n_195),
.B1(n_192),
.B2(n_198),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_195),
.B1(n_192),
.B2(n_186),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_198),
.B1(n_204),
.B2(n_179),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_253),
.B1(n_229),
.B2(n_193),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

OAI32xp33_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_209),
.A3(n_210),
.B1(n_214),
.B2(n_208),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_204),
.B1(n_193),
.B2(n_189),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_193),
.B1(n_184),
.B2(n_203),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_218),
.B1(n_217),
.B2(n_224),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_205),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_206),
.B(n_211),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_258),
.A2(n_286),
.B(n_129),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_225),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_136),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_243),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_261),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_230),
.B(n_226),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_266),
.B(n_277),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_218),
.B1(n_217),
.B2(n_224),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_217),
.B1(n_226),
.B2(n_219),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_231),
.A2(n_246),
.B(n_249),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_232),
.B(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_267),
.B(n_272),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_282),
.B1(n_285),
.B2(n_239),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_220),
.B1(n_227),
.B2(n_201),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_243),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_271),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_275),
.C(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_177),
.C(n_194),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_181),
.Y(n_277)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_279),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_148),
.A3(n_173),
.B1(n_227),
.B2(n_142),
.C1(n_151),
.C2(n_201),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_194),
.Y(n_280)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_267),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_151),
.B1(n_142),
.B2(n_168),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_187),
.B1(n_185),
.B2(n_129),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_239),
.B(n_185),
.Y(n_287)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_297),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_294),
.B1(n_296),
.B2(n_300),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_251),
.B(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_295),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_260),
.A2(n_242),
.B1(n_244),
.B2(n_187),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_242),
.B(n_157),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_187),
.B1(n_185),
.B2(n_157),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_305),
.C(n_315),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_260),
.A2(n_50),
.B1(n_128),
.B2(n_137),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_303),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_131),
.C(n_123),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_240),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_128),
.B1(n_1),
.B2(n_2),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_309),
.A2(n_274),
.B1(n_268),
.B2(n_284),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_311),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_264),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_312),
.A2(n_313),
.B1(n_271),
.B2(n_257),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_38),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_38),
.C(n_34),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_262),
.C(n_266),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_321),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_276),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_43),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_326),
.Y(n_346)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_333),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_265),
.C(n_272),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_339),
.C(n_299),
.Y(n_343)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_280),
.B1(n_286),
.B2(n_257),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_336),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_335),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_308),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_301),
.A2(n_279),
.B1(n_274),
.B2(n_287),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_338),
.A2(n_290),
.B1(n_295),
.B2(n_296),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_43),
.C(n_35),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_340),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_3),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_304),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_343),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_289),
.B(n_310),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_345),
.A2(n_330),
.B(n_333),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_315),
.C(n_316),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_358),
.C(n_364),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_352),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_338),
.A2(n_294),
.B1(n_310),
.B2(n_291),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_321),
.A2(n_291),
.B1(n_300),
.B2(n_309),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_329),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_313),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_359),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_312),
.C(n_292),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_43),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_363),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_362),
.A2(n_331),
.B1(n_324),
.B2(n_336),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_43),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_43),
.C(n_35),
.Y(n_364)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_368),
.Y(n_386)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_328),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_370),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_325),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_376),
.Y(n_396)
);

OAI21x1_ASAP7_75t_SL g372 ( 
.A1(n_356),
.A2(n_336),
.B(n_318),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_377),
.B(n_380),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_325),
.C(n_327),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_358),
.C(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_340),
.B1(n_329),
.B2(n_319),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_378),
.B(n_382),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_353),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_346),
.A2(n_341),
.B(n_339),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_337),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_357),
.A2(n_335),
.B(n_317),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_384),
.Y(n_397)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_387),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_370),
.B(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_388),
.B(n_371),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_343),
.C(n_347),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_399),
.C(n_393),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_365),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_393),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_359),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_369),
.B(n_377),
.Y(n_395)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_395),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_360),
.C(n_364),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_406),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_371),
.B1(n_383),
.B2(n_378),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_375),
.B(n_381),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_404),
.A2(n_405),
.B(n_408),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_397),
.A2(n_375),
.B(n_381),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_344),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_411),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_398),
.A2(n_366),
.B(n_363),
.Y(n_408)
);

AOI211xp5_ASAP7_75t_L g410 ( 
.A1(n_389),
.A2(n_362),
.B(n_5),
.C(n_6),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_410),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_4),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_4),
.B(n_5),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_412),
.A2(n_4),
.B(n_6),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_386),
.Y(n_413)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_390),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_417),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_399),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_35),
.C(n_11),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_400),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_420),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_35),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_423),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_422),
.A2(n_408),
.B(n_412),
.Y(n_427)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_418),
.A2(n_416),
.B(n_414),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_428),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_13),
.Y(n_436)
);

AOI21x1_ASAP7_75t_SL g431 ( 
.A1(n_418),
.A2(n_10),
.B(n_11),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_431),
.A2(n_432),
.B1(n_10),
.B2(n_13),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_436),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_424),
.A2(n_10),
.B(n_13),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_435),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_425),
.A2(n_426),
.B(n_432),
.Y(n_437)
);

AOI321xp33_ASAP7_75t_L g439 ( 
.A1(n_437),
.A2(n_14),
.A3(n_15),
.B1(n_35),
.B2(n_430),
.C(n_438),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_14),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_434),
.C(n_14),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_442),
.B(n_443),
.C(n_441),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_444),
.B(n_15),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_15),
.Y(n_446)
);


endmodule