module fake_netlist_6_2989_n_1716 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1716);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1716;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_28),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_35),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_47),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_108),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_62),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_77),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_18),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_45),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_19),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_80),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_34),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_29),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_48),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_100),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_75),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_38),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_48),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_61),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_105),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_68),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_112),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_140),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_142),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_45),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_57),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_49),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_95),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_5),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_41),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_51),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_34),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_23),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_83),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_26),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_126),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_154),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_17),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_0),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_79),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_26),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_13),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_86),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_87),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_23),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_29),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_66),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_127),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_39),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_4),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_44),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_113),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_125),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_40),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_20),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_33),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_88),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_47),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_40),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_150),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_21),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_38),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_133),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_114),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_43),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_134),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_19),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_93),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_22),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_41),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_22),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_73),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_53),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_72),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_54),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_81),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_10),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_3),
.Y(n_286)
);

BUFx2_ASAP7_75t_R g287 ( 
.A(n_60),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_25),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_106),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_56),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_17),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_14),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_145),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_74),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_31),
.Y(n_295)
);

BUFx2_ASAP7_75t_SL g296 ( 
.A(n_78),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_36),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_20),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_123),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_58),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_135),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_107),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_65),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_24),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_82),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_24),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_13),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_131),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_25),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_187),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_59),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_67),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_244),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_185),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_200),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_208),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_166),
.B(n_1),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_156),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_195),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_157),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_265),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_178),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_166),
.B(n_1),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_221),
.B(n_200),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_178),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_198),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_178),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_201),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_178),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_202),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_178),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_205),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_156),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_193),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_193),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_173),
.B(n_2),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_193),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_193),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_176),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_175),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_213),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_215),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_193),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_221),
.B(n_206),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_157),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_157),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_183),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_159),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_271),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_271),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_216),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_188),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_271),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_219),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_229),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_237),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_155),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_239),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_189),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_206),
.B(n_2),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_243),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_190),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_191),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_235),
.B(n_250),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_245),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_246),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_192),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_159),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_197),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_248),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_285),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_306),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_306),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_159),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_306),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_207),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_306),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_306),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_309),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_361),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_158),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_372),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_375),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_313),
.B(n_235),
.Y(n_406)
);

BUFx8_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_376),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_330),
.B(n_309),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_351),
.B(n_309),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_380),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_317),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_373),
.A2(n_222),
.B(n_171),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_382),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_389),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_313),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_316),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_332),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_314),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_309),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_312),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_334),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_334),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_336),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_314),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_336),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_R g438 ( 
.A(n_355),
.B(n_214),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_338),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_314),
.B(n_250),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_315),
.B(n_318),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_346),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_319),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_338),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_327),
.A2(n_311),
.B1(n_223),
.B2(n_231),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_348),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_342),
.B(n_217),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_348),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_431),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_325),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_349),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_423),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_429),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_349),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_429),
.B(n_387),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_429),
.B(n_165),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_418),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_360),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_429),
.B(n_423),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_429),
.B(n_423),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_442),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

BUFx4f_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_429),
.B(n_329),
.Y(n_486)
);

AO22x2_ASAP7_75t_L g487 ( 
.A1(n_406),
.A2(n_173),
.B1(n_276),
.B2(n_323),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_406),
.A2(n_309),
.B1(n_276),
.B2(n_222),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_391),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_424),
.B(n_360),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_443),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_423),
.B(n_363),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_414),
.B(n_425),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_390),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_406),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_392),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_392),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_392),
.B(n_321),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_441),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_432),
.B(n_363),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_418),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_406),
.B(n_440),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_444),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_406),
.B(n_264),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_347),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_431),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_458),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_440),
.B(n_436),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_454),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_458),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_436),
.B(n_365),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_444),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_459),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_440),
.B(n_264),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_345),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_446),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_440),
.B(n_365),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_440),
.B(n_284),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_430),
.B(n_284),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_411),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_454),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_430),
.B(n_301),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_410),
.B(n_367),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

INVx4_ASAP7_75t_SL g545 ( 
.A(n_454),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_419),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_399),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_410),
.B(n_322),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_412),
.B(n_367),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_412),
.B(n_369),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_434),
.B(n_369),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_409),
.B(n_374),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_437),
.A2(n_374),
.B1(n_378),
.B2(n_379),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_439),
.B(n_378),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_413),
.B(n_301),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_409),
.B(n_379),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_438),
.B(n_302),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_419),
.A2(n_240),
.B1(n_210),
.B2(n_266),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_449),
.B(n_383),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_409),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_419),
.B(n_368),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_409),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_419),
.B(n_326),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_462),
.B(n_383),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_453),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_409),
.B(n_326),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_459),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_454),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_398),
.A2(n_212),
.B1(n_303),
.B2(n_258),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_404),
.B(n_352),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_413),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_404),
.A2(n_211),
.B1(n_160),
.B2(n_174),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_405),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_438),
.B(n_302),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_405),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_400),
.B(n_161),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_460),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_402),
.B(n_353),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_460),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_413),
.B(n_203),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_451),
.B(n_255),
.C(n_253),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_402),
.B(n_381),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_448),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_416),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_415),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_460),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_402),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_415),
.A2(n_251),
.B1(n_238),
.B2(n_236),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_416),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_416),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_448),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_400),
.B(n_218),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_443),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_447),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_448),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_543),
.B(n_551),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_501),
.B(n_452),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_503),
.B(n_452),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_471),
.A2(n_428),
.B1(n_407),
.B2(n_220),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_484),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_549),
.B(n_428),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_502),
.B(n_452),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_484),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_475),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_513),
.A2(n_428),
.B1(n_261),
.B2(n_164),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_483),
.B(n_452),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_513),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_552),
.B(n_397),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_468),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_403),
.C(n_401),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_496),
.B(n_162),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_525),
.Y(n_625)
);

NOR3xp33_ASAP7_75t_L g626 ( 
.A(n_466),
.B(n_417),
.C(n_408),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_500),
.B(n_172),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_476),
.A2(n_407),
.B1(n_225),
.B2(n_226),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_490),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_493),
.B(n_420),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_495),
.B(n_287),
.Y(n_631)
);

AO22x1_ASAP7_75t_L g632 ( 
.A1(n_568),
.A2(n_407),
.B1(n_249),
.B2(n_242),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_486),
.B(n_568),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_565),
.B(n_186),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_422),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_519),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_549),
.B(n_394),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_536),
.A2(n_407),
.B1(n_247),
.B2(n_228),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_492),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_549),
.B(n_394),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_463),
.B(n_394),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_555),
.B(n_407),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_565),
.A2(n_296),
.B1(n_199),
.B2(n_230),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_204),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_523),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_578),
.B(n_163),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_578),
.B(n_163),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_475),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_491),
.B(n_447),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_481),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_540),
.A2(n_184),
.B1(n_288),
.B2(n_263),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_481),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_478),
.A2(n_421),
.B(n_396),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_562),
.A2(n_267),
.B1(n_227),
.B2(n_224),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_522),
.B(n_209),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_473),
.B(n_257),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_473),
.B(n_268),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_596),
.B(n_167),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_596),
.B(n_523),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_479),
.B(n_421),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_499),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_499),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_482),
.B(n_421),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_507),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_539),
.A2(n_272),
.B1(n_196),
.B2(n_252),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_472),
.A2(n_289),
.B1(n_180),
.B2(n_310),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_510),
.B(n_455),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_583),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_275),
.C(n_279),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_542),
.A2(n_286),
.B1(n_291),
.B2(n_292),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_504),
.B(n_396),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_540),
.B(n_396),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_507),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_505),
.B(n_396),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_523),
.B(n_167),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_523),
.B(n_233),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_554),
.B(n_168),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_556),
.B(n_455),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_518),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_518),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_558),
.B(n_168),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_520),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_563),
.B(n_169),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_560),
.B(n_169),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_520),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_569),
.B(n_274),
.C(n_262),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_516),
.B(n_170),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_516),
.A2(n_295),
.B1(n_179),
.B2(n_277),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_530),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_521),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_590),
.B(n_256),
.C(n_259),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_468),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_581),
.B(n_584),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_560),
.B(n_170),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_517),
.Y(n_698)
);

NOR2x1p5_ASAP7_75t_L g699 ( 
.A(n_587),
.B(n_498),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_521),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_582),
.B(n_180),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_527),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_515),
.A2(n_278),
.B1(n_280),
.B2(n_305),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_594),
.B(n_181),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_582),
.B(n_181),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_515),
.A2(n_269),
.B1(n_254),
.B2(n_194),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_531),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_506),
.B(n_182),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_587),
.B(n_182),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_498),
.B(n_234),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_477),
.B(n_234),
.Y(n_712)
);

NAND2x1_ASAP7_75t_L g713 ( 
.A(n_497),
.B(n_117),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_477),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_519),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_509),
.B(n_310),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_531),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_544),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_583),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_307),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_544),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_SL g722 ( 
.A(n_488),
.B(n_175),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_602),
.B(n_307),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_529),
.B(n_305),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_532),
.B(n_304),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_533),
.A2(n_217),
.B1(n_177),
.B2(n_299),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_535),
.B(n_304),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_571),
.B(n_289),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_550),
.B(n_559),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_R g730 ( 
.A1(n_605),
.A2(n_177),
.B1(n_232),
.B2(n_281),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_570),
.B(n_300),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_485),
.A2(n_217),
.B(n_300),
.C(n_283),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_606),
.B(n_290),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_573),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_572),
.B(n_299),
.Y(n_735)
);

OAI221xp5_ASAP7_75t_L g736 ( 
.A1(n_577),
.A2(n_260),
.B1(n_297),
.B2(n_298),
.C(n_281),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_485),
.A2(n_290),
.B1(n_282),
.B2(n_294),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_574),
.B(n_294),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_589),
.A2(n_298),
.B1(n_297),
.B2(n_232),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_576),
.B(n_293),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_600),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_573),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_586),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_586),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_547),
.A2(n_293),
.B1(n_283),
.B2(n_282),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_547),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_588),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_547),
.B(n_3),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_603),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_588),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_593),
.B(n_69),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_538),
.B(n_84),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_517),
.B(n_55),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_517),
.B(n_85),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_534),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_595),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_606),
.B(n_52),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_487),
.A2(n_89),
.B1(n_153),
.B2(n_149),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_595),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_526),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_526),
.B(n_147),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_564),
.B(n_143),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_564),
.B(n_139),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_495),
.B(n_6),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_564),
.B(n_136),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_607),
.A2(n_604),
.B(n_585),
.C(n_599),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_611),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_615),
.B(n_495),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_671),
.B(n_534),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_639),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_645),
.A2(n_512),
.B(n_497),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_619),
.B(n_548),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_645),
.A2(n_512),
.B(n_524),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_645),
.A2(n_524),
.B(n_561),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_612),
.B(n_546),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_622),
.B(n_487),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_713),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_633),
.A2(n_464),
.B(n_474),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_611),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_671),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_614),
.B(n_548),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_SL g783 ( 
.A(n_631),
.B(n_583),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_620),
.B(n_546),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_634),
.A2(n_464),
.B(n_511),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_723),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_SL g787 ( 
.A1(n_752),
.A2(n_601),
.B(n_464),
.C(n_470),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_616),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_614),
.B(n_619),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_641),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_686),
.B(n_546),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_674),
.A2(n_575),
.B(n_567),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_748),
.A2(n_630),
.B1(n_657),
.B2(n_635),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_694),
.B(n_691),
.C(n_764),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_677),
.A2(n_575),
.B(n_557),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_621),
.B(n_548),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_675),
.B(n_465),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_663),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_714),
.B(n_690),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_675),
.B(n_585),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_701),
.A2(n_585),
.B(n_598),
.C(n_579),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_613),
.A2(n_609),
.B(n_608),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_625),
.B(n_597),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_621),
.B(n_537),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_610),
.B(n_537),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_637),
.B(n_537),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_650),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_637),
.B(n_537),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_719),
.Y(n_809)
);

INVx11_ASAP7_75t_L g810 ( 
.A(n_719),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_711),
.A2(n_598),
.B(n_579),
.C(n_580),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_640),
.B(n_548),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_636),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_643),
.A2(n_746),
.B1(n_654),
.B2(n_656),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_698),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_640),
.B(n_566),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_663),
.B(n_566),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_658),
.A2(n_566),
.B1(n_530),
.B2(n_579),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_746),
.A2(n_679),
.B(n_618),
.Y(n_819)
);

BUFx12f_ASAP7_75t_L g820 ( 
.A(n_715),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_712),
.B(n_566),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_666),
.B(n_530),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_699),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_666),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_751),
.A2(n_511),
.B(n_530),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_648),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_L g827 ( 
.A1(n_710),
.A2(n_735),
.B(n_736),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_696),
.B(n_606),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_646),
.B(n_606),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_698),
.A2(n_606),
.B1(n_592),
.B2(n_541),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_735),
.B(n_649),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_650),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_729),
.A2(n_541),
.B(n_592),
.Y(n_833)
);

AOI21x1_ASAP7_75t_L g834 ( 
.A1(n_644),
.A2(n_545),
.B(n_592),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_692),
.A2(n_541),
.B(n_592),
.Y(n_835)
);

OAI321xp33_ASAP7_75t_L g836 ( 
.A1(n_739),
.A2(n_651),
.A3(n_617),
.B1(n_726),
.B2(n_642),
.C(n_628),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_659),
.A2(n_684),
.B1(n_680),
.B2(n_661),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_722),
.A2(n_545),
.B1(n_7),
.B2(n_8),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_692),
.A2(n_545),
.B(n_130),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_698),
.A2(n_545),
.B(n_124),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_667),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_760),
.A2(n_627),
.B(n_624),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_741),
.B(n_6),
.Y(n_843)
);

CKINVDCx10_ASAP7_75t_R g844 ( 
.A(n_636),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_667),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_638),
.B(n_119),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_749),
.B(n_8),
.Y(n_847)
);

CKINVDCx11_ASAP7_75t_R g848 ( 
.A(n_715),
.Y(n_848)
);

BUFx8_ASAP7_75t_SL g849 ( 
.A(n_709),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_737),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_760),
.B(n_118),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_670),
.B(n_11),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_681),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_722),
.A2(n_16),
.B1(n_30),
.B2(n_32),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_730),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_705),
.A2(n_103),
.B1(n_99),
.B2(n_96),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_745),
.A2(n_37),
.B(n_42),
.C(n_43),
.Y(n_857)
);

CKINVDCx6p67_ASAP7_75t_R g858 ( 
.A(n_647),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_SL g859 ( 
.A(n_660),
.B(n_44),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_682),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_672),
.B(n_46),
.C(n_50),
.Y(n_861)
);

AO32x2_ASAP7_75t_L g862 ( 
.A1(n_669),
.A2(n_50),
.A3(n_51),
.B1(n_732),
.B2(n_632),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_716),
.Y(n_863)
);

BUFx4f_ASAP7_75t_L g864 ( 
.A(n_682),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_753),
.A2(n_765),
.B(n_763),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_724),
.B(n_740),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_689),
.B(n_623),
.Y(n_867)
);

BUFx4f_ASAP7_75t_L g868 ( 
.A(n_683),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_683),
.A2(n_734),
.B(n_721),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_727),
.B(n_721),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_754),
.A2(n_762),
.B(n_761),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_720),
.A2(n_731),
.B1(n_725),
.B2(n_738),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_SL g873 ( 
.A(n_758),
.B(n_626),
.C(n_673),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_653),
.A2(n_706),
.B(n_687),
.C(n_697),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_685),
.B(n_734),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_713),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_755),
.B(n_668),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_757),
.B(n_733),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_685),
.A2(n_718),
.B(n_717),
.C(n_688),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_728),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_707),
.A2(n_703),
.B1(n_717),
.B2(n_718),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_688),
.A2(n_708),
.B(n_652),
.C(n_655),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_678),
.B(n_632),
.C(n_733),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_759),
.A2(n_662),
.B1(n_664),
.B2(n_665),
.Y(n_884)
);

AO21x1_ASAP7_75t_L g885 ( 
.A1(n_757),
.A2(n_676),
.B(n_693),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_700),
.B(n_702),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_702),
.B(n_704),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_704),
.A2(n_708),
.B1(n_759),
.B2(n_742),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_742),
.A2(n_743),
.B1(n_744),
.B2(n_747),
.Y(n_889)
);

AOI21x1_ASAP7_75t_L g890 ( 
.A1(n_743),
.A2(n_744),
.B(n_747),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_750),
.A2(n_756),
.B(n_755),
.Y(n_891)
);

AOI22x1_ASAP7_75t_L g892 ( 
.A1(n_629),
.A2(n_622),
.B1(n_695),
.B2(n_619),
.Y(n_892)
);

NAND2x1_ASAP7_75t_L g893 ( 
.A(n_692),
.B(n_469),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_607),
.B(n_629),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_611),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_633),
.A2(n_547),
.B(n_485),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_715),
.B(n_395),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_622),
.A2(n_695),
.B1(n_619),
.B2(n_633),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_645),
.A2(n_469),
.B(n_513),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_622),
.A2(n_695),
.B1(n_619),
.B2(n_633),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_607),
.B(n_629),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_698),
.A2(n_480),
.B(n_478),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_607),
.A2(n_619),
.B1(n_695),
.B2(n_622),
.Y(n_903)
);

AOI22x1_ASAP7_75t_L g904 ( 
.A1(n_629),
.A2(n_622),
.B1(n_695),
.B2(n_619),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_607),
.A2(n_619),
.B(n_629),
.C(n_701),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_629),
.A2(n_607),
.B(n_633),
.C(n_634),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_633),
.A2(n_547),
.B(n_485),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_645),
.A2(n_469),
.B(n_513),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_611),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_629),
.A2(n_607),
.B(n_633),
.C(n_634),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_607),
.A2(n_619),
.B(n_629),
.C(n_701),
.Y(n_911)
);

BUFx12f_ASAP7_75t_L g912 ( 
.A(n_671),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_607),
.B(n_629),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_645),
.A2(n_469),
.B(n_513),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_645),
.A2(n_469),
.B(n_513),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_634),
.A2(n_513),
.B(n_490),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_645),
.A2(n_469),
.B(n_513),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_611),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_645),
.A2(n_469),
.B(n_513),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_622),
.A2(n_695),
.B1(n_619),
.B2(n_633),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_615),
.B(n_607),
.Y(n_921)
);

O2A1O1Ixp5_ASAP7_75t_L g922 ( 
.A1(n_607),
.A2(n_486),
.B(n_542),
.C(n_539),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_SL g923 ( 
.A1(n_752),
.A2(n_633),
.B(n_634),
.C(n_753),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_622),
.A2(n_695),
.B1(n_619),
.B2(n_633),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_607),
.B(n_615),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_607),
.B(n_629),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_607),
.B(n_615),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_L g928 ( 
.A1(n_607),
.A2(n_486),
.B(n_542),
.C(n_539),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_633),
.A2(n_547),
.B(n_485),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_645),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_713),
.B(n_513),
.Y(n_931)
);

AOI33xp33_ASAP7_75t_L g932 ( 
.A1(n_691),
.A2(n_451),
.A3(n_651),
.B1(n_457),
.B2(n_596),
.B3(n_288),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_607),
.B(n_629),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_930),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_930),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_923),
.A2(n_900),
.B(n_898),
.Y(n_936)
);

OAI22x1_ASAP7_75t_L g937 ( 
.A1(n_921),
.A2(n_784),
.B1(n_793),
.B2(n_791),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_920),
.A2(n_924),
.B(n_907),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_933),
.B(n_894),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_SL g940 ( 
.A1(n_901),
.A2(n_926),
.B(n_913),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_831),
.A2(n_921),
.B1(n_866),
.B2(n_863),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_SL g942 ( 
.A1(n_906),
.A2(n_910),
.B(n_896),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_883),
.A2(n_777),
.B(n_846),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_792),
.A2(n_834),
.B(n_795),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_930),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_929),
.A2(n_911),
.B(n_905),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_770),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_813),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_860),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_903),
.B(n_925),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_860),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_802),
.A2(n_875),
.B(n_871),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_883),
.A2(n_857),
.B(n_850),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_826),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_791),
.A2(n_827),
.B(n_786),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_842),
.A2(n_779),
.B(n_785),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_927),
.B(n_798),
.Y(n_957)
);

NAND2x1_ASAP7_75t_L g958 ( 
.A(n_930),
.B(n_815),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_922),
.A2(n_928),
.B(n_814),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_817),
.A2(n_822),
.B(n_828),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_844),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_878),
.A2(n_808),
.B(n_816),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_807),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_878),
.A2(n_806),
.B(n_812),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_772),
.B(n_799),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_897),
.Y(n_966)
);

INVx5_ASAP7_75t_L g967 ( 
.A(n_778),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_773),
.A2(n_892),
.B(n_904),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_771),
.A2(n_774),
.B(n_775),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_L g970 ( 
.A1(n_855),
.A2(n_836),
.B1(n_854),
.B2(n_794),
.C(n_873),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_832),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_823),
.Y(n_972)
);

OAI22x1_ASAP7_75t_L g973 ( 
.A1(n_786),
.A2(n_852),
.B1(n_768),
.B2(n_799),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_824),
.B(n_790),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_931),
.A2(n_914),
.B(n_908),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_931),
.A2(n_899),
.B(n_919),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_915),
.A2(n_917),
.B(n_888),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_815),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_772),
.B(n_870),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_841),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_767),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_801),
.A2(n_865),
.B(n_869),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_838),
.A2(n_794),
.B(n_854),
.C(n_932),
.Y(n_983)
);

OAI22x1_ASAP7_75t_L g984 ( 
.A1(n_768),
.A2(n_776),
.B1(n_797),
.B2(n_823),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_922),
.A2(n_928),
.B(n_766),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_789),
.B(n_821),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_889),
.A2(n_893),
.B(n_887),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_803),
.B(n_877),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_848),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_891),
.A2(n_874),
.B(n_879),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_821),
.B(n_872),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_809),
.B(n_880),
.Y(n_992)
);

OAI21x1_ASAP7_75t_SL g993 ( 
.A1(n_885),
.A2(n_838),
.B(n_839),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_845),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_855),
.A2(n_859),
.B(n_861),
.C(n_776),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_780),
.B(n_895),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_864),
.B(n_868),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_909),
.B(n_918),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_796),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_835),
.A2(n_782),
.B(n_833),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_811),
.A2(n_800),
.B(n_882),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_864),
.B(n_868),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_820),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_858),
.B(n_853),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_884),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_787),
.A2(n_881),
.B(n_778),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_830),
.A2(n_840),
.B(n_804),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_818),
.A2(n_886),
.B(n_805),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_778),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_867),
.B(n_873),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_837),
.B(n_829),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_912),
.Y(n_1012)
);

BUFx4f_ASAP7_75t_L g1013 ( 
.A(n_851),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_851),
.Y(n_1014)
);

AO21x2_ASAP7_75t_L g1015 ( 
.A1(n_829),
.A2(n_843),
.B(n_847),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_778),
.A2(n_876),
.B(n_856),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_862),
.A2(n_769),
.B(n_810),
.Y(n_1017)
);

AO31x2_ASAP7_75t_L g1018 ( 
.A1(n_862),
.A2(n_783),
.A3(n_849),
.B(n_781),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_862),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_862),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_894),
.B(n_901),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_793),
.B(n_894),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_770),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_770),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_894),
.A2(n_901),
.B1(n_926),
.B2(n_913),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_860),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_860),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_831),
.B(n_921),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_890),
.A2(n_819),
.B(n_916),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_788),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_770),
.B(n_671),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_894),
.B(n_901),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_770),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_813),
.B(n_639),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_770),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_930),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_R g1043 ( 
.A(n_912),
.B(n_671),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_793),
.B(n_894),
.Y(n_1044)
);

AO21x2_ASAP7_75t_L g1045 ( 
.A1(n_779),
.A2(n_907),
.B(n_896),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_831),
.A2(n_793),
.B1(n_607),
.B2(n_921),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_894),
.B(n_901),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_SL g1048 ( 
.A(n_783),
.B(n_395),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_894),
.B(n_901),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_860),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_902),
.A2(n_890),
.B(n_825),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_902),
.A2(n_890),
.B(n_825),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_813),
.B(n_639),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_831),
.A2(n_793),
.B1(n_607),
.B2(n_921),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_902),
.A2(n_890),
.B(n_825),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_902),
.A2(n_890),
.B(n_825),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_894),
.B(n_901),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_894),
.A2(n_901),
.B(n_926),
.C(n_913),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_905),
.A2(n_911),
.B(n_922),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_894),
.B(n_901),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_894),
.B(n_901),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_923),
.A2(n_633),
.B(n_898),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_954),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_947),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_934),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1024),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_982),
.A2(n_956),
.B(n_942),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_934),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1020),
.A2(n_970),
.B1(n_1066),
.B2(n_1065),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_980),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1010),
.A2(n_970),
.B1(n_937),
.B2(n_988),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_994),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_1025),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1063),
.B(n_1026),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1010),
.A2(n_1048),
.B1(n_1029),
.B2(n_1056),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1039),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_938),
.A2(n_991),
.B(n_968),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_934),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1038),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_L g1085 ( 
.A(n_955),
.B(n_1046),
.C(n_995),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_983),
.A2(n_1063),
.B(n_995),
.C(n_940),
.Y(n_1086)
);

CKINVDCx8_ASAP7_75t_R g1087 ( 
.A(n_989),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_941),
.B(n_1021),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_949),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_985),
.A2(n_1064),
.B(n_1006),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_951),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_1036),
.Y(n_1092)
);

BUFx10_ASAP7_75t_L g1093 ( 
.A(n_961),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_963),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_1023),
.A2(n_1044),
.B(n_1011),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_938),
.A2(n_1016),
.B(n_1067),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1055),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1034),
.B(n_1047),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_L g1099 ( 
.A(n_983),
.B(n_1023),
.C(n_1044),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1006),
.A2(n_1067),
.B(n_1042),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_948),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_939),
.C(n_950),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1022),
.A2(n_1035),
.B(n_1061),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_1014),
.B(n_934),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_939),
.B(n_965),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1004),
.B(n_979),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1022),
.A2(n_1040),
.B(n_1060),
.Y(n_1107)
);

NOR2x1p5_ASAP7_75t_L g1108 ( 
.A(n_1003),
.B(n_1012),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_992),
.B(n_1014),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_SL g1110 ( 
.A1(n_1020),
.A2(n_1013),
.B1(n_1003),
.B2(n_1017),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1027),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_986),
.B(n_999),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1028),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_971),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_992),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_972),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_1050),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_945),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1032),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_962),
.B(n_964),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1013),
.B(n_957),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_962),
.B(n_964),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_960),
.B(n_1005),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_966),
.A2(n_1019),
.B1(n_1033),
.B2(n_993),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_981),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_981),
.B(n_973),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_974),
.B(n_997),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_960),
.B(n_1015),
.Y(n_1128)
);

CKINVDCx8_ASAP7_75t_R g1129 ( 
.A(n_1033),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_984),
.B(n_1018),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_967),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1033),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_1012),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_996),
.Y(n_1134)
);

INVx3_ASAP7_75t_SL g1135 ( 
.A(n_945),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_SL g1136 ( 
.A(n_967),
.B(n_1009),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1018),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1018),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1015),
.B(n_943),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_935),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_935),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_959),
.A2(n_997),
.B(n_1002),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_967),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1030),
.A2(n_1040),
.B(n_1053),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_998),
.B(n_1002),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_L g1146 ( 
.A(n_1009),
.B(n_1041),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1041),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1018),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_978),
.B(n_958),
.Y(n_1149)
);

INVx8_ASAP7_75t_L g1150 ( 
.A(n_1009),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_L g1151 ( 
.A(n_1009),
.B(n_978),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_953),
.B(n_1019),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1019),
.A2(n_990),
.B1(n_1001),
.B2(n_1043),
.Y(n_1153)
);

INVx3_ASAP7_75t_SL g1154 ( 
.A(n_1019),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1031),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1008),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_946),
.B(n_1045),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_975),
.B(n_976),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_936),
.A2(n_1060),
.B(n_1058),
.C(n_1053),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_936),
.B(n_1058),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1007),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1035),
.B(n_1051),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_SL g1163 ( 
.A(n_1045),
.B(n_952),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_987),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_969),
.B(n_977),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1000),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1037),
.B(n_1051),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_1042),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1052),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1054),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_944),
.B(n_1057),
.C(n_1059),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_954),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_992),
.B(n_772),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1063),
.B(n_894),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_947),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1029),
.B(n_831),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1010),
.A2(n_853),
.B1(n_670),
.B2(n_681),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_954),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_983),
.A2(n_970),
.B(n_1063),
.C(n_911),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1029),
.B(n_831),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_954),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_947),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_954),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_1038),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_947),
.Y(n_1185)
);

OR2x6_ASAP7_75t_L g1186 ( 
.A(n_1033),
.B(n_997),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1029),
.B(n_831),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_982),
.A2(n_469),
.B(n_645),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_982),
.A2(n_469),
.B(n_645),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_954),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1029),
.B(n_831),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_947),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_1048),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1013),
.B(n_631),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1038),
.Y(n_1195)
);

AO21x1_ASAP7_75t_L g1196 ( 
.A1(n_1010),
.A2(n_991),
.B(n_1023),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1029),
.B(n_831),
.Y(n_1197)
);

BUFx10_ASAP7_75t_L g1198 ( 
.A(n_961),
.Y(n_1198)
);

BUFx4_ASAP7_75t_SL g1199 ( 
.A(n_1012),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_947),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1199),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1123),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1085),
.A2(n_1177),
.B1(n_1076),
.B2(n_1153),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1075),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1087),
.B(n_1193),
.Y(n_1205)
);

AO21x2_ASAP7_75t_L g1206 ( 
.A1(n_1144),
.A2(n_1107),
.B(n_1103),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1150),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1077),
.Y(n_1208)
);

BUFx10_ASAP7_75t_L g1209 ( 
.A(n_1108),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1172),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1085),
.A2(n_1153),
.B1(n_1074),
.B2(n_1099),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1074),
.A2(n_1099),
.B1(n_1196),
.B2(n_1088),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1096),
.B(n_1072),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1178),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1150),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1159),
.A2(n_1162),
.B(n_1082),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1181),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1183),
.Y(n_1218)
);

BUFx12f_ASAP7_75t_L g1219 ( 
.A(n_1093),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1190),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1080),
.A2(n_1180),
.B1(n_1197),
.B2(n_1187),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1194),
.A2(n_1106),
.B1(n_1191),
.B2(n_1176),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1200),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1194),
.A2(n_1098),
.B1(n_1127),
.B2(n_1079),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1134),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1101),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1101),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1168),
.B(n_1136),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1102),
.A2(n_1174),
.B(n_1098),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1157),
.B(n_1120),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_1090),
.B(n_1167),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1069),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1139),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1185),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1093),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1089),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1150),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1174),
.A2(n_1086),
.B(n_1142),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1091),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1084),
.A2(n_1195),
.B1(n_1186),
.B2(n_1112),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1112),
.B(n_1105),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1126),
.A2(n_1195),
.B1(n_1084),
.B2(n_1148),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1111),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1113),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1125),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1121),
.A2(n_1097),
.B1(n_1184),
.B2(n_1105),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1152),
.B(n_1130),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1094),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1198),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1137),
.A2(n_1138),
.B1(n_1186),
.B2(n_1090),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1083),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1114),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1156),
.B(n_1160),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1119),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1198),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1095),
.A2(n_1142),
.B1(n_1110),
.B2(n_1124),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1117),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1173),
.A2(n_1186),
.B1(n_1109),
.B2(n_1145),
.Y(n_1258)
);

AND2x4_ASAP7_75t_SL g1259 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1117),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1133),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1083),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1070),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1154),
.B(n_1122),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1070),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1120),
.B(n_1122),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1109),
.B(n_1128),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1070),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1083),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1173),
.A2(n_1175),
.B1(n_1071),
.B2(n_1116),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1092),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1073),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1170),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1132),
.A2(n_1192),
.B1(n_1182),
.B2(n_1115),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1129),
.A2(n_1147),
.B1(n_1078),
.B2(n_1081),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1135),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1149),
.B(n_1131),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1140),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1156),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1179),
.A2(n_1104),
.B1(n_1146),
.B2(n_1151),
.Y(n_1280)
);

NOR2x1_ASAP7_75t_R g1281 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1104),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1131),
.B(n_1143),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1104),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1118),
.A2(n_1165),
.B1(n_1158),
.B2(n_1161),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1165),
.A2(n_1164),
.B1(n_1166),
.B2(n_1188),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1163),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1169),
.Y(n_1288)
);

CKINVDCx6p67_ASAP7_75t_R g1289 ( 
.A(n_1189),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1171),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1171),
.Y(n_1291)
);

NOR2x1_ASAP7_75t_SL g1292 ( 
.A(n_1168),
.B(n_967),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1087),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1194),
.A2(n_784),
.B1(n_631),
.B2(n_783),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1085),
.A2(n_1010),
.B1(n_970),
.B2(n_794),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1154),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1076),
.B(n_1010),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1068),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1085),
.A2(n_1010),
.B1(n_970),
.B2(n_794),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1144),
.A2(n_1107),
.B(n_1103),
.Y(n_1300)
);

AO21x1_ASAP7_75t_SL g1301 ( 
.A1(n_1079),
.A2(n_1139),
.B(n_1174),
.Y(n_1301)
);

BUFx10_ASAP7_75t_L g1302 ( 
.A(n_1108),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1200),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1076),
.B(n_1010),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1068),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1200),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1144),
.A2(n_1159),
.B(n_1100),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1199),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1068),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1068),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_1098),
.B1(n_1046),
.B2(n_1056),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1155),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1226),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1247),
.B(n_1267),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1295),
.A2(n_1299),
.B(n_1212),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1205),
.B(n_1232),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1227),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1247),
.B(n_1267),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1257),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1230),
.B(n_1266),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1266),
.B(n_1241),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1260),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1230),
.B(n_1297),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1296),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1264),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1297),
.B(n_1304),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1234),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1307),
.A2(n_1290),
.B(n_1253),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1307),
.A2(n_1253),
.B(n_1286),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1229),
.A2(n_1238),
.B(n_1233),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1253),
.A2(n_1287),
.B(n_1216),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1304),
.B(n_1264),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1277),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1211),
.A2(n_1256),
.B(n_1291),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1301),
.B(n_1231),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1245),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1202),
.B(n_1288),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1277),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1291),
.A2(n_1202),
.B(n_1312),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1225),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1216),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1296),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1225),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1231),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1206),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1300),
.Y(n_1346)
);

INVx5_ASAP7_75t_SL g1347 ( 
.A(n_1213),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1246),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1279),
.B(n_1285),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1213),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1294),
.B(n_1271),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1213),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1214),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1213),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1220),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1224),
.B(n_1311),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1220),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1273),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1208),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1210),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1217),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1218),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1292),
.A2(n_1228),
.B(n_1280),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1204),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1204),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1240),
.B(n_1273),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1236),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1239),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1223),
.B(n_1303),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1243),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1293),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1203),
.B(n_1242),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1244),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1289),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1310),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1293),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1301),
.B(n_1250),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1289),
.Y(n_1378)
);

INVxp33_ASAP7_75t_L g1379 ( 
.A(n_1275),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1298),
.A2(n_1309),
.B(n_1305),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1255),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1221),
.B(n_1222),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1335),
.B(n_1320),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1329),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1339),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1348),
.B(n_1258),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1339),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1335),
.B(n_1254),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1378),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1329),
.Y(n_1390)
);

AOI221xp5_ASAP7_75t_L g1391 ( 
.A1(n_1315),
.A2(n_1274),
.B1(n_1270),
.B2(n_1254),
.C(n_1252),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1320),
.B(n_1248),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1378),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1341),
.B(n_1344),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1321),
.B(n_1323),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1323),
.B(n_1268),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1350),
.B(n_1263),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1350),
.B(n_1265),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1350),
.B(n_1272),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1328),
.B(n_1352),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1321),
.B(n_1284),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_1330),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1352),
.B(n_1282),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1352),
.B(n_1207),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1354),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1315),
.A2(n_1278),
.B1(n_1255),
.B2(n_1276),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1326),
.B(n_1283),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1378),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1356),
.A2(n_1334),
.B1(n_1372),
.B2(n_1379),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1330),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1326),
.B(n_1269),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1330),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1314),
.B(n_1251),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1345),
.B(n_1276),
.Y(n_1414)
);

OAI211xp5_ASAP7_75t_L g1415 ( 
.A1(n_1356),
.A2(n_1249),
.B(n_1235),
.C(n_1308),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1346),
.B(n_1223),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1330),
.Y(n_1417)
);

NAND4xp25_ASAP7_75t_L g1418 ( 
.A(n_1409),
.B(n_1351),
.C(n_1317),
.D(n_1372),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1409),
.B(n_1378),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1406),
.A2(n_1334),
.B1(n_1382),
.B2(n_1332),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1395),
.B(n_1332),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1406),
.A2(n_1382),
.B(n_1366),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1386),
.A2(n_1366),
.B(n_1377),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1383),
.B(n_1325),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1391),
.B(n_1334),
.C(n_1363),
.Y(n_1425)
);

AOI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1386),
.A2(n_1317),
.B1(n_1327),
.B2(n_1313),
.C(n_1336),
.Y(n_1426)
);

AOI221x1_ASAP7_75t_SL g1427 ( 
.A1(n_1401),
.A2(n_1316),
.B1(n_1362),
.B2(n_1359),
.C(n_1373),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1401),
.B(n_1392),
.Y(n_1428)
);

OAI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1391),
.A2(n_1334),
.B1(n_1358),
.B2(n_1374),
.C(n_1363),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1414),
.B(n_1319),
.C(n_1322),
.Y(n_1430)
);

OAI221xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1415),
.A2(n_1377),
.B1(n_1358),
.B2(n_1412),
.C(n_1402),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1415),
.A2(n_1347),
.B1(n_1378),
.B2(n_1354),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1407),
.A2(n_1336),
.B1(n_1370),
.B2(n_1367),
.C(n_1375),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1392),
.B(n_1338),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1414),
.B(n_1378),
.C(n_1343),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1414),
.B(n_1340),
.C(n_1365),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1416),
.B(n_1364),
.C(n_1337),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1392),
.B(n_1338),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1411),
.A2(n_1381),
.B1(n_1324),
.B2(n_1342),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1411),
.A2(n_1324),
.B1(n_1342),
.B2(n_1369),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1416),
.B(n_1337),
.C(n_1359),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1392),
.B(n_1314),
.Y(n_1442)
);

OAI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1416),
.A2(n_1374),
.B1(n_1324),
.B2(n_1342),
.C(n_1303),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1407),
.B(n_1318),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1383),
.B(n_1318),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1404),
.B(n_1374),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1410),
.B(n_1362),
.C(n_1373),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1403),
.A2(n_1278),
.B1(n_1374),
.B2(n_1347),
.Y(n_1448)
);

AOI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1402),
.A2(n_1333),
.B1(n_1368),
.B2(n_1360),
.C(n_1361),
.Y(n_1449)
);

NAND4xp25_ASAP7_75t_L g1450 ( 
.A(n_1399),
.B(n_1360),
.C(n_1361),
.D(n_1368),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1410),
.B(n_1355),
.C(n_1357),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1452)
);

AOI211xp5_ASAP7_75t_L g1453 ( 
.A1(n_1384),
.A2(n_1349),
.B(n_1360),
.C(n_1361),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1413),
.B(n_1388),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1396),
.B(n_1368),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1456)
);

NAND3xp33_ASAP7_75t_L g1457 ( 
.A(n_1417),
.B(n_1353),
.C(n_1355),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1397),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1399),
.B(n_1380),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1396),
.B(n_1380),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1417),
.B(n_1357),
.C(n_1353),
.Y(n_1462)
);

NOR3xp33_ASAP7_75t_L g1463 ( 
.A(n_1408),
.B(n_1376),
.C(n_1281),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1394),
.B(n_1331),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1461),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1421),
.B(n_1371),
.Y(n_1466)
);

BUFx2_ASAP7_75t_SL g1467 ( 
.A(n_1446),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1460),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1427),
.B(n_1397),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1454),
.B(n_1394),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1460),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1458),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1435),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1447),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1451),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1457),
.Y(n_1476)
);

NAND2x1_ASAP7_75t_L g1477 ( 
.A(n_1462),
.B(n_1385),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1464),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1464),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1446),
.B(n_1400),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1441),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1482)
);

NAND2x1p5_ASAP7_75t_L g1483 ( 
.A(n_1419),
.B(n_1385),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1428),
.B(n_1385),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1455),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1434),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1453),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1438),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1437),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1450),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1452),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1445),
.B(n_1387),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1430),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1456),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1442),
.Y(n_1495)
);

NOR2x1_ASAP7_75t_L g1496 ( 
.A(n_1425),
.B(n_1408),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1444),
.B(n_1387),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1456),
.B(n_1405),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1433),
.B(n_1398),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1436),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1418),
.B(n_1306),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1459),
.B(n_1405),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1496),
.B(n_1459),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1475),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1500),
.B(n_1426),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1490),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1472),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1490),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1481),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1469),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1475),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1489),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1476),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1476),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1473),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1492),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1500),
.B(n_1423),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1492),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1468),
.B(n_1419),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1400),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1467),
.B(n_1480),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1474),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1478),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1474),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1468),
.B(n_1399),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1501),
.A2(n_1432),
.B1(n_1422),
.B2(n_1429),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1485),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1485),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1489),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1478),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1408),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1497),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1479),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_SL g1536 ( 
.A(n_1473),
.B(n_1431),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1497),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1482),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1479),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1470),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1514),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1493),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1507),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1507),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1536),
.A2(n_1477),
.B(n_1473),
.Y(n_1545)
);

INVx3_ASAP7_75t_SL g1546 ( 
.A(n_1533),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1523),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1517),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1506),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1508),
.Y(n_1550)
);

NOR2x1_ASAP7_75t_L g1551 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1531),
.B(n_1504),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1471),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1526),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1512),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1519),
.B(n_1499),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1513),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1513),
.B(n_1471),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1509),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1515),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1512),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1521),
.B(n_1484),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1516),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1509),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1516),
.B(n_1466),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1510),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1521),
.B(n_1484),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1525),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1510),
.Y(n_1571)
);

AOI32xp33_ASAP7_75t_L g1572 ( 
.A1(n_1522),
.A2(n_1494),
.A3(n_1491),
.B1(n_1502),
.B2(n_1498),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1573)
);

NAND2x1_ASAP7_75t_L g1574 ( 
.A(n_1503),
.B(n_1533),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1518),
.B(n_1495),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1529),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1525),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1528),
.B(n_1491),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1503),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1522),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1559),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1548),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1503),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1545),
.A2(n_1483),
.B1(n_1420),
.B2(n_1477),
.C(n_1533),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.B(n_1534),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1559),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1550),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1541),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1566),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1582),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1554),
.B(n_1530),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1235),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1578),
.B(n_1483),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1567),
.B(n_1249),
.Y(n_1600)
);

AOI222xp33_ASAP7_75t_L g1601 ( 
.A1(n_1578),
.A2(n_1420),
.B1(n_1412),
.B2(n_1449),
.C1(n_1439),
.C2(n_1448),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1582),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1556),
.B(n_1543),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1568),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1555),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1542),
.B(n_1261),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1568),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1552),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1544),
.B(n_1530),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1547),
.B(n_1534),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1563),
.B(n_1537),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1557),
.A2(n_1537),
.B(n_1520),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1555),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

INVx5_ASAP7_75t_L g1615 ( 
.A(n_1563),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1558),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1560),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1562),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1562),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1590),
.A2(n_1561),
.B(n_1565),
.C(n_1571),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1587),
.A2(n_1553),
.B(n_1572),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1583),
.Y(n_1622)
);

AOI32xp33_ASAP7_75t_L g1623 ( 
.A1(n_1590),
.A2(n_1494),
.A3(n_1580),
.B1(n_1576),
.B2(n_1564),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1601),
.A2(n_1463),
.B(n_1569),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1601),
.A2(n_1384),
.B1(n_1390),
.B2(n_1533),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1585),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1584),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1591),
.B(n_1538),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_1575),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1587),
.A2(n_1581),
.B(n_1579),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1592),
.A2(n_1585),
.B(n_1598),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1611),
.B(n_1586),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1615),
.Y(n_1634)
);

OAI32xp33_ASAP7_75t_L g1635 ( 
.A1(n_1586),
.A2(n_1573),
.A3(n_1577),
.B1(n_1570),
.B2(n_1538),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1588),
.A2(n_1440),
.B1(n_1443),
.B2(n_1408),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1594),
.A2(n_1577),
.B1(n_1570),
.B2(n_1488),
.C(n_1486),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1589),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1595),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1615),
.B(n_1614),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1589),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1603),
.A2(n_1261),
.B(n_1201),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1594),
.B(n_1602),
.C(n_1608),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1593),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1593),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1642),
.B(n_1615),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1639),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1639),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_L g1650 ( 
.A(n_1626),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1624),
.A2(n_1600),
.B(n_1597),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1634),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1640),
.B(n_1614),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1622),
.B(n_1595),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1625),
.A2(n_1616),
.B1(n_1599),
.B2(n_1603),
.C(n_1604),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1629),
.B(n_1588),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1634),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1643),
.B(n_1606),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1631),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1632),
.B(n_1610),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1599),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1641),
.B(n_1644),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1645),
.B(n_1620),
.Y(n_1665)
);

AND4x1_ASAP7_75t_L g1666 ( 
.A(n_1654),
.B(n_1660),
.C(n_1653),
.D(n_1655),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1649),
.B(n_1628),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1665),
.A2(n_1640),
.B(n_1621),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1665),
.A2(n_1625),
.B(n_1635),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1662),
.A2(n_1630),
.B(n_1636),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1656),
.A2(n_1623),
.B(n_1637),
.C(n_1604),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1648),
.B(n_1610),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1651),
.B(n_1607),
.C(n_1617),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1658),
.A2(n_1607),
.B1(n_1617),
.B2(n_1609),
.C(n_1596),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1663),
.A2(n_1615),
.B1(n_1609),
.B2(n_1612),
.C(n_1596),
.Y(n_1676)
);

NAND4xp75_ASAP7_75t_L g1677 ( 
.A(n_1668),
.B(n_1646),
.C(n_1647),
.D(n_1652),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1667),
.B(n_1659),
.Y(n_1678)
);

AND5x1_ASAP7_75t_L g1679 ( 
.A(n_1669),
.B(n_1650),
.C(n_1615),
.D(n_1663),
.E(n_1664),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1672),
.Y(n_1680)
);

AOI211x1_ASAP7_75t_L g1681 ( 
.A1(n_1666),
.A2(n_1670),
.B(n_1675),
.C(n_1664),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1671),
.B(n_1673),
.C(n_1674),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1676),
.B(n_1657),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_L g1684 ( 
.A(n_1666),
.B(n_1661),
.C(n_1615),
.Y(n_1684)
);

NAND4xp75_ASAP7_75t_L g1685 ( 
.A(n_1668),
.B(n_1619),
.C(n_1618),
.D(n_1613),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1682),
.A2(n_1612),
.B1(n_1618),
.B2(n_1613),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1681),
.A2(n_1619),
.B1(n_1618),
.B2(n_1613),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1683),
.A2(n_1619),
.B(n_1605),
.C(n_1612),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_L g1689 ( 
.A(n_1684),
.B(n_1605),
.C(n_1306),
.D(n_1308),
.Y(n_1689)
);

OAI211xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1678),
.A2(n_1605),
.B(n_1612),
.C(n_1488),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1687),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1686),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1688),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1689),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1690),
.A2(n_1677),
.B1(n_1685),
.B2(n_1680),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1688),
.A2(n_1679),
.B1(n_1201),
.B2(n_1219),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1695),
.A2(n_1696),
.B(n_1693),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1691),
.A2(n_1219),
.B(n_1209),
.C(n_1302),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1692),
.B(n_1262),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1694),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1691),
.Y(n_1701)
);

NOR2xp67_ASAP7_75t_L g1702 ( 
.A(n_1701),
.B(n_1262),
.Y(n_1702)
);

AOI31xp33_ASAP7_75t_L g1703 ( 
.A1(n_1697),
.A2(n_1209),
.A3(n_1302),
.B(n_1237),
.Y(n_1703)
);

NOR2x1p5_ASAP7_75t_L g1704 ( 
.A(n_1698),
.B(n_1209),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1700),
.B1(n_1699),
.B2(n_1539),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1705),
.B(n_1702),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1706),
.B(n_1703),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1706),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1302),
.B1(n_1532),
.B2(n_1539),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1707),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1710),
.B(n_1532),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1709),
.A2(n_1535),
.B(n_1486),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1711),
.B(n_1262),
.C(n_1215),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1713),
.B(n_1712),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1714),
.A2(n_1535),
.B1(n_1259),
.B2(n_1215),
.Y(n_1715)
);

AOI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1527),
.B(n_1389),
.C(n_1393),
.Y(n_1716)
);


endmodule