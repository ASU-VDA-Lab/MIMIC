module real_aes_7794_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_602;
wire n_552;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_90), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g735 ( .A(n_0), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_1), .A2(n_143), .B(n_147), .C(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g196 ( .A(n_2), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_3), .A2(n_138), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_4), .B(n_160), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g164 ( .A1(n_5), .A2(n_138), .B(n_165), .Y(n_164) );
AND2x6_ASAP7_75t_L g143 ( .A(n_6), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_7), .A2(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_8), .B(n_40), .Y(n_108) );
INVx1_ASAP7_75t_L g533 ( .A(n_9), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_10), .B(n_169), .Y(n_512) );
INVx1_ASAP7_75t_L g171 ( .A(n_11), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_12), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g136 ( .A(n_13), .Y(n_136) );
INVx1_ASAP7_75t_L g252 ( .A(n_14), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_15), .A2(n_155), .B(n_253), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_16), .B(n_160), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_17), .B(n_152), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_18), .B(n_138), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_19), .B(n_561), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_20), .A2(n_179), .B(n_238), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_21), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_22), .B(n_169), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_23), .A2(n_250), .B(n_251), .C(n_253), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_24), .B(n_169), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_25), .Y(n_457) );
INVx1_ASAP7_75t_L g483 ( .A(n_26), .Y(n_483) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_28), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_29), .B(n_169), .Y(n_198) );
INVx1_ASAP7_75t_L g558 ( .A(n_30), .Y(n_558) );
INVx1_ASAP7_75t_L g185 ( .A(n_31), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_32), .A2(n_92), .B1(n_752), .B2(n_753), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_32), .Y(n_753) );
INVx2_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_34), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_35), .A2(n_156), .B(n_238), .C(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g559 ( .A(n_36), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_37), .A2(n_143), .B(n_147), .C(n_210), .Y(n_209) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_38), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_39), .A2(n_147), .B(n_482), .C(n_487), .Y(n_481) );
INVx1_ASAP7_75t_L g183 ( .A(n_41), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_42), .A2(n_49), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_42), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_43), .A2(n_63), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_43), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_44), .A2(n_728), .B1(n_729), .B2(n_732), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_44), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_45), .A2(n_168), .B(n_214), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_46), .B(n_169), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_47), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_48), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_49), .Y(n_748) );
INVx1_ASAP7_75t_L g498 ( .A(n_50), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_51), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_52), .B(n_138), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_53), .A2(n_147), .B1(n_179), .B2(n_181), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_54), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_55), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_56), .A2(n_156), .B(n_168), .C(n_170), .Y(n_167) );
CKINVDCx14_ASAP7_75t_R g530 ( .A(n_57), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_58), .Y(n_228) );
INVx1_ASAP7_75t_L g166 ( .A(n_59), .Y(n_166) );
INVx1_ASAP7_75t_L g144 ( .A(n_60), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_61), .Y(n_739) );
INVx1_ASAP7_75t_L g135 ( .A(n_62), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_63), .Y(n_730) );
INVx1_ASAP7_75t_SL g476 ( .A(n_64), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_65), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_66), .B(n_160), .Y(n_502) );
INVx1_ASAP7_75t_L g460 ( .A(n_67), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_68), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_SL g151 ( .A1(n_69), .A2(n_152), .B(n_153), .C(n_156), .Y(n_151) );
INVxp67_ASAP7_75t_L g154 ( .A(n_70), .Y(n_154) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_72), .A2(n_138), .B(n_529), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_73), .A2(n_726), .B1(n_727), .B2(n_733), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_73), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_74), .A2(n_105), .B1(n_114), .B2(n_764), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_75), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_76), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_77), .A2(n_138), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g221 ( .A(n_78), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_79), .A2(n_246), .B(n_554), .Y(n_553) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_80), .Y(n_480) );
INVx1_ASAP7_75t_L g518 ( .A(n_81), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_82), .A2(n_143), .B(n_147), .C(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_83), .A2(n_138), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g521 ( .A(n_84), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_85), .B(n_197), .Y(n_211) );
INVx2_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g511 ( .A(n_87), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_88), .B(n_152), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_89), .A2(n_143), .B(n_147), .C(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
OR2x2_ASAP7_75t_L g759 ( .A(n_90), .B(n_738), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_91), .A2(n_147), .B(n_459), .C(n_463), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_92), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_92), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_93), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_94), .A2(n_143), .B(n_147), .C(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_95), .Y(n_242) );
INVx1_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_97), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_98), .B(n_197), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_99), .B(n_131), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_100), .B(n_131), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_101), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_102), .A2(n_138), .B(n_145), .Y(n_137) );
INVx2_ASAP7_75t_L g501 ( .A(n_103), .Y(n_501) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx6p67_ASAP7_75t_R g764 ( .A(n_107), .Y(n_764) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g734 ( .A(n_108), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO221x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_740), .B1(n_745), .B2(n_755), .C(n_760), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_734), .B1(n_736), .B2(n_739), .Y(n_115) );
XOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_725), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B1(n_447), .B2(n_448), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g447 ( .A(n_120), .Y(n_447) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_120), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND4x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_365), .C(n_412), .D(n_432), .Y(n_123) );
NOR3xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_295), .C(n_320), .Y(n_124) );
OAI211xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_203), .B(n_255), .C(n_285), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_174), .Y(n_127) );
INVx3_ASAP7_75t_SL g337 ( .A(n_128), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_128), .B(n_268), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_128), .B(n_190), .Y(n_418) );
AND2x2_ASAP7_75t_L g441 ( .A(n_128), .B(n_307), .Y(n_441) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_162), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g259 ( .A(n_130), .B(n_163), .Y(n_259) );
INVx3_ASAP7_75t_L g272 ( .A(n_130), .Y(n_272) );
AND2x2_ASAP7_75t_L g277 ( .A(n_130), .B(n_162), .Y(n_277) );
OR2x2_ASAP7_75t_L g328 ( .A(n_130), .B(n_269), .Y(n_328) );
BUFx2_ASAP7_75t_L g348 ( .A(n_130), .Y(n_348) );
AND2x2_ASAP7_75t_L g358 ( .A(n_130), .B(n_269), .Y(n_358) );
AND2x2_ASAP7_75t_L g364 ( .A(n_130), .B(n_175), .Y(n_364) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_137), .B(n_159), .Y(n_130) );
INVx4_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_131), .Y(n_470) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_133), .B(n_134), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx2_ASAP7_75t_L g246 ( .A(n_138), .Y(n_246) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_139), .B(n_143), .Y(n_187) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g486 ( .A(n_140), .Y(n_486) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
INVx1_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVx1_ASAP7_75t_L g149 ( .A(n_142), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
INVx4_ASAP7_75t_SL g158 ( .A(n_143), .Y(n_158) );
BUFx3_ASAP7_75t_L g487 ( .A(n_143), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_150), .B(n_151), .C(n_158), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_146), .A2(n_158), .B(n_166), .C(n_167), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_146), .A2(n_158), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_146), .A2(n_158), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_146), .A2(n_158), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_146), .A2(n_158), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_146), .A2(n_158), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g554 ( .A1(n_146), .A2(n_158), .B(n_555), .C(n_556), .Y(n_554) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx3_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_155), .B(n_171), .Y(n_170) );
INVx5_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_155), .B(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_157), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_178), .B1(n_186), .B2(n_187), .Y(n_177) );
INVx1_ASAP7_75t_L g463 ( .A(n_158), .Y(n_463) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_160), .A2(n_164), .B(n_172), .Y(n_163) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g217 ( .A(n_161), .B(n_218), .Y(n_217) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_161), .A2(n_456), .B(n_464), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_161), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_161), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_163), .B(n_269), .Y(n_283) );
INVx2_ASAP7_75t_L g293 ( .A(n_163), .Y(n_293) );
AND2x2_ASAP7_75t_L g306 ( .A(n_163), .B(n_272), .Y(n_306) );
OR2x2_ASAP7_75t_L g317 ( .A(n_163), .B(n_269), .Y(n_317) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_163), .B(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g375 ( .A(n_163), .Y(n_375) );
AND2x2_ASAP7_75t_L g421 ( .A(n_163), .B(n_175), .Y(n_421) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g238 ( .A(n_169), .Y(n_238) );
INVx1_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
INVx2_ASAP7_75t_L g232 ( .A(n_173), .Y(n_232) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_173), .A2(n_245), .B(n_254), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_173), .A2(n_187), .B(n_480), .C(n_481), .Y(n_479) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_173), .A2(n_528), .B(n_534), .Y(n_527) );
INVx3_ASAP7_75t_SL g294 ( .A(n_174), .Y(n_294) );
OR2x2_ASAP7_75t_L g347 ( .A(n_174), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
INVx3_ASAP7_75t_L g269 ( .A(n_175), .Y(n_269) );
AND2x2_ASAP7_75t_L g336 ( .A(n_175), .B(n_191), .Y(n_336) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_175), .Y(n_404) );
AOI33xp33_ASAP7_75t_L g408 ( .A1(n_175), .A2(n_337), .A3(n_344), .B1(n_353), .B2(n_409), .B3(n_410), .Y(n_408) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_188), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_176), .B(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_176), .A2(n_192), .B(n_200), .Y(n_191) );
INVx2_ASAP7_75t_L g216 ( .A(n_176), .Y(n_216) );
INVx2_ASAP7_75t_L g199 ( .A(n_179), .Y(n_199) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_181) );
INVx2_ASAP7_75t_L g184 ( .A(n_182), .Y(n_184) );
INVx4_ASAP7_75t_L g250 ( .A(n_182), .Y(n_250) );
INVx2_ASAP7_75t_L g461 ( .A(n_184), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_187), .A2(n_193), .B(n_194), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_187), .A2(n_221), .B(n_222), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_187), .A2(n_457), .B(n_458), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_187), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g257 ( .A(n_190), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_190), .B(n_272), .Y(n_271) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_190), .B(n_332), .C(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g357 ( .A(n_190), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_190), .B(n_364), .Y(n_367) );
AND2x2_ASAP7_75t_L g420 ( .A(n_190), .B(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g276 ( .A(n_191), .Y(n_276) );
OR2x2_ASAP7_75t_L g370 ( .A(n_191), .B(n_269), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_197), .A2(n_483), .B(n_484), .C(n_485), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_197), .A2(n_250), .B1(n_558), .B2(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_202), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_202), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_202), .A2(n_507), .B(n_513), .Y(n_506) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_229), .Y(n_203) );
AOI32xp33_ASAP7_75t_L g321 ( .A1(n_204), .A2(n_322), .A3(n_324), .B1(n_326), .B2(n_329), .Y(n_321) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_204), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g424 ( .A(n_204), .Y(n_424) );
INVx4_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g356 ( .A(n_205), .B(n_340), .Y(n_356) );
AND2x2_ASAP7_75t_L g376 ( .A(n_205), .B(n_302), .Y(n_376) );
AND2x2_ASAP7_75t_L g444 ( .A(n_205), .B(n_362), .Y(n_444) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_219), .Y(n_205) );
INVx3_ASAP7_75t_L g265 ( .A(n_206), .Y(n_265) );
AND2x2_ASAP7_75t_L g279 ( .A(n_206), .B(n_263), .Y(n_279) );
OR2x2_ASAP7_75t_L g284 ( .A(n_206), .B(n_262), .Y(n_284) );
INVx1_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
AND2x2_ASAP7_75t_L g299 ( .A(n_206), .B(n_273), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_206), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_206), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g354 ( .A(n_206), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_206), .B(n_439), .Y(n_438) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AOI21xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_209), .B(n_216), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_213), .A2(n_224), .B(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_213), .A2(n_460), .B(n_461), .C(n_462), .Y(n_459) );
O2A1O1Ixp5_ASAP7_75t_L g510 ( .A1(n_213), .A2(n_461), .B(n_511), .C(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
INVx1_ASAP7_75t_L g226 ( .A(n_216), .Y(n_226) );
INVx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
AND2x2_ASAP7_75t_L g309 ( .A(n_219), .B(n_230), .Y(n_309) );
AND2x2_ASAP7_75t_L g319 ( .A(n_219), .B(n_244), .Y(n_319) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_226), .B(n_227), .Y(n_219) );
INVx1_ASAP7_75t_L g552 ( .A(n_226), .Y(n_552) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_226), .A2(n_569), .B(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g439 ( .A(n_229), .Y(n_439) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_243), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_230), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g280 ( .A(n_230), .Y(n_280) );
AND2x2_ASAP7_75t_L g324 ( .A(n_230), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g340 ( .A(n_230), .B(n_303), .Y(n_340) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
AND2x2_ASAP7_75t_L g302 ( .A(n_231), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g353 ( .A(n_231), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_231), .B(n_263), .Y(n_385) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_241), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_232), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g561 ( .A(n_232), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_239), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_238), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g264 ( .A(n_243), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g325 ( .A(n_243), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_243), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g362 ( .A(n_243), .Y(n_362) );
INVx1_ASAP7_75t_L g395 ( .A(n_243), .Y(n_395) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g273 ( .A(n_244), .B(n_263), .Y(n_273) );
INVx1_ASAP7_75t_L g303 ( .A(n_244), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_250), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_250), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_250), .B(n_521), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_260), .B1(n_266), .B2(n_273), .C(n_274), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_257), .B(n_277), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_257), .B(n_340), .Y(n_417) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_259), .B(n_307), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_259), .B(n_268), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_259), .B(n_282), .Y(n_411) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
AND2x2_ASAP7_75t_L g308 ( .A(n_264), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g386 ( .A(n_264), .Y(n_386) );
AND2x2_ASAP7_75t_L g318 ( .A(n_265), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_265), .B(n_288), .Y(n_334) );
AND2x2_ASAP7_75t_L g398 ( .A(n_265), .B(n_324), .Y(n_398) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g307 ( .A(n_269), .B(n_276), .Y(n_307) );
AND2x2_ASAP7_75t_L g403 ( .A(n_270), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_272), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_273), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_273), .B(n_280), .Y(n_368) );
AND2x2_ASAP7_75t_L g388 ( .A(n_273), .B(n_288), .Y(n_388) );
AND2x2_ASAP7_75t_L g409 ( .A(n_273), .B(n_353), .Y(n_409) );
OAI32xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .A3(n_280), .B1(n_281), .B2(n_284), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_SL g282 ( .A(n_276), .Y(n_282) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_276), .B(n_306), .Y(n_323) );
OR2x2_ASAP7_75t_L g327 ( .A(n_276), .B(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_276), .B(n_375), .Y(n_428) );
INVx1_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_278), .A2(n_369), .B1(n_415), .B2(n_418), .C(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g286 ( .A(n_279), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g329 ( .A(n_279), .B(n_302), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_279), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g407 ( .A(n_279), .B(n_340), .Y(n_407) );
INVxp67_ASAP7_75t_L g343 ( .A(n_280), .Y(n_343) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g413 ( .A(n_282), .B(n_400), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_282), .B(n_363), .Y(n_436) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_284), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g429 ( .A(n_284), .B(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_289), .B(n_292), .Y(n_285) );
AND2x2_ASAP7_75t_L g298 ( .A(n_287), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g382 ( .A(n_291), .B(n_302), .Y(n_382) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g400 ( .A(n_293), .B(n_358), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_293), .B(n_357), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_294), .B(n_306), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_300), .C(n_310), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_296), .A2(n_331), .B1(n_335), .B2(n_338), .C(n_341), .Y(n_330) );
AOI31xp33_ASAP7_75t_L g425 ( .A1(n_296), .A2(n_426), .A3(n_427), .B(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B1(n_306), .B2(n_308), .Y(n_300) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g426 ( .A(n_306), .Y(n_426) );
INVx1_ASAP7_75t_L g389 ( .A(n_307), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g432 ( .A1(n_309), .A2(n_433), .B(n_435), .C(n_437), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_314), .B2(n_318), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_315), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI221xp5_ASAP7_75t_SL g405 ( .A1(n_317), .A2(n_351), .B1(n_370), .B2(n_406), .C(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
INVx1_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g320 ( .A(n_321), .B(n_330), .C(n_345), .Y(n_320) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_322), .A2(n_372), .B(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_324), .B(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g431 ( .A(n_325), .Y(n_431) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_352), .Y(n_369) );
INVx1_ASAP7_75t_L g344 ( .A(n_333), .Y(n_344) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g342 ( .A(n_336), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_336), .B(n_374), .Y(n_373) );
NOR4xp25_ASAP7_75t_L g341 ( .A(n_337), .B(n_342), .C(n_343), .D(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI222xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_350), .B1(n_356), .B2(n_357), .C1(n_359), .C2(n_363), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g443 ( .A(n_347), .Y(n_443) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_359), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI21xp5_ASAP7_75t_SL g419 ( .A1(n_364), .A2(n_420), .B(n_422), .Y(n_419) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_377), .C(n_390), .D(n_405), .Y(n_365) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B1(n_369), .B2(n_370), .C(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g446 ( .A(n_367), .Y(n_446) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_374), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
OAI222xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .B1(n_383), .B2(n_384), .C1(n_387), .C2(n_389), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI211xp5_ASAP7_75t_L g412 ( .A1(n_382), .A2(n_413), .B(n_414), .C(n_425), .Y(n_412) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OAI222xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_396), .B1(n_397), .B2(n_399), .C1(n_401), .C2(n_402), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_407), .A2(n_410), .B1(n_443), .B2(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_440), .B(n_442), .C(n_445), .Y(n_437) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
XNOR2xp5_ASAP7_75t_L g746 ( .A(n_448), .B(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_449), .B(n_680), .Y(n_448) );
NOR4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_617), .C(n_651), .D(n_667), .Y(n_449) );
NAND4xp25_ASAP7_75t_SL g450 ( .A(n_451), .B(n_547), .C(n_581), .D(n_597), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_490), .B1(n_523), .B2(n_535), .C1(n_540), .C2(n_546), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI31xp33_ASAP7_75t_L g713 ( .A1(n_453), .A2(n_714), .A3(n_715), .B(n_717), .Y(n_713) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_466), .Y(n_453) );
AND2x2_ASAP7_75t_L g688 ( .A(n_454), .B(n_468), .Y(n_688) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_SL g539 ( .A(n_455), .Y(n_539) );
AND2x2_ASAP7_75t_L g546 ( .A(n_455), .B(n_478), .Y(n_546) );
AND2x2_ASAP7_75t_L g602 ( .A(n_455), .B(n_469), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_466), .B(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_467), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_467), .B(n_550), .Y(n_592) );
AND2x2_ASAP7_75t_L g685 ( .A(n_467), .B(n_625), .Y(n_685) );
OAI321xp33_ASAP7_75t_L g719 ( .A1(n_467), .A2(n_539), .A3(n_692), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g723 ( .A(n_467), .B(n_526), .C(n_632), .D(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g587 ( .A(n_468), .B(n_537), .Y(n_587) );
AND2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_539), .Y(n_606) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g538 ( .A(n_469), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g562 ( .A(n_469), .B(n_478), .Y(n_562) );
AND2x2_ASAP7_75t_L g648 ( .A(n_469), .B(n_537), .Y(n_648) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_477), .Y(n_469) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_470), .A2(n_496), .B(n_502), .Y(n_495) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_470), .A2(n_516), .B(n_522), .Y(n_515) );
INVx3_ASAP7_75t_SL g537 ( .A(n_478), .Y(n_537) );
AND2x2_ASAP7_75t_L g580 ( .A(n_478), .B(n_567), .Y(n_580) );
OR2x2_ASAP7_75t_L g613 ( .A(n_478), .B(n_539), .Y(n_613) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_478), .Y(n_620) );
AND2x2_ASAP7_75t_L g649 ( .A(n_478), .B(n_538), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_478), .B(n_622), .Y(n_664) );
AND2x2_ASAP7_75t_L g696 ( .A(n_478), .B(n_688), .Y(n_696) );
AND2x2_ASAP7_75t_L g705 ( .A(n_478), .B(n_551), .Y(n_705) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_486), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
INVx1_ASAP7_75t_SL g673 ( .A(n_492), .Y(n_673) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g542 ( .A(n_493), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g525 ( .A(n_494), .B(n_505), .Y(n_525) );
AND2x2_ASAP7_75t_L g609 ( .A(n_494), .B(n_527), .Y(n_609) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g579 ( .A(n_495), .B(n_515), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_495), .B(n_527), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_495), .B(n_527), .Y(n_616) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_495), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_503), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_503), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g589 ( .A(n_504), .B(n_590), .Y(n_589) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_504), .A2(n_579), .A3(n_585), .B1(n_616), .B2(n_666), .C1(n_676), .C2(n_678), .Y(n_675) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_515), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_505), .B(n_526), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_505), .B(n_527), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_505), .B(n_543), .Y(n_596) );
AND2x2_ASAP7_75t_L g650 ( .A(n_505), .B(n_616), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_505), .Y(n_654) );
AND2x2_ASAP7_75t_L g666 ( .A(n_505), .B(n_515), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_505), .B(n_542), .Y(n_698) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g563 ( .A(n_506), .B(n_515), .Y(n_563) );
BUFx3_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
AND3x2_ASAP7_75t_L g659 ( .A(n_506), .B(n_639), .C(n_660), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_515), .B(n_525), .C(n_526), .Y(n_524) );
INVx1_ASAP7_75t_SL g543 ( .A(n_515), .Y(n_543) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_515), .Y(n_644) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g638 ( .A(n_525), .B(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g645 ( .A(n_525), .Y(n_645) );
AND2x2_ASAP7_75t_L g683 ( .A(n_526), .B(n_661), .Y(n_683) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g564 ( .A(n_527), .Y(n_564) );
AND2x2_ASAP7_75t_L g639 ( .A(n_527), .B(n_543), .Y(n_639) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
OR2x2_ASAP7_75t_L g583 ( .A(n_537), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g702 ( .A(n_537), .B(n_602), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_537), .B(n_539), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_538), .B(n_551), .Y(n_657) );
AND2x2_ASAP7_75t_L g704 ( .A(n_538), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g567 ( .A(n_539), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g584 ( .A(n_539), .B(n_551), .Y(n_584) );
INVx1_ASAP7_75t_L g594 ( .A(n_539), .Y(n_594) );
AND2x2_ASAP7_75t_L g625 ( .A(n_539), .B(n_551), .Y(n_625) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_541), .A2(n_668), .B1(n_672), .B2(n_674), .C(n_675), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_544), .Y(n_541) );
AND2x2_ASAP7_75t_L g571 ( .A(n_542), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_545), .B(n_578), .Y(n_721) );
AOI322xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_563), .A3(n_564), .B1(n_565), .B2(n_571), .C1(n_573), .C2(n_580), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_562), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_550), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_550), .B(n_612), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_550), .A2(n_562), .B(n_636), .C(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_550), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_550), .B(n_606), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_550), .B(n_688), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_550), .B(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_551), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_551), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g677 ( .A(n_551), .B(n_564), .Y(n_677) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_560), .Y(n_551) );
INVx1_ASAP7_75t_L g569 ( .A(n_553), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_560), .Y(n_570) );
INVx1_ASAP7_75t_L g652 ( .A(n_562), .Y(n_652) );
OAI31xp33_ASAP7_75t_L g662 ( .A1(n_562), .A2(n_587), .A3(n_663), .B(n_665), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_562), .B(n_568), .Y(n_714) );
INVx1_ASAP7_75t_SL g575 ( .A(n_563), .Y(n_575) );
AND2x2_ASAP7_75t_L g608 ( .A(n_563), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g689 ( .A(n_563), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g574 ( .A(n_564), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g599 ( .A(n_564), .Y(n_599) );
AND2x2_ASAP7_75t_L g626 ( .A(n_564), .B(n_579), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_564), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g718 ( .A(n_564), .B(n_666), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_566), .B(n_636), .Y(n_709) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g605 ( .A(n_568), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g623 ( .A(n_568), .Y(n_623) );
NAND2xp33_ASAP7_75t_SL g573 ( .A(n_574), .B(n_576), .Y(n_573) );
OAI211xp5_ASAP7_75t_SL g617 ( .A1(n_575), .A2(n_618), .B(n_624), .C(n_640), .Y(n_617) );
OR2x2_ASAP7_75t_L g692 ( .A(n_575), .B(n_673), .Y(n_692) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
CKINVDCx16_ASAP7_75t_R g629 ( .A(n_577), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_577), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g598 ( .A(n_579), .B(n_599), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_588), .C(n_591), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g632 ( .A(n_584), .Y(n_632) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_587), .B(n_625), .Y(n_630) );
INVx1_ASAP7_75t_L g636 ( .A(n_587), .Y(n_636) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g595 ( .A(n_590), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g628 ( .A(n_590), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g690 ( .A(n_590), .Y(n_690) );
AOI21xp33_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B(n_595), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_593), .A2(n_604), .B(n_607), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_603), .C(n_610), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_598), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_601), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g614 ( .A(n_602), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_604), .A2(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_609), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g634 ( .A(n_609), .Y(n_634) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_614), .B(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g665 ( .A(n_616), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_622), .B(n_648), .Y(n_674) );
AND2x2_ASAP7_75t_L g687 ( .A(n_622), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g701 ( .A(n_622), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g711 ( .A(n_622), .B(n_649), .Y(n_711) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_627), .C(n_635), .Y(n_624) );
INVx1_ASAP7_75t_L g671 ( .A(n_625), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B1(n_631), .B2(n_633), .Y(n_627) );
OR2x2_ASAP7_75t_L g633 ( .A(n_629), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_629), .B(n_690), .Y(n_712) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g706 ( .A(n_639), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_646), .B1(n_649), .B2(n_650), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g724 ( .A(n_644), .Y(n_724) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g670 ( .A(n_648), .Y(n_670) );
OAI211xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_655), .C(n_662), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_670), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR5xp2_ASAP7_75t_L g680 ( .A(n_681), .B(n_699), .C(n_707), .D(n_713), .E(n_719), .Y(n_680) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_684), .B(n_686), .C(n_693), .Y(n_681) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_691), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_696), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B(n_706), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g722 ( .A(n_702), .Y(n_722) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g738 ( .A(n_734), .Y(n_738) );
INVx3_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g756 ( .A(n_744), .Y(n_756) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_750), .B1(n_751), .B2(n_754), .Y(n_745) );
INVx1_ASAP7_75t_L g754 ( .A(n_746), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g763 ( .A(n_759), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule