module real_jpeg_23236_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_8;
wire n_4;
wire n_6;
wire n_7;
wire n_9;

OAI21xp5_ASAP7_75t_SL g4 ( 
.A1(n_0),
.A2(n_5),
.B(n_8),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

OR2x2_ASAP7_75t_SL g6 ( 
.A(n_2),
.B(n_7),
.Y(n_6)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g3 ( 
.A(n_4),
.Y(n_3)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_6),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);


endmodule