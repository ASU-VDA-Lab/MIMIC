module fake_jpeg_11365_n_182 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_8),
.B(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_17),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_41),
.Y(n_66)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_45),
.Y(n_82)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_2),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_55),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_7),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_12),
.B(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_71),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_75),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_19),
.B1(n_23),
.B2(n_13),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_79),
.B(n_94),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_19),
.B1(n_23),
.B2(n_13),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_15),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_15),
.B1(n_22),
.B2(n_30),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_89),
.B1(n_76),
.B2(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_93),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_6),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_35),
.B1(n_58),
.B2(n_40),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_117),
.B1(n_77),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_48),
.B1(n_36),
.B2(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_116),
.B1(n_90),
.B2(n_98),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_107),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_102),
.B(n_101),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_93),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_67),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_81),
.B1(n_67),
.B2(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_66),
.B1(n_62),
.B2(n_74),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_66),
.C(n_62),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_114),
.C(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_116),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_113),
.B1(n_108),
.B2(n_100),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_84),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_136),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_114),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_143),
.B1(n_126),
.B2(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_141),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_148),
.C(n_135),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_145),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_155),
.B(n_157),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_136),
.B1(n_126),
.B2(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_129),
.B1(n_132),
.B2(n_122),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_131),
.C(n_123),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_130),
.C(n_121),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_140),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_164),
.C(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_147),
.B1(n_142),
.B2(n_120),
.Y(n_165)
);

XOR2x1_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_148),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_152),
.C(n_125),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_160),
.B1(n_163),
.B2(n_162),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_100),
.B1(n_109),
.B2(n_97),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_166),
.A2(n_143),
.B(n_125),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_173),
.C(n_172),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_170),
.C(n_176),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_109),
.C(n_106),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);


endmodule