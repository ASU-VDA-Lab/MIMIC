module fake_netlist_6_4855_n_2834 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2834);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2834;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_1371;
wire n_1285;
wire n_873;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_2247;
wire n_544;
wire n_1711;
wire n_1078;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_1986;
wire n_2300;
wire n_699;
wire n_564;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_572;
wire n_1909;
wire n_813;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_586;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1950;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_835;
wire n_850;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_627;
wire n_1767;
wire n_595;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_738;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_745;
wire n_1142;
wire n_1475;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_716;
wire n_2354;
wire n_884;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_811;
wire n_1207;
wire n_683;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2289;
wire n_1733;
wire n_2315;
wire n_1077;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1832;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_2049;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_828;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1818;
wire n_1108;
wire n_710;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_1637;
wire n_934;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_1548;
wire n_799;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_2533;
wire n_569;
wire n_1672;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1794;
wire n_1962;
wire n_786;
wire n_1236;
wire n_1650;
wire n_2398;
wire n_1725;
wire n_1928;
wire n_1559;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_2671;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_2062;
wire n_660;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_1476;
wire n_841;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1848;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_761;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_839;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_779;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1890;
wire n_1632;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_629;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1742;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_489),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_422),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_283),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_33),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_377),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_417),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_465),
.Y(n_530)
);

BUFx8_ASAP7_75t_SL g531 ( 
.A(n_145),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_135),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_370),
.Y(n_533)
);

BUFx8_ASAP7_75t_SL g534 ( 
.A(n_74),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_203),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_518),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_263),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_71),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_437),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_276),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_24),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_480),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_218),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_108),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_412),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_491),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_401),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_375),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_490),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_259),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_426),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_331),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_289),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_390),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_250),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_511),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_325),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_319),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_363),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_346),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_128),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_81),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_394),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_408),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_481),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_378),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_344),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_325),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_176),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_508),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_348),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_477),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_430),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_257),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_396),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_165),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_118),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_462),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_292),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_424),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_171),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_131),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_287),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_523),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_291),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_155),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_493),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_226),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_503),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_243),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_134),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_198),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_200),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_117),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_79),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_152),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_71),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_215),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_203),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_139),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_90),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_520),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_201),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_291),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_82),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_45),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_442),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_510),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_517),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_485),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_443),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_310),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_134),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_371),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_389),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_56),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_484),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_305),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_104),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_55),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_359),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_129),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_139),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_411),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_435),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_204),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_14),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_259),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_14),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_385),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_403),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_447),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_441),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_177),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_402),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_497),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_45),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_174),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_43),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_227),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_338),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_275),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_391),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_55),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_157),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_197),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_308),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_504),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_229),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_519),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_432),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_415),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_218),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_507),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_316),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_82),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_260),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_7),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_181),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_170),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_65),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_84),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_107),
.Y(n_669)
);

BUFx8_ASAP7_75t_SL g670 ( 
.A(n_93),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_420),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_329),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_232),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_143),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_388),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_487),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_227),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_248),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_150),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_399),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_486),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_404),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_353),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_335),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_253),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_23),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_468),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_56),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_305),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_226),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_474),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_414),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_317),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_285),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_386),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_309),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_400),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_289),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_418),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_406),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_171),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_236),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_248),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_293),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_74),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_73),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_100),
.Y(n_707)
);

CKINVDCx16_ASAP7_75t_R g708 ( 
.A(n_103),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_8),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_460),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_445),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_284),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_405),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_448),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_279),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_81),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_364),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_482),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_427),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_483),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_202),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_431),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_296),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_46),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_409),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_367),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_327),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_306),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_228),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_250),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_43),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_264),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_101),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_360),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_132),
.Y(n_735)
);

CKINVDCx14_ASAP7_75t_R g736 ( 
.A(n_108),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_18),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_349),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_243),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_398),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_242),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_152),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_331),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_84),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_463),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_450),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_310),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_369),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_433),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_221),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_454),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_181),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_332),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_80),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_160),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_281),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_379),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_183),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_425),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_215),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_211),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_340),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_476),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_155),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_355),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_146),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_374),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_73),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_416),
.Y(n_769)
);

CKINVDCx16_ASAP7_75t_R g770 ( 
.A(n_136),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_65),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_88),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_154),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_6),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_423),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_434),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_372),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_351),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_3),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_316),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_275),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_479),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_438),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_27),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_410),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_464),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_189),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_499),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_86),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_365),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_333),
.Y(n_791)
);

CKINVDCx16_ASAP7_75t_R g792 ( 
.A(n_488),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_492),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_494),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_478),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_214),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_104),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_354),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_24),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_53),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_357),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_393),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_102),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_358),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_228),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_366),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_236),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_211),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_428),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_513),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_469),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_220),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_306),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_119),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_38),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_35),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_83),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_459),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_516),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_88),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_41),
.Y(n_821)
);

CKINVDCx16_ASAP7_75t_R g822 ( 
.A(n_270),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_380),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_97),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_381),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_160),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_356),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_472),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_234),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_273),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_270),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_31),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_470),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_170),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_281),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_295),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_19),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_522),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_475),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_180),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_51),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_502),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_495),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_326),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_35),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_384),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_392),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_2),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_262),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_59),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_22),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_376),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_57),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_148),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_53),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_110),
.Y(n_856)
);

INVxp33_ASAP7_75t_SL g857 ( 
.A(n_509),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_42),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_240),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_473),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_268),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_237),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_440),
.Y(n_863)
);

CKINVDCx16_ASAP7_75t_R g864 ( 
.A(n_290),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_167),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_15),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_287),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_361),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_458),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_514),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_206),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_383),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_261),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_457),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_146),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_57),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_397),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_207),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_278),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_252),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_329),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_436),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_336),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_505),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_191),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_347),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_373),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_230),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_242),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_64),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_141),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_413),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_163),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_145),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_174),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_324),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_466),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_261),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_300),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_444),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_109),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_449),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_368),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_162),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_421),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_39),
.Y(n_906)
);

BUFx10_ASAP7_75t_L g907 ( 
.A(n_147),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_515),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_362),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_209),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_419),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_382),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_254),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_303),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_133),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_157),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_395),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_68),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_467),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_387),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_96),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_180),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_456),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_521),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_352),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_461),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_25),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_452),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_164),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_201),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_246),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_197),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_37),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_193),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_506),
.Y(n_935)
);

BUFx10_ASAP7_75t_L g936 ( 
.A(n_115),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_407),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_41),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_92),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_39),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_498),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_312),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_29),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_271),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_115),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_446),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_138),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_500),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_512),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_496),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_114),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_36),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_89),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_165),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_297),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_471),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_194),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_304),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_896),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_896),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_563),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_563),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_531),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_531),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_534),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_711),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_613),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_534),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_563),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_563),
.Y(n_970)
);

BUFx2_ASAP7_75t_SL g971 ( 
.A(n_524),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_670),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_737),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_737),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_737),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_739),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_670),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_739),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_739),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_739),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_551),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_755),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_755),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_755),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_643),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_585),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_755),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_774),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_696),
.Y(n_989)
);

CKINVDCx16_ASAP7_75t_R g990 ( 
.A(n_708),
.Y(n_990)
);

INVxp33_ASAP7_75t_L g991 ( 
.A(n_544),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_774),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_525),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_774),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_774),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_770),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_585),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_817),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_817),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_817),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_817),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_822),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_736),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_537),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_554),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_831),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_864),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_558),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_867),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_571),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_687),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_613),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_579),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_698),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_580),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_553),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_591),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_593),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_553),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_526),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_527),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_532),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_549),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_600),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_603),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_614),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_609),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_610),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_546),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_535),
.Y(n_1030)
);

INVxp67_ASAP7_75t_SL g1031 ( 
.A(n_614),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_539),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_1006),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_981),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_993),
.B(n_576),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1029),
.B(n_1012),
.Y(n_1036)
);

BUFx8_ASAP7_75t_L g1037 ( 
.A(n_965),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_969),
.Y(n_1038)
);

BUFx8_ASAP7_75t_L g1039 ( 
.A(n_967),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_969),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_974),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_974),
.Y(n_1042)
);

BUFx8_ASAP7_75t_L g1043 ( 
.A(n_967),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_978),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_1006),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_1011),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_983),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1007),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_1011),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_983),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_981),
.B(n_1003),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1026),
.B(n_636),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_985),
.A2(n_792),
.B1(n_857),
.B2(n_548),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_1003),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_961),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_962),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_970),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_986),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_1007),
.Y(n_1059)
);

AND2x6_ASAP7_75t_L g1060 ( 
.A(n_973),
.B(n_791),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_975),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_976),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_979),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1031),
.B(n_958),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_980),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_982),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_984),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_987),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_988),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_992),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_966),
.B(n_857),
.Y(n_1071)
);

BUFx12f_ASAP7_75t_L g1072 ( 
.A(n_968),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_994),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_995),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_998),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_999),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_1000),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_1001),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_1004),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1005),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1008),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1010),
.Y(n_1082)
);

CKINVDCx6p67_ASAP7_75t_R g1083 ( 
.A(n_972),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1013),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1015),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1023),
.B(n_636),
.Y(n_1086)
);

OA21x2_ASAP7_75t_L g1087 ( 
.A1(n_1017),
.A2(n_638),
.B(n_573),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_959),
.B(n_960),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1018),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_1023),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1046),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1088),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1088),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_1046),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1046),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1090),
.B(n_996),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_1058),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1080),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_1090),
.B(n_1020),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1034),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1080),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1082),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1036),
.B(n_549),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1052),
.B(n_990),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_1046),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_1054),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_1054),
.B(n_1021),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1090),
.B(n_1002),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1072),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1072),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1082),
.Y(n_1112)
);

INVxp33_ASAP7_75t_L g1113 ( 
.A(n_1053),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1084),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1043),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1084),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1046),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1035),
.B(n_872),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1079),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1083),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1079),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1043),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1079),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_1033),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1081),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1083),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1081),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1085),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1041),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1041),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1071),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1037),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1043),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1037),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1085),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1089),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1037),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1042),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1037),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_1033),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1039),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1039),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1039),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1043),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1045),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1045),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1059),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1059),
.Y(n_1148)
);

OAI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1113),
.A2(n_1131),
.B1(n_1103),
.B2(n_1118),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1129),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1129),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1119),
.B(n_1064),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1098),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1113),
.A2(n_989),
.B1(n_604),
.B2(n_944),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1130),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1091),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1092),
.A2(n_548),
.B1(n_565),
.B2(n_524),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1099),
.B(n_1064),
.Y(n_1158)
);

AND2x6_ASAP7_75t_L g1159 ( 
.A(n_1115),
.B(n_791),
.Y(n_1159)
);

XOR2xp5_ASAP7_75t_L g1160 ( 
.A(n_1097),
.B(n_986),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1130),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1096),
.B(n_971),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1105),
.B(n_1009),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1101),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1121),
.B(n_1087),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1138),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1138),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1102),
.B(n_1089),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1123),
.B(n_1114),
.C(n_1112),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1109),
.B(n_1048),
.Y(n_1170)
);

NAND2x1p5_ASAP7_75t_L g1171 ( 
.A(n_1115),
.B(n_1051),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_1091),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1116),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1093),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1125),
.Y(n_1175)
);

BUFx4f_ASAP7_75t_L g1176 ( 
.A(n_1127),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1133),
.B(n_1021),
.Y(n_1177)
);

BUFx4f_ASAP7_75t_L g1178 ( 
.A(n_1128),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1135),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1095),
.Y(n_1180)
);

AND2x6_ASAP7_75t_L g1181 ( 
.A(n_1133),
.B(n_791),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1136),
.A2(n_565),
.B1(n_641),
.B2(n_608),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1095),
.B(n_1024),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1091),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1091),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1095),
.A2(n_1087),
.B1(n_1060),
.B2(n_638),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1117),
.B(n_1025),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1117),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1117),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1094),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_1094),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1145),
.B(n_1022),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1104),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1094),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1106),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_SL g1196 ( 
.A(n_1122),
.B(n_608),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1146),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1147),
.B(n_1086),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1122),
.B(n_641),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1147),
.Y(n_1200)
);

NAND2xp33_ASAP7_75t_L g1201 ( 
.A(n_1148),
.B(n_1060),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1144),
.A2(n_718),
.B1(n_775),
.B2(n_697),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1148),
.Y(n_1203)
);

NAND2xp33_ASAP7_75t_L g1204 ( 
.A(n_1108),
.B(n_1060),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1141),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1097),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1142),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1124),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1143),
.B(n_1022),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1132),
.B(n_1087),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1134),
.B(n_1087),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1107),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1137),
.B(n_753),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1139),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1100),
.B(n_963),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1124),
.B(n_1030),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1140),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1140),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1100),
.A2(n_1060),
.B1(n_682),
.B2(n_749),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1120),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1110),
.B(n_1030),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1111),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1126),
.B(n_1032),
.Y(n_1223)
);

AND2x2_ASAP7_75t_SL g1224 ( 
.A(n_1096),
.B(n_964),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1131),
.B(n_1032),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1174),
.B(n_1028),
.Y(n_1226)
);

AO22x2_ASAP7_75t_L g1227 ( 
.A1(n_1154),
.A2(n_601),
.B1(n_944),
.B2(n_604),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1156),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1170),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1150),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1153),
.B(n_706),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_1212),
.B(n_1016),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1208),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1156),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1162),
.B(n_1225),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1155),
.Y(n_1236)
);

AND2x6_ASAP7_75t_L g1237 ( 
.A(n_1210),
.B(n_573),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1156),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1151),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1151),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1161),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1217),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1161),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1166),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1167),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1164),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1173),
.B(n_730),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1152),
.A2(n_749),
.B1(n_842),
.B2(n_682),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1168),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1152),
.A2(n_946),
.B1(n_956),
.B2(n_842),
.Y(n_1250)
);

NAND2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1200),
.B(n_753),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1168),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1179),
.Y(n_1253)
);

OR2x2_ASAP7_75t_SL g1254 ( 
.A(n_1197),
.B(n_1014),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1149),
.B(n_528),
.Y(n_1255)
);

BUFx8_ASAP7_75t_L g1256 ( 
.A(n_1205),
.Y(n_1256)
);

AO22x2_ASAP7_75t_L g1257 ( 
.A1(n_1154),
.A2(n_601),
.B1(n_958),
.B2(n_667),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1169),
.A2(n_946),
.B1(n_956),
.B2(n_872),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1183),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1192),
.B(n_968),
.C(n_1019),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1183),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1187),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1187),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1206),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1175),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1180),
.Y(n_1266)
);

OR2x2_ASAP7_75t_SL g1267 ( 
.A(n_1203),
.B(n_997),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1180),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1169),
.B(n_1158),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1214),
.B(n_885),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1198),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1202),
.B(n_997),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_SL g1273 ( 
.A(n_1205),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1200),
.B(n_783),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1214),
.B(n_1055),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1163),
.B(n_1027),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1188),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1189),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1216),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1218),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1157),
.B(n_1027),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1195),
.B(n_530),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_991),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1176),
.B(n_697),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1178),
.B(n_533),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1165),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1196),
.A2(n_572),
.B1(n_577),
.B2(n_559),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1165),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1186),
.B(n_1184),
.Y(n_1289)
);

INVx5_ASAP7_75t_L g1290 ( 
.A(n_1205),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1218),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1160),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1190),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1199),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1194),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1224),
.B(n_1210),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1211),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1185),
.B(n_783),
.Y(n_1298)
);

AND2x2_ASAP7_75t_SL g1299 ( 
.A(n_1196),
.B(n_564),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1172),
.Y(n_1300)
);

AO22x2_ASAP7_75t_L g1301 ( 
.A1(n_1182),
.A2(n_1211),
.B1(n_624),
.B2(n_690),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1185),
.B(n_912),
.Y(n_1302)
);

AO22x2_ASAP7_75t_L g1303 ( 
.A1(n_1182),
.A2(n_871),
.B1(n_901),
.B2(n_678),
.Y(n_1303)
);

AOI211xp5_ASAP7_75t_L g1304 ( 
.A1(n_1223),
.A2(n_991),
.B(n_914),
.C(n_650),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1207),
.B(n_1055),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1172),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1219),
.A2(n_1060),
.B1(n_540),
.B2(n_543),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1207),
.B(n_1056),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1159),
.B(n_1181),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1159),
.A2(n_1181),
.B1(n_1201),
.B2(n_1204),
.Y(n_1310)
);

AO22x2_ASAP7_75t_L g1311 ( 
.A1(n_1220),
.A2(n_628),
.B1(n_664),
.B2(n_564),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1221),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1191),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1191),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1191),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1159),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1213),
.B(n_1023),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1159),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1181),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1181),
.B(n_538),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1171),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1177),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1209),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1212),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1222),
.Y(n_1325)
);

AO21x1_ASAP7_75t_L g1326 ( 
.A1(n_1255),
.A2(n_561),
.B(n_547),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1290),
.Y(n_1327)
);

BUFx2_ASAP7_75t_SL g1328 ( 
.A(n_1290),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1290),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1286),
.A2(n_1060),
.B(n_568),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1286),
.A2(n_1060),
.B(n_569),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1289),
.A2(n_1049),
.B(n_775),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1288),
.A2(n_582),
.B(n_562),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1310),
.A2(n_798),
.B1(n_846),
.B2(n_718),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1234),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1235),
.B(n_1193),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1271),
.B(n_798),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1297),
.B(n_846),
.Y(n_1338)
);

CKINVDCx10_ASAP7_75t_R g1339 ( 
.A(n_1273),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1256),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1288),
.A2(n_617),
.B(n_606),
.Y(n_1341)
);

BUFx12f_ASAP7_75t_L g1342 ( 
.A(n_1256),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1296),
.A2(n_581),
.B1(n_584),
.B2(n_557),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_L g1344 ( 
.A(n_1325),
.B(n_589),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1229),
.B(n_972),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1277),
.A2(n_1293),
.B(n_1278),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1309),
.A2(n_1049),
.B(n_810),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1246),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1228),
.A2(n_1049),
.B(n_869),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1269),
.A2(n_1306),
.B(n_1300),
.Y(n_1350)
);

BUFx12f_ASAP7_75t_L g1351 ( 
.A(n_1280),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1234),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1269),
.A2(n_635),
.B1(n_645),
.B2(n_609),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1306),
.A2(n_1049),
.B(n_897),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1312),
.A2(n_637),
.B(n_657),
.C(n_647),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1279),
.A2(n_645),
.B1(n_646),
.B2(n_635),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1284),
.A2(n_594),
.B1(n_616),
.B2(n_592),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1282),
.A2(n_536),
.B(n_687),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1231),
.B(n_1247),
.Y(n_1359)
);

OAI321xp33_ASAP7_75t_L g1360 ( 
.A1(n_1281),
.A2(n_913),
.A3(n_611),
.B1(n_947),
.B2(n_814),
.C(n_652),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1291),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1233),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1231),
.B(n_1074),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1307),
.A2(n_717),
.B(n_687),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1299),
.B(n_550),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1237),
.A2(n_680),
.B(n_675),
.Y(n_1366)
);

BUFx4f_ASAP7_75t_L g1367 ( 
.A(n_1325),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1292),
.B(n_620),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1247),
.B(n_1056),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1237),
.A2(n_719),
.B(n_713),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1249),
.A2(n_672),
.B1(n_673),
.B2(n_646),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1323),
.B(n_550),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1237),
.A2(n_748),
.B(n_734),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1254),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1242),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1316),
.A2(n_717),
.B(n_687),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1276),
.B(n_977),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1316),
.A2(n_765),
.B(n_717),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1318),
.A2(n_765),
.B(n_717),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1265),
.B(n_1070),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1230),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1252),
.B(n_1070),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1301),
.A2(n_928),
.B1(n_762),
.B2(n_767),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1318),
.A2(n_776),
.B(n_765),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1226),
.B(n_1253),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1230),
.Y(n_1387)
);

O2A1O1Ixp5_ASAP7_75t_L g1388 ( 
.A1(n_1320),
.A2(n_769),
.B(n_793),
.C(n_759),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1272),
.B(n_977),
.Y(n_1389)
);

OAI21xp33_ASAP7_75t_L g1390 ( 
.A1(n_1283),
.A2(n_673),
.B(n_672),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1226),
.B(n_1261),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1319),
.A2(n_776),
.B(n_765),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1319),
.A2(n_782),
.B(n_776),
.Y(n_1393)
);

NOR2xp67_ASAP7_75t_L g1394 ( 
.A(n_1324),
.B(n_621),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1264),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1263),
.B(n_1237),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1285),
.B(n_1259),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1321),
.A2(n_804),
.B(n_809),
.C(n_802),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1270),
.B(n_1215),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1234),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1262),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1236),
.A2(n_818),
.B(n_811),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1321),
.B(n_1074),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1248),
.A2(n_833),
.B(n_825),
.Y(n_1404)
);

AO22x1_ASAP7_75t_L g1405 ( 
.A1(n_1270),
.A2(n_1324),
.B1(n_1294),
.B2(n_1317),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1303),
.A2(n_694),
.B1(n_704),
.B2(n_677),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1238),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1301),
.B(n_1075),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1266),
.A2(n_782),
.B(n_776),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1268),
.A2(n_919),
.B(n_782),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1244),
.B(n_1076),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1245),
.B(n_1057),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1239),
.A2(n_919),
.B(n_782),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1304),
.B(n_1215),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1275),
.A2(n_1308),
.B1(n_1305),
.B2(n_1232),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1240),
.A2(n_925),
.B(n_919),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1241),
.A2(n_925),
.B(n_919),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1275),
.B(n_552),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1341),
.A2(n_1260),
.B(n_1250),
.C(n_1258),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1350),
.A2(n_1331),
.B(n_1330),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1335),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1339),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1348),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_R g1424 ( 
.A(n_1351),
.B(n_1238),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1336),
.B(n_1303),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1334),
.B(n_1257),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1378),
.B(n_1308),
.C(n_1305),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1338),
.B(n_1257),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1337),
.B(n_1227),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1359),
.B(n_1227),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1361),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1367),
.B(n_1251),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1376),
.Y(n_1433)
);

INVx3_ASAP7_75t_SL g1434 ( 
.A(n_1340),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1397),
.A2(n_1238),
.B1(n_1267),
.B2(n_1313),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1360),
.A2(n_1365),
.B(n_1287),
.C(n_1373),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1367),
.B(n_1274),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1362),
.B(n_1215),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1382),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1407),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1387),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1389),
.B(n_1243),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1415),
.A2(n_1313),
.B1(n_1315),
.B2(n_1314),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1330),
.A2(n_1331),
.B(n_1332),
.Y(n_1445)
);

OAI22x1_ASAP7_75t_L g1446 ( 
.A1(n_1414),
.A2(n_1311),
.B1(n_1302),
.B2(n_1298),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1390),
.B(n_1311),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1407),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1407),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1327),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1346),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1347),
.A2(n_1333),
.B(n_1396),
.Y(n_1452)
);

O2A1O1Ixp5_ASAP7_75t_L g1453 ( 
.A1(n_1333),
.A2(n_1295),
.B(n_882),
.C(n_883),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1329),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1395),
.Y(n_1455)
);

OR2x6_ASAP7_75t_SL g1456 ( 
.A(n_1353),
.B(n_1356),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1368),
.A2(n_694),
.B1(n_704),
.B2(n_677),
.Y(n_1457)
);

AOI21xp33_ASAP7_75t_L g1458 ( 
.A1(n_1345),
.A2(n_942),
.B(n_800),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1406),
.A2(n_555),
.B1(n_588),
.B2(n_529),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1335),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1352),
.B(n_1038),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1372),
.B(n_773),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1411),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1383),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_SL g1466 ( 
.A(n_1360),
.B(n_572),
.C(n_559),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1328),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1399),
.B(n_773),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1402),
.A2(n_900),
.B(n_911),
.C(n_863),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1381),
.Y(n_1471)
);

AO21x1_ASAP7_75t_L g1472 ( 
.A1(n_1371),
.A2(n_920),
.B(n_917),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1405),
.A2(n_941),
.B(n_925),
.Y(n_1473)
);

AOI21x1_ASAP7_75t_SL g1474 ( 
.A1(n_1408),
.A2(n_555),
.B(n_529),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1403),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1369),
.B(n_800),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1344),
.B(n_862),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1363),
.B(n_1370),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1352),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1402),
.A2(n_941),
.B(n_937),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1375),
.Y(n_1481)
);

O2A1O1Ixp5_ASAP7_75t_L g1482 ( 
.A1(n_1326),
.A2(n_1371),
.B(n_1374),
.C(n_1388),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1394),
.B(n_1062),
.Y(n_1483)
);

OA22x2_ASAP7_75t_L g1484 ( 
.A1(n_1418),
.A2(n_743),
.B1(n_943),
.B2(n_577),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1400),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1374),
.A2(n_941),
.B(n_630),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1400),
.Y(n_1487)
);

OAI21xp33_ASAP7_75t_L g1488 ( 
.A1(n_1384),
.A2(n_942),
.B(n_862),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1366),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1357),
.B(n_552),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1354),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1364),
.A2(n_627),
.B(n_623),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1355),
.A2(n_619),
.B(n_633),
.C(n_626),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1343),
.A2(n_566),
.B1(n_567),
.B2(n_560),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1342),
.B(n_1398),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1404),
.A2(n_566),
.B1(n_567),
.B2(n_560),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1404),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1377),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1349),
.A2(n_1358),
.B(n_1379),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1380),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1409),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_SL g1502 ( 
.A(n_1385),
.B(n_943),
.C(n_743),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1392),
.B(n_1063),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1393),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1410),
.B(n_529),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1413),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1416),
.B(n_1063),
.Y(n_1507)
);

O2A1O1Ixp5_ASAP7_75t_SL g1508 ( 
.A1(n_1417),
.A2(n_648),
.B(n_659),
.C(n_644),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_SL g1509 ( 
.A1(n_1378),
.A2(n_1069),
.B(n_1067),
.C(n_1065),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1334),
.A2(n_574),
.B1(n_575),
.B2(n_570),
.Y(n_1510)
);

NOR2xp67_ASAP7_75t_SL g1511 ( 
.A(n_1342),
.B(n_951),
.Y(n_1511)
);

O2A1O1Ixp5_ASAP7_75t_L g1512 ( 
.A1(n_1341),
.A2(n_664),
.B(n_669),
.C(n_628),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1348),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1341),
.A2(n_928),
.B(n_685),
.C(n_686),
.Y(n_1514)
);

NAND2xp33_ASAP7_75t_L g1515 ( 
.A(n_1359),
.B(n_570),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1439),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1442),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1423),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1513),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1431),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1449),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1450),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1450),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1451),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1450),
.Y(n_1525)
);

INVx8_ASAP7_75t_L g1526 ( 
.A(n_1449),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1422),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1449),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1424),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1471),
.B(n_1475),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1454),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1465),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1497),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1488),
.A2(n_848),
.B1(n_891),
.B2(n_553),
.Y(n_1534)
);

INVx5_ASAP7_75t_L g1535 ( 
.A(n_1440),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1487),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1467),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1485),
.Y(n_1538)
);

CKINVDCx8_ASAP7_75t_R g1539 ( 
.A(n_1440),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1461),
.Y(n_1540)
);

INVx6_ASAP7_75t_L g1541 ( 
.A(n_1461),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1429),
.B(n_1447),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1454),
.Y(n_1543)
);

INVx3_ASAP7_75t_SL g1544 ( 
.A(n_1434),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1432),
.B(n_1065),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1425),
.B(n_1443),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1455),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1461),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1441),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1454),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1440),
.Y(n_1551)
);

BUFx2_ASAP7_75t_R g1552 ( 
.A(n_1456),
.Y(n_1552)
);

INVx6_ASAP7_75t_L g1553 ( 
.A(n_1448),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1448),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1421),
.B(n_1075),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1448),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1479),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1488),
.A2(n_891),
.B1(n_898),
.B2(n_848),
.Y(n_1558)
);

INVx8_ASAP7_75t_L g1559 ( 
.A(n_1421),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1468),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1427),
.B(n_1076),
.Y(n_1561)
);

INVx6_ASAP7_75t_L g1562 ( 
.A(n_1438),
.Y(n_1562)
);

CKINVDCx16_ASAP7_75t_R g1563 ( 
.A(n_1481),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1479),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1459),
.Y(n_1565)
);

INVxp67_ASAP7_75t_SL g1566 ( 
.A(n_1420),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1433),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1430),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1437),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1495),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1466),
.B(n_1428),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1462),
.Y(n_1572)
);

INVx4_ASAP7_75t_L g1573 ( 
.A(n_1501),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1435),
.Y(n_1574)
);

AO21x1_ASAP7_75t_L g1575 ( 
.A1(n_1445),
.A2(n_689),
.B(n_663),
.Y(n_1575)
);

BUFx12f_ASAP7_75t_L g1576 ( 
.A(n_1500),
.Y(n_1576)
);

INVx5_ASAP7_75t_SL g1577 ( 
.A(n_1498),
.Y(n_1577)
);

BUFx4_ASAP7_75t_SL g1578 ( 
.A(n_1464),
.Y(n_1578)
);

BUFx8_ASAP7_75t_SL g1579 ( 
.A(n_1426),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1511),
.Y(n_1580)
);

BUFx8_ASAP7_75t_L g1581 ( 
.A(n_1491),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1484),
.Y(n_1582)
);

INVx5_ASAP7_75t_L g1583 ( 
.A(n_1504),
.Y(n_1583)
);

BUFx2_ASAP7_75t_SL g1584 ( 
.A(n_1477),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1476),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1469),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1478),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1446),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1490),
.B(n_555),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1457),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1489),
.B(n_1061),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1483),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1444),
.Y(n_1593)
);

BUFx4_ASAP7_75t_SL g1594 ( 
.A(n_1506),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1463),
.Y(n_1595)
);

NAND2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1504),
.B(n_1038),
.Y(n_1596)
);

CKINVDCx16_ASAP7_75t_R g1597 ( 
.A(n_1510),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1590),
.A2(n_1460),
.B1(n_1458),
.B2(n_1496),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1532),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1595),
.B(n_1436),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1596),
.A2(n_1499),
.B(n_1452),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1534),
.A2(n_1558),
.B1(n_1590),
.B2(n_1589),
.C(n_954),
.Y(n_1602)
);

CKINVDCx8_ASAP7_75t_R g1603 ( 
.A(n_1584),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1524),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1537),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1592),
.A2(n_1419),
.B(n_1482),
.Y(n_1606)
);

AOI222xp33_ASAP7_75t_L g1607 ( 
.A1(n_1534),
.A2(n_907),
.B1(n_891),
.B2(n_936),
.C1(n_898),
.C2(n_848),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1516),
.Y(n_1608)
);

AOI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1558),
.A2(n_954),
.B1(n_952),
.B2(n_951),
.C(n_1493),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1518),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1566),
.A2(n_1480),
.B(n_1453),
.C(n_1486),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1521),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1519),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1536),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1560),
.B(n_1473),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1575),
.A2(n_1512),
.B(n_1508),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1591),
.A2(n_1474),
.B(n_1503),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1533),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1517),
.Y(n_1619)
);

NAND2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1573),
.B(n_1505),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1533),
.A2(n_1472),
.B(n_1470),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1564),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1574),
.B(n_1597),
.Y(n_1623)
);

OAI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1574),
.A2(n_1592),
.B1(n_1549),
.B2(n_1573),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1593),
.A2(n_1514),
.B(n_1507),
.Y(n_1625)
);

AO32x2_ASAP7_75t_L g1626 ( 
.A1(n_1588),
.A2(n_1509),
.A3(n_1502),
.B1(n_936),
.B2(n_907),
.Y(n_1626)
);

INVx6_ASAP7_75t_L g1627 ( 
.A(n_1526),
.Y(n_1627)
);

AOI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1591),
.A2(n_1492),
.B(n_1040),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1546),
.B(n_588),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1579),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1568),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1557),
.A2(n_1068),
.B(n_1040),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1574),
.A2(n_907),
.B1(n_936),
.B2(n_898),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1568),
.B(n_1494),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1569),
.B(n_1494),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1530),
.Y(n_1636)
);

BUFx10_ASAP7_75t_L g1637 ( 
.A(n_1547),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1552),
.A2(n_952),
.B1(n_542),
.B2(n_545),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1530),
.Y(n_1639)
);

CKINVDCx14_ASAP7_75t_R g1640 ( 
.A(n_1527),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1576),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1522),
.Y(n_1642)
);

AO21x2_ASAP7_75t_L g1643 ( 
.A1(n_1561),
.A2(n_1515),
.B(n_709),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1583),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1555),
.A2(n_1047),
.B(n_1044),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1587),
.A2(n_1050),
.B(n_1047),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1565),
.Y(n_1647)
);

OA21x2_ASAP7_75t_L g1648 ( 
.A1(n_1542),
.A2(n_1050),
.B(n_701),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1571),
.B(n_588),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1521),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1583),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1547),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1604),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1647),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1582),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1644),
.B(n_1583),
.Y(n_1656)
);

INVx5_ASAP7_75t_L g1657 ( 
.A(n_1644),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1613),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1614),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1647),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1651),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1618),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1631),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1618),
.B(n_1565),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1651),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1601),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1646),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1639),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1615),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1648),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1648),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1615),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1648),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1606),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1627),
.Y(n_1676)
);

BUFx8_ASAP7_75t_SL g1677 ( 
.A(n_1652),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1599),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1625),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1600),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1602),
.A2(n_1570),
.B1(n_1585),
.B2(n_1586),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1605),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1608),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1625),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1640),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1619),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1625),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1621),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1617),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1598),
.A2(n_1552),
.B1(n_1585),
.B2(n_1520),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1627),
.Y(n_1691)
);

INVx6_ASAP7_75t_L g1692 ( 
.A(n_1627),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1622),
.B(n_1583),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1621),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1621),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1612),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1626),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1616),
.A2(n_1538),
.B(n_701),
.Y(n_1698)
);

OR2x6_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1526),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1600),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1658),
.Y(n_1701)
);

OR2x4_ASAP7_75t_L g1702 ( 
.A(n_1664),
.B(n_1623),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_R g1703 ( 
.A(n_1685),
.B(n_1630),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_SL g1704 ( 
.A1(n_1690),
.A2(n_1602),
.B(n_1630),
.C(n_1623),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1658),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1658),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1660),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1659),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1670),
.B(n_1637),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1661),
.Y(n_1711)
);

NAND2xp33_ASAP7_75t_SL g1712 ( 
.A(n_1690),
.B(n_1594),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1677),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1691),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1686),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1675),
.A2(n_1598),
.B1(n_1607),
.B2(n_1609),
.Y(n_1716)
);

OR2x6_ASAP7_75t_L g1717 ( 
.A(n_1673),
.B(n_1526),
.Y(n_1717)
);

BUFx12f_ASAP7_75t_L g1718 ( 
.A(n_1676),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1659),
.Y(n_1719)
);

CKINVDCx16_ASAP7_75t_R g1720 ( 
.A(n_1680),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1655),
.B(n_1637),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1655),
.B(n_1520),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1673),
.B(n_1594),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1659),
.Y(n_1724)
);

NOR3xp33_ASAP7_75t_SL g1725 ( 
.A(n_1681),
.B(n_1620),
.C(n_1563),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1692),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_R g1727 ( 
.A(n_1692),
.B(n_1640),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1653),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1691),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1691),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1662),
.Y(n_1732)
);

OR2x2_ASAP7_75t_SL g1733 ( 
.A(n_1692),
.B(n_1664),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1653),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1692),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1661),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1665),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_R g1738 ( 
.A(n_1692),
.B(n_1603),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_R g1739 ( 
.A(n_1676),
.B(n_1544),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1673),
.A2(n_1620),
.B1(n_1609),
.B2(n_1581),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1665),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1686),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1669),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1669),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1696),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1678),
.B(n_1624),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1678),
.B(n_1634),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1661),
.B(n_1642),
.Y(n_1748)
);

AO21x2_ASAP7_75t_L g1749 ( 
.A1(n_1688),
.A2(n_1695),
.B(n_1689),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1661),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1686),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1732),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1705),
.Y(n_1753)
);

BUFx8_ASAP7_75t_L g1754 ( 
.A(n_1718),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1732),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1728),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1733),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1699),
.B(n_1657),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1734),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1720),
.B(n_1697),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1700),
.B(n_1682),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1708),
.B(n_1697),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1707),
.B(n_1662),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1727),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1727),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1723),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1737),
.Y(n_1767)
);

AO21x2_ASAP7_75t_L g1768 ( 
.A1(n_1749),
.A2(n_1689),
.B(n_1694),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1705),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1706),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1750),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1746),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1723),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1682),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1703),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1711),
.A2(n_1684),
.B(n_1679),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1741),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1731),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_L g1780 ( 
.A(n_1723),
.B(n_1673),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1729),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1750),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1743),
.Y(n_1783)
);

AO21x2_ASAP7_75t_L g1784 ( 
.A1(n_1768),
.A2(n_1749),
.B(n_1694),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1752),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1755),
.Y(n_1786)
);

AO21x2_ASAP7_75t_L g1787 ( 
.A1(n_1768),
.A2(n_1776),
.B(n_1769),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1772),
.B(n_1702),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1763),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1768),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1764),
.Y(n_1792)
);

INVxp67_ASAP7_75t_L g1793 ( 
.A(n_1761),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1757),
.A2(n_1716),
.B(n_1704),
.C(n_1633),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1753),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1753),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1760),
.B(n_1702),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1775),
.A2(n_1716),
.B(n_1704),
.C(n_1633),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1707),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1769),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1762),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1760),
.B(n_1744),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1770),
.Y(n_1803)
);

NOR2xp67_ASAP7_75t_L g1804 ( 
.A(n_1758),
.B(n_1657),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1776),
.A2(n_1687),
.B(n_1701),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1780),
.A2(n_1712),
.B(n_1740),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1770),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1756),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1762),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1764),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1758),
.B(n_1699),
.Y(n_1811)
);

A2O1A1Ixp33_ASAP7_75t_L g1812 ( 
.A1(n_1765),
.A2(n_1725),
.B(n_1649),
.C(n_1638),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1779),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1759),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1810),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1810),
.B(n_1765),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1812),
.A2(n_1725),
.B1(n_1773),
.B2(n_1766),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1789),
.B(n_1774),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1793),
.B(n_1788),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1791),
.B(n_1781),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1808),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1792),
.B(n_1758),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1808),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1792),
.B(n_1766),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1794),
.A2(n_712),
.B1(n_723),
.B2(n_715),
.C(n_705),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1810),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1787),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1787),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1791),
.B(n_1783),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1787),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1804),
.B(n_1766),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1811),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_L g1833 ( 
.A(n_1798),
.B(n_1581),
.C(n_724),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1805),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1813),
.B(n_1713),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1789),
.A2(n_727),
.B1(n_735),
.B2(n_729),
.C(n_728),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1805),
.Y(n_1837)
);

INVxp67_ASAP7_75t_SL g1838 ( 
.A(n_1797),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1799),
.B(n_1778),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1790),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1811),
.B(n_1766),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1790),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1784),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1811),
.B(n_1766),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1808),
.Y(n_1845)
);

INVxp67_ASAP7_75t_SL g1846 ( 
.A(n_1799),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1814),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1815),
.Y(n_1848)
);

INVxp67_ASAP7_75t_SL g1849 ( 
.A(n_1826),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1847),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1824),
.B(n_1811),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1824),
.B(n_1804),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1817),
.B(n_1806),
.Y(n_1853)
);

OR2x6_ASAP7_75t_L g1854 ( 
.A(n_1815),
.B(n_1773),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1847),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1819),
.B(n_1802),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1835),
.B(n_1779),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1841),
.B(n_1801),
.Y(n_1858)
);

XOR2xp5_ASAP7_75t_L g1859 ( 
.A(n_1833),
.B(n_1714),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1841),
.B(n_1809),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1829),
.B(n_1785),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1844),
.B(n_1785),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1844),
.B(n_1786),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1821),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1816),
.B(n_1786),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1816),
.B(n_1814),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1821),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1815),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1839),
.B(n_1803),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1823),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1823),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1839),
.B(n_1803),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1816),
.B(n_1795),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1830),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1822),
.B(n_1795),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1838),
.B(n_1820),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1830),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1849),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1851),
.B(n_1832),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1868),
.B(n_1846),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1877),
.B(n_1832),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1862),
.B(n_1818),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1850),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1854),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1858),
.B(n_1822),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1856),
.B(n_1818),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1851),
.B(n_1831),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1854),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1861),
.B(n_1845),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1855),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1858),
.B(n_1831),
.Y(n_1892)
);

OAI21xp33_ASAP7_75t_L g1893 ( 
.A1(n_1853),
.A2(n_1833),
.B(n_1836),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1864),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1867),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1870),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1860),
.B(n_1831),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1862),
.B(n_1825),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1857),
.B(n_1754),
.Y(n_1899)
);

CKINVDCx16_ASAP7_75t_R g1900 ( 
.A(n_1857),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1854),
.Y(n_1901)
);

OAI21xp33_ASAP7_75t_SL g1902 ( 
.A1(n_1853),
.A2(n_1837),
.B(n_1834),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1859),
.B(n_1754),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1863),
.B(n_1796),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1860),
.B(n_1831),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1854),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1848),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1871),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1875),
.Y(n_1909)
);

BUFx2_ASAP7_75t_SL g1910 ( 
.A(n_1848),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1863),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1866),
.B(n_1703),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1866),
.B(n_1773),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1869),
.B(n_1795),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1872),
.B(n_1796),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1865),
.B(n_1773),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1865),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1873),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1873),
.B(n_1721),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1876),
.B(n_1796),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1876),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1852),
.B(n_1767),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1907),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1879),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1892),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1881),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1893),
.B(n_849),
.C(n_724),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1897),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1893),
.B(n_1852),
.Y(n_1929)
);

AOI33xp33_ASAP7_75t_L g1930 ( 
.A1(n_1911),
.A2(n_779),
.A3(n_796),
.B1(n_805),
.B2(n_803),
.B3(n_758),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1881),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1918),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1888),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1921),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1894),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1912),
.B(n_1874),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1886),
.B(n_1874),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1898),
.B(n_1878),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1895),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1896),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1900),
.B(n_1878),
.C(n_1629),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1917),
.B(n_1800),
.Y(n_1942)
);

OAI33xp33_ASAP7_75t_L g1943 ( 
.A1(n_1898),
.A2(n_1843),
.A3(n_1842),
.B1(n_1840),
.B2(n_832),
.B3(n_821),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1882),
.B(n_1807),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1883),
.B(n_1807),
.Y(n_1945)
);

NOR2x1_ASAP7_75t_L g1946 ( 
.A(n_1910),
.B(n_1830),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1908),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1889),
.A2(n_1880),
.B1(n_1887),
.B2(n_1905),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1916),
.B(n_1544),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1885),
.Y(n_1950)
);

BUFx2_ASAP7_75t_SL g1951 ( 
.A(n_1889),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1899),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1885),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1909),
.Y(n_1954)
);

NAND2x1_ASAP7_75t_L g1955 ( 
.A(n_1913),
.B(n_1834),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1903),
.B(n_1773),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1884),
.B(n_1807),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1901),
.Y(n_1958)
);

NAND2x1_ASAP7_75t_SL g1959 ( 
.A(n_1906),
.B(n_1834),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1883),
.B(n_1800),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1891),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1890),
.Y(n_1962)
);

INVx4_ASAP7_75t_L g1963 ( 
.A(n_1920),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1919),
.B(n_1754),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1904),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1922),
.B(n_1739),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1914),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1915),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1904),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1902),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1892),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1879),
.B(n_1840),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1907),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1912),
.B(n_1739),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1879),
.B(n_1842),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1879),
.B(n_1777),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1907),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1907),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1907),
.Y(n_1979)
);

INVx1_ASAP7_75t_SL g1980 ( 
.A(n_1910),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1907),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1892),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1892),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_1907),
.Y(n_1984)
);

AO21x2_ASAP7_75t_L g1985 ( 
.A1(n_1898),
.A2(n_1843),
.B(n_1828),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1907),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1952),
.B(n_1580),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1977),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1951),
.B(n_1567),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1959),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1953),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1980),
.B(n_1827),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1956),
.B(n_1730),
.Y(n_1993)
);

OAI31xp33_ASAP7_75t_L g1994 ( 
.A1(n_1970),
.A2(n_1837),
.A3(n_1827),
.B(n_1828),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1980),
.B(n_813),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1984),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1929),
.B(n_1837),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1986),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1953),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1950),
.B(n_826),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1964),
.B(n_1926),
.Y(n_2001)
);

AND2x2_ASAP7_75t_SL g2002 ( 
.A(n_1941),
.B(n_1585),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1948),
.B(n_836),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1958),
.Y(n_2004)
);

CKINVDCx16_ASAP7_75t_R g2005 ( 
.A(n_1948),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1925),
.B(n_845),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1974),
.B(n_1529),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1949),
.B(n_1771),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_L g2009 ( 
.A(n_1927),
.B(n_732),
.C(n_669),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1946),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1928),
.B(n_851),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1971),
.B(n_855),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1982),
.B(n_875),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1933),
.B(n_1771),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1923),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1983),
.B(n_1782),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1973),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1936),
.B(n_1782),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_SL g2019 ( 
.A(n_1963),
.B(n_1579),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1955),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1962),
.B(n_876),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1978),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1936),
.B(n_1748),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1963),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1979),
.B(n_1726),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1981),
.Y(n_2026)
);

AOI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_1943),
.A2(n_890),
.B1(n_899),
.B2(n_881),
.C(n_878),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1931),
.B(n_1586),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1962),
.B(n_1523),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_1938),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1937),
.B(n_1805),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1965),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1932),
.B(n_1525),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1924),
.Y(n_2034)
);

CKINVDCx16_ASAP7_75t_R g2035 ( 
.A(n_1966),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1967),
.B(n_1699),
.Y(n_2036)
);

NOR3xp33_ASAP7_75t_SL g2037 ( 
.A(n_1972),
.B(n_556),
.C(n_541),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1968),
.B(n_1735),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1934),
.Y(n_2039)
);

NAND2x1_ASAP7_75t_L g2040 ( 
.A(n_1935),
.B(n_1805),
.Y(n_2040)
);

NOR2x1p5_ASAP7_75t_L g2041 ( 
.A(n_1927),
.B(n_1586),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1965),
.B(n_1738),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_1944),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1939),
.B(n_1562),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1945),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1969),
.B(n_1738),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1930),
.B(n_906),
.Y(n_2047)
);

NAND2x1_ASAP7_75t_L g2048 ( 
.A(n_1940),
.B(n_1717),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1947),
.B(n_916),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_1972),
.B(n_927),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1985),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1975),
.Y(n_2052)
);

OR2x6_ASAP7_75t_L g2053 ( 
.A(n_1954),
.B(n_1531),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1985),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1961),
.B(n_931),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1975),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1976),
.B(n_932),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1942),
.B(n_1717),
.Y(n_2058)
);

INVxp67_ASAP7_75t_L g2059 ( 
.A(n_1957),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1960),
.B(n_1957),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1977),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1952),
.B(n_1562),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1951),
.B(n_934),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1959),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1977),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1956),
.B(n_1717),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1977),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1956),
.B(n_1745),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1980),
.B(n_1543),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1977),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1951),
.B(n_940),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1956),
.B(n_1745),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1956),
.B(n_1745),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2032),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_2005),
.B(n_2019),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1993),
.B(n_1550),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1999),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2035),
.A2(n_1745),
.B1(n_1657),
.B2(n_1736),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2051),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2016),
.B(n_945),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2051),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2007),
.B(n_955),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_2069),
.B(n_1657),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_1987),
.Y(n_2084)
);

OAI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2030),
.A2(n_957),
.B1(n_849),
.B2(n_921),
.C(n_840),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2054),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1991),
.B(n_583),
.Y(n_2087)
);

NAND2x1_ASAP7_75t_L g2088 ( 
.A(n_1990),
.B(n_1528),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2004),
.B(n_586),
.Y(n_2089)
);

INVx1_ASAP7_75t_SL g2090 ( 
.A(n_1989),
.Y(n_2090)
);

INVxp33_ASAP7_75t_L g2091 ( 
.A(n_2001),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2038),
.B(n_732),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2024),
.B(n_1996),
.Y(n_2093)
);

INVx1_ASAP7_75t_SL g2094 ( 
.A(n_2043),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1998),
.B(n_587),
.Y(n_2095)
);

INVx1_ASAP7_75t_SL g2096 ( 
.A(n_2069),
.Y(n_2096)
);

OAI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_2036),
.A2(n_1635),
.B(n_921),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2054),
.A2(n_840),
.B1(n_953),
.B2(n_629),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2042),
.A2(n_953),
.B(n_595),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2066),
.A2(n_1635),
.B1(n_1784),
.B2(n_786),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2064),
.A2(n_1657),
.B1(n_1736),
.B2(n_1711),
.Y(n_2101)
);

INVxp67_ASAP7_75t_SL g2102 ( 
.A(n_1988),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2058),
.A2(n_1784),
.B1(n_786),
.B2(n_615),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1988),
.Y(n_2104)
);

NAND4xp25_ASAP7_75t_L g2105 ( 
.A(n_2061),
.B(n_1545),
.C(n_1578),
.D(n_1696),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2065),
.Y(n_2106)
);

OAI321xp33_ASAP7_75t_L g2107 ( 
.A1(n_2067),
.A2(n_2070),
.A3(n_2026),
.B1(n_2017),
.B2(n_2022),
.C(n_2015),
.Y(n_2107)
);

NAND2x1p5_ASAP7_75t_L g2108 ( 
.A(n_2029),
.B(n_1521),
.Y(n_2108)
);

AOI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_2010),
.A2(n_597),
.B1(n_598),
.B2(n_596),
.C(n_590),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_2020),
.Y(n_2110)
);

AOI21xp33_ASAP7_75t_L g2111 ( 
.A1(n_2048),
.A2(n_602),
.B(n_599),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1992),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2046),
.B(n_1562),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_SL g2114 ( 
.A(n_2029),
.B(n_1539),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_2018),
.Y(n_2115)
);

AOI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_2052),
.A2(n_612),
.B1(n_618),
.B2(n_607),
.C(n_605),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2063),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_2014),
.Y(n_2118)
);

AOI21xp33_ASAP7_75t_L g2119 ( 
.A1(n_2003),
.A2(n_625),
.B(n_622),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2033),
.B(n_632),
.Y(n_2120)
);

AOI221xp5_ASAP7_75t_SL g2121 ( 
.A1(n_2059),
.A2(n_1612),
.B1(n_1650),
.B2(n_1569),
.C(n_1578),
.Y(n_2121)
);

NAND3xp33_ASAP7_75t_SL g2122 ( 
.A(n_2037),
.B(n_640),
.C(n_634),
.Y(n_2122)
);

AOI21xp33_ASAP7_75t_L g2123 ( 
.A1(n_2006),
.A2(n_653),
.B(n_651),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2033),
.B(n_655),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2068),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2045),
.B(n_0),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2072),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2025),
.B(n_661),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2071),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_2014),
.Y(n_2130)
);

OR2x6_ASAP7_75t_L g2131 ( 
.A(n_1995),
.B(n_1545),
.Y(n_2131)
);

NAND3x2_ASAP7_75t_L g2132 ( 
.A(n_1997),
.B(n_1572),
.C(n_1693),
.Y(n_2132)
);

O2A1O1Ixp33_ASAP7_75t_L g2133 ( 
.A1(n_2056),
.A2(n_1643),
.B(n_1611),
.C(n_1548),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2002),
.A2(n_1657),
.B1(n_1719),
.B2(n_1696),
.Y(n_2134)
);

AOI31xp33_ASAP7_75t_L g2135 ( 
.A1(n_2009),
.A2(n_665),
.A3(n_666),
.B(n_662),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2000),
.Y(n_2136)
);

NAND3x2_ASAP7_75t_L g2137 ( 
.A(n_2060),
.B(n_1693),
.C(n_1656),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_SL g2138 ( 
.A1(n_2028),
.A2(n_1569),
.B(n_1693),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_2034),
.B(n_0),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_2053),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2057),
.Y(n_2141)
);

AOI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2041),
.A2(n_741),
.B1(n_752),
.B2(n_721),
.Y(n_2142)
);

AOI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_1994),
.A2(n_2039),
.B1(n_2025),
.B2(n_2021),
.C(n_2012),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_2053),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2044),
.A2(n_674),
.B(n_668),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2073),
.A2(n_688),
.B(n_679),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2011),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2023),
.B(n_1622),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2013),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2047),
.B(n_2062),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2049),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2050),
.B(n_693),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_2055),
.B(n_1),
.Y(n_2153)
);

NAND2xp33_ASAP7_75t_SL g2154 ( 
.A(n_2008),
.B(n_2040),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2027),
.B(n_702),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2031),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2032),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2032),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2032),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2032),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2005),
.B(n_703),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2032),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1999),
.Y(n_2163)
);

AOI221x1_ASAP7_75t_L g2164 ( 
.A1(n_2054),
.A2(n_1528),
.B1(n_1548),
.B2(n_1540),
.C(n_1612),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2032),
.Y(n_2165)
);

OR2x2_ASAP7_75t_L g2166 ( 
.A(n_2005),
.B(n_1),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2032),
.Y(n_2167)
);

AOI21xp33_ASAP7_75t_L g2168 ( 
.A1(n_2030),
.A2(n_716),
.B(n_707),
.Y(n_2168)
);

INVx1_ASAP7_75t_SL g2169 ( 
.A(n_2030),
.Y(n_2169)
);

AOI31xp33_ASAP7_75t_L g2170 ( 
.A1(n_2030),
.A2(n_733),
.A3(n_742),
.B(n_731),
.Y(n_2170)
);

NAND3xp33_ASAP7_75t_L g2171 ( 
.A(n_2005),
.B(n_747),
.C(n_744),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2032),
.Y(n_2172)
);

CKINVDCx20_ASAP7_75t_R g2173 ( 
.A(n_2035),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_2019),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2032),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2005),
.B(n_2),
.Y(n_2176)
);

INVxp67_ASAP7_75t_L g2177 ( 
.A(n_2019),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2019),
.Y(n_2178)
);

AOI21xp33_ASAP7_75t_L g2179 ( 
.A1(n_2030),
.A2(n_754),
.B(n_750),
.Y(n_2179)
);

AND2x4_ASAP7_75t_SL g2180 ( 
.A(n_2069),
.B(n_1612),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2032),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2032),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2005),
.B(n_756),
.Y(n_2183)
);

AOI32xp33_ASAP7_75t_L g2184 ( 
.A1(n_2054),
.A2(n_1696),
.A3(n_764),
.B1(n_766),
.B2(n_761),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2005),
.A2(n_797),
.B1(n_816),
.B2(n_768),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2005),
.B(n_760),
.Y(n_2186)
);

OAI222xp33_ASAP7_75t_L g2187 ( 
.A1(n_2005),
.A2(n_1657),
.B1(n_1666),
.B2(n_1656),
.C1(n_1683),
.C2(n_1693),
.Y(n_2187)
);

AOI21xp33_ASAP7_75t_L g2188 ( 
.A1(n_2030),
.A2(n_772),
.B(n_771),
.Y(n_2188)
);

OAI332xp33_ASAP7_75t_L g2189 ( 
.A1(n_2005),
.A2(n_8),
.A3(n_7),
.B1(n_5),
.B2(n_9),
.B3(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_2189)
);

AND2x2_ASAP7_75t_SL g2190 ( 
.A(n_2005),
.B(n_1650),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2005),
.B(n_4),
.Y(n_2191)
);

INVx2_ASAP7_75t_SL g2192 ( 
.A(n_2020),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2032),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1999),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2005),
.A2(n_1706),
.B1(n_1724),
.B2(n_1709),
.Y(n_2195)
);

BUFx2_ASAP7_75t_L g2196 ( 
.A(n_2032),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1993),
.B(n_1715),
.Y(n_2197)
);

BUFx2_ASAP7_75t_L g2198 ( 
.A(n_2032),
.Y(n_2198)
);

AOI32xp33_ASAP7_75t_L g2199 ( 
.A1(n_2054),
.A2(n_784),
.A3(n_787),
.B1(n_781),
.B2(n_780),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2032),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2032),
.Y(n_2201)
);

OAI21xp33_ASAP7_75t_L g2202 ( 
.A1(n_2001),
.A2(n_1666),
.B(n_799),
.Y(n_2202)
);

CKINVDCx20_ASAP7_75t_R g2203 ( 
.A(n_2035),
.Y(n_2203)
);

A2O1A1Ixp33_ASAP7_75t_L g2204 ( 
.A1(n_2054),
.A2(n_807),
.B(n_808),
.C(n_789),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2005),
.B(n_812),
.Y(n_2205)
);

OAI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2030),
.A2(n_824),
.B1(n_829),
.B2(n_820),
.C(n_815),
.Y(n_2206)
);

NAND3xp33_ASAP7_75t_L g2207 ( 
.A(n_2005),
.B(n_834),
.C(n_830),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2005),
.B(n_835),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2032),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2032),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1993),
.B(n_1742),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_1993),
.B(n_1742),
.Y(n_2212)
);

NAND3xp33_ASAP7_75t_L g2213 ( 
.A(n_2005),
.B(n_841),
.C(n_837),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1993),
.B(n_1751),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2005),
.B(n_844),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2032),
.Y(n_2216)
);

NOR3xp33_ASAP7_75t_L g2217 ( 
.A(n_2005),
.B(n_853),
.C(n_850),
.Y(n_2217)
);

A2O1A1Ixp33_ASAP7_75t_L g2218 ( 
.A1(n_2054),
.A2(n_856),
.B(n_858),
.C(n_854),
.Y(n_2218)
);

OAI22xp33_ASAP7_75t_L g2219 ( 
.A1(n_2005),
.A2(n_1650),
.B1(n_1535),
.B2(n_1751),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2032),
.Y(n_2220)
);

BUFx3_ASAP7_75t_L g2221 ( 
.A(n_2069),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2005),
.B(n_859),
.Y(n_2222)
);

AOI21xp33_ASAP7_75t_L g2223 ( 
.A1(n_2030),
.A2(n_865),
.B(n_861),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_2173),
.B(n_866),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2130),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2203),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2196),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2190),
.B(n_873),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2198),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2077),
.B(n_879),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2181),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2210),
.Y(n_2232)
);

INVxp67_ASAP7_75t_SL g2233 ( 
.A(n_2075),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2163),
.B(n_880),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2091),
.B(n_888),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2086),
.Y(n_2236)
);

OAI21xp33_ASAP7_75t_L g2237 ( 
.A1(n_2174),
.A2(n_893),
.B(n_889),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2166),
.B(n_894),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2102),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2079),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2096),
.B(n_895),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2081),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2130),
.B(n_904),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2176),
.B(n_5),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2221),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2074),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2194),
.B(n_910),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2118),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2169),
.B(n_915),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2157),
.Y(n_2250)
);

NOR3xp33_ASAP7_75t_L g2251 ( 
.A(n_2177),
.B(n_922),
.C(n_918),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2158),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_SL g2253 ( 
.A(n_2094),
.B(n_1650),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2191),
.B(n_9),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2192),
.B(n_929),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2090),
.B(n_10),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2159),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2160),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2110),
.B(n_930),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2162),
.B(n_10),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2161),
.A2(n_938),
.B(n_933),
.Y(n_2261)
);

INVx1_ASAP7_75t_SL g2262 ( 
.A(n_2115),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2165),
.B(n_939),
.Y(n_2263)
);

NOR2xp67_ASAP7_75t_L g2264 ( 
.A(n_2167),
.B(n_11),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2172),
.B(n_1709),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2175),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2125),
.B(n_1724),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2185),
.B(n_1535),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2127),
.B(n_11),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2178),
.B(n_12),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2182),
.B(n_12),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2193),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2200),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_2201),
.B(n_2209),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2216),
.B(n_13),
.Y(n_2275)
);

NAND3xp33_ASAP7_75t_L g2276 ( 
.A(n_2185),
.B(n_575),
.C(n_574),
.Y(n_2276)
);

INVx1_ASAP7_75t_SL g2277 ( 
.A(n_2180),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2220),
.B(n_13),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2076),
.B(n_15),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_2217),
.B(n_1535),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2093),
.B(n_16),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2112),
.B(n_16),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2189),
.B(n_17),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2104),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2126),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2139),
.Y(n_2286)
);

NAND4xp25_ASAP7_75t_SL g2287 ( 
.A(n_2121),
.B(n_1611),
.C(n_1687),
.D(n_19),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2108),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2082),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2117),
.B(n_17),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2129),
.B(n_18),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2080),
.B(n_20),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2106),
.B(n_20),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2088),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2140),
.B(n_21),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2144),
.B(n_21),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2131),
.B(n_22),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2156),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2183),
.B(n_23),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2114),
.B(n_1535),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2092),
.B(n_25),
.Y(n_2301)
);

OAI21xp5_ASAP7_75t_SL g2302 ( 
.A1(n_2084),
.A2(n_1540),
.B(n_1656),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2153),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2087),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2137),
.A2(n_1541),
.B1(n_1553),
.B2(n_1679),
.Y(n_2305)
);

AOI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2186),
.A2(n_1643),
.B(n_757),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2128),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2150),
.B(n_26),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2131),
.B(n_26),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2113),
.B(n_27),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_2154),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2141),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2148),
.B(n_28),
.Y(n_2313)
);

XNOR2xp5_ASAP7_75t_L g2314 ( 
.A(n_2105),
.B(n_28),
.Y(n_2314)
);

INVxp67_ASAP7_75t_L g2315 ( 
.A(n_2205),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2170),
.B(n_29),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2208),
.B(n_2215),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2142),
.B(n_30),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2195),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2222),
.B(n_30),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2147),
.Y(n_2321)
);

BUFx2_ASAP7_75t_SL g2322 ( 
.A(n_2142),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2149),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2136),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2151),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_SL g2326 ( 
.A1(n_2171),
.A2(n_1656),
.B(n_1555),
.Y(n_2326)
);

NAND2x1p5_ASAP7_75t_L g2327 ( 
.A(n_2083),
.B(n_1556),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2120),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2143),
.B(n_31),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_L g2330 ( 
.A(n_2107),
.B(n_757),
.C(n_578),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2124),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2089),
.Y(n_2332)
);

INVxp67_ASAP7_75t_L g2333 ( 
.A(n_2207),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2197),
.B(n_32),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2184),
.B(n_32),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2213),
.B(n_33),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2097),
.B(n_34),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2146),
.B(n_34),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2095),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2211),
.B(n_36),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2152),
.Y(n_2341)
);

OR2x2_ASAP7_75t_L g2342 ( 
.A(n_2132),
.B(n_37),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2225),
.Y(n_2343)
);

AOI221xp5_ASAP7_75t_L g2344 ( 
.A1(n_2311),
.A2(n_2219),
.B1(n_2199),
.B2(n_2099),
.C(n_2085),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2226),
.B(n_2109),
.Y(n_2345)
);

INVxp33_ASAP7_75t_L g2346 ( 
.A(n_2224),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2248),
.B(n_2145),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2225),
.B(n_2155),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2264),
.B(n_2202),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2262),
.B(n_2212),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2227),
.B(n_2122),
.Y(n_2351)
);

OR2x6_ASAP7_75t_L g2352 ( 
.A(n_2229),
.B(n_2204),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2274),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_2239),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2231),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2294),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2232),
.B(n_2206),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2283),
.B(n_2116),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2253),
.B(n_2078),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2256),
.Y(n_2360)
);

AOI21xp33_ASAP7_75t_L g2361 ( 
.A1(n_2233),
.A2(n_2103),
.B(n_2100),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2244),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2254),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2245),
.B(n_2168),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2298),
.B(n_2279),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2278),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2329),
.A2(n_2138),
.B1(n_2098),
.B2(n_2218),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2270),
.B(n_2214),
.Y(n_2368)
);

CKINVDCx6p67_ASAP7_75t_R g2369 ( 
.A(n_2249),
.Y(n_2369)
);

NAND2x1p5_ASAP7_75t_L g2370 ( 
.A(n_2294),
.B(n_2098),
.Y(n_2370)
);

NOR2x1_ASAP7_75t_L g2371 ( 
.A(n_2298),
.B(n_2135),
.Y(n_2371)
);

INVxp67_ASAP7_75t_SL g2372 ( 
.A(n_2316),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2334),
.B(n_2179),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2260),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2288),
.B(n_2134),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_SL g2376 ( 
.A(n_2277),
.B(n_2111),
.Y(n_2376)
);

OAI31xp33_ASAP7_75t_L g2377 ( 
.A1(n_2287),
.A2(n_2187),
.A3(n_2223),
.B(n_2188),
.Y(n_2377)
);

INVx2_ASAP7_75t_SL g2378 ( 
.A(n_2297),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2269),
.B(n_2123),
.Y(n_2379)
);

NOR2x1_ASAP7_75t_L g2380 ( 
.A(n_2282),
.B(n_2101),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2293),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2340),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2313),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2295),
.B(n_2119),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2296),
.B(n_38),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2286),
.B(n_2133),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2314),
.A2(n_2164),
.B1(n_1541),
.B2(n_1553),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2281),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2309),
.B(n_40),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2310),
.B(n_40),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_SL g2391 ( 
.A(n_2285),
.B(n_1541),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2292),
.Y(n_2392)
);

INVx2_ASAP7_75t_SL g2393 ( 
.A(n_2290),
.Y(n_2393)
);

INVx2_ASAP7_75t_SL g2394 ( 
.A(n_2291),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2319),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2289),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2246),
.B(n_42),
.Y(n_2397)
);

INVx3_ASAP7_75t_L g2398 ( 
.A(n_2327),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2271),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2250),
.B(n_2252),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2257),
.B(n_44),
.Y(n_2401)
);

INVxp67_ASAP7_75t_L g2402 ( 
.A(n_2322),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2299),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2275),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2301),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2320),
.Y(n_2406)
);

OAI31xp33_ASAP7_75t_SL g2407 ( 
.A1(n_2300),
.A2(n_2266),
.A3(n_2272),
.B(n_2258),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2317),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2273),
.B(n_44),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2303),
.B(n_615),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2308),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2236),
.Y(n_2412)
);

OAI21xp33_ASAP7_75t_L g2413 ( 
.A1(n_2326),
.A2(n_1667),
.B(n_1679),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2315),
.B(n_46),
.Y(n_2414)
);

NAND2xp33_ASAP7_75t_SL g2415 ( 
.A(n_2342),
.B(n_1551),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2230),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2240),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2333),
.B(n_47),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2234),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2247),
.Y(n_2420)
);

INVxp67_ASAP7_75t_SL g2421 ( 
.A(n_2228),
.Y(n_2421)
);

NAND3xp33_ASAP7_75t_SL g2422 ( 
.A(n_2251),
.B(n_948),
.C(n_578),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2238),
.B(n_47),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2336),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2284),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2337),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2267),
.Y(n_2427)
);

NAND2x1_ASAP7_75t_SL g2428 ( 
.A(n_2312),
.B(n_48),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2307),
.B(n_48),
.Y(n_2429)
);

INVxp67_ASAP7_75t_L g2430 ( 
.A(n_2235),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2255),
.Y(n_2431)
);

INVxp67_ASAP7_75t_L g2432 ( 
.A(n_2318),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2338),
.B(n_49),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2242),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2243),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2241),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2328),
.B(n_49),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2331),
.B(n_2341),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2259),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2341),
.B(n_50),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2339),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2339),
.B(n_50),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2332),
.B(n_51),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2304),
.B(n_52),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2321),
.B(n_2323),
.Y(n_2445)
);

NAND2x1_ASAP7_75t_L g2446 ( 
.A(n_2324),
.B(n_1553),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2325),
.B(n_52),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2263),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2265),
.Y(n_2449)
);

NOR2x1p5_ASAP7_75t_L g2450 ( 
.A(n_2335),
.B(n_1551),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2276),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2237),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2330),
.B(n_615),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2268),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2280),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_2302),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2261),
.B(n_54),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_2306),
.B(n_54),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2305),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2226),
.B(n_58),
.Y(n_2460)
);

NAND3xp33_ASAP7_75t_L g2461 ( 
.A(n_2311),
.B(n_949),
.C(n_948),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2226),
.B(n_58),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2226),
.B(n_59),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2225),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2226),
.B(n_60),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2225),
.Y(n_2466)
);

NAND2xp33_ASAP7_75t_SL g2467 ( 
.A(n_2225),
.B(n_1551),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2226),
.B(n_60),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2225),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2225),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2226),
.B(n_61),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2226),
.B(n_61),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2225),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2226),
.B(n_62),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2225),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2225),
.Y(n_2476)
);

INVx2_ASAP7_75t_SL g2477 ( 
.A(n_2225),
.Y(n_2477)
);

INVx1_ASAP7_75t_SL g2478 ( 
.A(n_2226),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2226),
.B(n_62),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2225),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2226),
.B(n_63),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2226),
.B(n_63),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2225),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2226),
.B(n_64),
.Y(n_2484)
);

INVx1_ASAP7_75t_SL g2485 ( 
.A(n_2226),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2226),
.B(n_66),
.Y(n_2486)
);

INVxp67_ASAP7_75t_L g2487 ( 
.A(n_2253),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2226),
.B(n_66),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_2226),
.B(n_786),
.Y(n_2489)
);

NAND2x1p5_ASAP7_75t_L g2490 ( 
.A(n_2226),
.B(n_1554),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2226),
.B(n_67),
.Y(n_2491)
);

AOI322xp5_ASAP7_75t_L g2492 ( 
.A1(n_2395),
.A2(n_1626),
.A3(n_1687),
.B1(n_1684),
.B2(n_1679),
.C1(n_69),
.C2(n_75),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2478),
.B(n_67),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2485),
.B(n_68),
.Y(n_2494)
);

NAND3xp33_ASAP7_75t_L g2495 ( 
.A(n_2407),
.B(n_950),
.C(n_949),
.Y(n_2495)
);

NAND5xp2_ASAP7_75t_L g2496 ( 
.A(n_2376),
.B(n_72),
.C(n_69),
.D(n_70),
.E(n_75),
.Y(n_2496)
);

AOI211xp5_ASAP7_75t_SL g2497 ( 
.A1(n_2402),
.A2(n_76),
.B(n_70),
.C(n_72),
.Y(n_2497)
);

OAI221xp5_ASAP7_75t_L g2498 ( 
.A1(n_2377),
.A2(n_2477),
.B1(n_2469),
.B2(n_2470),
.C(n_2466),
.Y(n_2498)
);

OAI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2487),
.A2(n_1667),
.B1(n_1684),
.B2(n_1554),
.Y(n_2499)
);

NOR3xp33_ASAP7_75t_L g2500 ( 
.A(n_2351),
.B(n_950),
.C(n_639),
.Y(n_2500)
);

AOI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2489),
.A2(n_642),
.B(n_631),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2428),
.Y(n_2502)
);

NAND4xp25_ASAP7_75t_L g2503 ( 
.A(n_2345),
.B(n_2344),
.C(n_2358),
.D(n_2350),
.Y(n_2503)
);

OAI211xp5_ASAP7_75t_SL g2504 ( 
.A1(n_2361),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_2504)
);

OAI211xp5_ASAP7_75t_L g2505 ( 
.A1(n_2354),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_2505)
);

NAND4xp25_ASAP7_75t_L g2506 ( 
.A(n_2364),
.B(n_85),
.C(n_80),
.D(n_83),
.Y(n_2506)
);

AND4x1_ASAP7_75t_L g2507 ( 
.A(n_2468),
.B(n_87),
.C(n_85),
.D(n_86),
.Y(n_2507)
);

OAI221xp5_ASAP7_75t_SL g2508 ( 
.A1(n_2353),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.C(n_91),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2483),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_2343),
.B(n_1554),
.Y(n_2510)
);

NAND4xp25_ASAP7_75t_L g2511 ( 
.A(n_2371),
.B(n_93),
.C(n_91),
.D(n_92),
.Y(n_2511)
);

NOR3xp33_ASAP7_75t_SL g2512 ( 
.A(n_2365),
.B(n_654),
.C(n_649),
.Y(n_2512)
);

AOI221x1_ASAP7_75t_L g2513 ( 
.A1(n_2483),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.C(n_97),
.Y(n_2513)
);

AOI221xp5_ASAP7_75t_L g2514 ( 
.A1(n_2415),
.A2(n_660),
.B1(n_671),
.B2(n_658),
.C(n_656),
.Y(n_2514)
);

NAND3x1_ASAP7_75t_L g2515 ( 
.A(n_2464),
.B(n_94),
.C(n_95),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2475),
.Y(n_2516)
);

NOR3xp33_ASAP7_75t_SL g2517 ( 
.A(n_2375),
.B(n_681),
.C(n_676),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2473),
.B(n_98),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2474),
.A2(n_2378),
.B1(n_2394),
.B2(n_2393),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_L g2520 ( 
.A(n_2476),
.B(n_684),
.C(n_683),
.Y(n_2520)
);

NOR3xp33_ASAP7_75t_L g2521 ( 
.A(n_2348),
.B(n_692),
.C(n_691),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2383),
.A2(n_1667),
.B1(n_1684),
.B2(n_1577),
.Y(n_2522)
);

OAI31xp33_ASAP7_75t_L g2523 ( 
.A1(n_2480),
.A2(n_100),
.A3(n_98),
.B(n_99),
.Y(n_2523)
);

OA21x2_ASAP7_75t_L g2524 ( 
.A1(n_2356),
.A2(n_1632),
.B(n_99),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2398),
.B(n_1564),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2463),
.B(n_2471),
.Y(n_2526)
);

INVxp67_ASAP7_75t_L g2527 ( 
.A(n_2460),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2472),
.Y(n_2528)
);

NOR3xp33_ASAP7_75t_L g2529 ( 
.A(n_2349),
.B(n_699),
.C(n_695),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_L g2530 ( 
.A(n_2391),
.B(n_710),
.C(n_700),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2481),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2482),
.B(n_101),
.Y(n_2532)
);

HB1xp67_ASAP7_75t_L g2533 ( 
.A(n_2370),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2484),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2486),
.B(n_2488),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2390),
.Y(n_2536)
);

OAI21xp33_ASAP7_75t_L g2537 ( 
.A1(n_2346),
.A2(n_1667),
.B(n_1564),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2462),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2490),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2368),
.B(n_102),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_SL g2541 ( 
.A1(n_2398),
.A2(n_106),
.B1(n_103),
.B2(n_105),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2401),
.B(n_105),
.Y(n_2542)
);

OAI22xp5_ASAP7_75t_L g2543 ( 
.A1(n_2369),
.A2(n_1577),
.B1(n_1559),
.B2(n_1671),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2382),
.B(n_106),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2366),
.B(n_107),
.Y(n_2545)
);

NAND4xp25_ASAP7_75t_SL g2546 ( 
.A(n_2355),
.B(n_111),
.C(n_109),
.D(n_110),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2362),
.B(n_111),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2410),
.A2(n_720),
.B(n_714),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2465),
.Y(n_2549)
);

NAND3x1_ASAP7_75t_SL g2550 ( 
.A(n_2380),
.B(n_112),
.C(n_113),
.Y(n_2550)
);

NOR2x1_ASAP7_75t_L g2551 ( 
.A(n_2360),
.B(n_112),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2479),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2372),
.A2(n_1559),
.B1(n_1577),
.B2(n_1698),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2491),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2389),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2408),
.B(n_113),
.Y(n_2556)
);

NOR2xp33_ASAP7_75t_L g2557 ( 
.A(n_2363),
.B(n_114),
.Y(n_2557)
);

AOI221xp5_ASAP7_75t_SL g2558 ( 
.A1(n_2359),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.C(n_119),
.Y(n_2558)
);

NAND4xp25_ASAP7_75t_L g2559 ( 
.A(n_2373),
.B(n_121),
.C(n_116),
.D(n_120),
.Y(n_2559)
);

AOI211xp5_ASAP7_75t_L g2560 ( 
.A1(n_2367),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2429),
.B(n_122),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2443),
.B(n_123),
.Y(n_2562)
);

NOR3xp33_ASAP7_75t_L g2563 ( 
.A(n_2432),
.B(n_725),
.C(n_722),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_2446),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2374),
.B(n_1559),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2385),
.Y(n_2566)
);

OAI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2400),
.A2(n_738),
.B(n_726),
.Y(n_2567)
);

NAND4xp25_ASAP7_75t_L g2568 ( 
.A(n_2396),
.B(n_125),
.C(n_123),
.D(n_124),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2459),
.A2(n_2347),
.B1(n_2424),
.B2(n_2418),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_2381),
.B(n_2388),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2455),
.A2(n_1698),
.B1(n_745),
.B2(n_746),
.Y(n_2571)
);

NAND3xp33_ASAP7_75t_L g2572 ( 
.A(n_2412),
.B(n_751),
.C(n_740),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2433),
.Y(n_2573)
);

BUFx2_ASAP7_75t_L g2574 ( 
.A(n_2352),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2426),
.A2(n_1698),
.B1(n_777),
.B2(n_778),
.Y(n_2575)
);

NAND3xp33_ASAP7_75t_SL g2576 ( 
.A(n_2357),
.B(n_785),
.C(n_763),
.Y(n_2576)
);

AOI211xp5_ASAP7_75t_L g2577 ( 
.A1(n_2454),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2397),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2447),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2550),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2493),
.B(n_2533),
.Y(n_2581)
);

XOR2x1_ASAP7_75t_L g2582 ( 
.A(n_2502),
.B(n_2417),
.Y(n_2582)
);

OAI211xp5_ASAP7_75t_L g2583 ( 
.A1(n_2519),
.A2(n_2445),
.B(n_2386),
.C(n_2434),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2558),
.B(n_2387),
.Y(n_2584)
);

AOI21xp33_ASAP7_75t_L g2585 ( 
.A1(n_2498),
.A2(n_2352),
.B(n_2384),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_SL g2586 ( 
.A1(n_2569),
.A2(n_2456),
.B(n_2419),
.Y(n_2586)
);

AOI221xp5_ASAP7_75t_SL g2587 ( 
.A1(n_2503),
.A2(n_2425),
.B1(n_2417),
.B2(n_2438),
.C(n_2451),
.Y(n_2587)
);

AOI322xp5_ASAP7_75t_L g2588 ( 
.A1(n_2574),
.A2(n_2452),
.A3(n_2411),
.B1(n_2392),
.B2(n_2420),
.C1(n_2416),
.C2(n_2405),
.Y(n_2588)
);

OAI21xp33_ASAP7_75t_SL g2589 ( 
.A1(n_2535),
.A2(n_2379),
.B(n_2421),
.Y(n_2589)
);

AOI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_2570),
.A2(n_2453),
.B(n_2440),
.Y(n_2590)
);

OAI211xp5_ASAP7_75t_SL g2591 ( 
.A1(n_2527),
.A2(n_2404),
.B(n_2399),
.C(n_2403),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2497),
.B(n_2409),
.Y(n_2592)
);

NAND4xp25_ASAP7_75t_L g2593 ( 
.A(n_2526),
.B(n_2456),
.C(n_2406),
.D(n_2430),
.Y(n_2593)
);

AOI21xp33_ASAP7_75t_L g2594 ( 
.A1(n_2534),
.A2(n_2441),
.B(n_2399),
.Y(n_2594)
);

AOI222xp33_ASAP7_75t_L g2595 ( 
.A1(n_2516),
.A2(n_2509),
.B1(n_2536),
.B2(n_2552),
.C1(n_2549),
.C2(n_2538),
.Y(n_2595)
);

OAI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2551),
.A2(n_2427),
.B(n_2461),
.Y(n_2596)
);

AOI211xp5_ASAP7_75t_L g2597 ( 
.A1(n_2504),
.A2(n_2436),
.B(n_2449),
.C(n_2422),
.Y(n_2597)
);

AOI322xp5_ASAP7_75t_L g2598 ( 
.A1(n_2554),
.A2(n_2528),
.A3(n_2531),
.B1(n_2539),
.B2(n_2573),
.C1(n_2555),
.C2(n_2566),
.Y(n_2598)
);

OAI211xp5_ASAP7_75t_L g2599 ( 
.A1(n_2564),
.A2(n_2467),
.B(n_2435),
.C(n_2431),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2544),
.B(n_2556),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2515),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2541),
.Y(n_2602)
);

AOI21xp33_ASAP7_75t_L g2603 ( 
.A1(n_2578),
.A2(n_2448),
.B(n_2439),
.Y(n_2603)
);

AOI211xp5_ASAP7_75t_SL g2604 ( 
.A1(n_2505),
.A2(n_2458),
.B(n_2414),
.C(n_2442),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_L g2605 ( 
.A1(n_2579),
.A2(n_2450),
.B1(n_2413),
.B2(n_2457),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2507),
.B(n_2437),
.Y(n_2606)
);

O2A1O1Ixp33_ASAP7_75t_L g2607 ( 
.A1(n_2511),
.A2(n_2444),
.B(n_2423),
.C(n_128),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_R g2608 ( 
.A(n_2546),
.B(n_2576),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2494),
.A2(n_2518),
.B1(n_2557),
.B2(n_2540),
.Y(n_2609)
);

AOI211xp5_ASAP7_75t_SL g2610 ( 
.A1(n_2508),
.A2(n_2547),
.B(n_2545),
.C(n_2577),
.Y(n_2610)
);

AOI211xp5_ASAP7_75t_L g2611 ( 
.A1(n_2565),
.A2(n_129),
.B(n_126),
.C(n_127),
.Y(n_2611)
);

OAI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2517),
.A2(n_790),
.B(n_788),
.Y(n_2612)
);

AOI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2532),
.A2(n_795),
.B(n_794),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2524),
.Y(n_2614)
);

AOI211xp5_ASAP7_75t_L g2615 ( 
.A1(n_2496),
.A2(n_131),
.B(n_127),
.C(n_130),
.Y(n_2615)
);

AOI211xp5_ASAP7_75t_L g2616 ( 
.A1(n_2525),
.A2(n_133),
.B(n_130),
.C(n_132),
.Y(n_2616)
);

OAI21xp33_ASAP7_75t_L g2617 ( 
.A1(n_2512),
.A2(n_806),
.B(n_801),
.Y(n_2617)
);

AOI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2510),
.A2(n_827),
.B1(n_828),
.B2(n_823),
.C(n_819),
.Y(n_2618)
);

AOI211xp5_ASAP7_75t_L g2619 ( 
.A1(n_2495),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2542),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2513),
.B(n_2523),
.Y(n_2621)
);

AOI211xp5_ASAP7_75t_L g2622 ( 
.A1(n_2568),
.A2(n_2500),
.B(n_2559),
.C(n_2506),
.Y(n_2622)
);

AOI211xp5_ASAP7_75t_L g2623 ( 
.A1(n_2529),
.A2(n_140),
.B(n_137),
.C(n_138),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2560),
.B(n_140),
.Y(n_2624)
);

AOI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2537),
.A2(n_843),
.B1(n_847),
.B2(n_839),
.C(n_838),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2561),
.Y(n_2626)
);

AOI221xp5_ASAP7_75t_L g2627 ( 
.A1(n_2543),
.A2(n_868),
.B1(n_870),
.B2(n_860),
.C(n_852),
.Y(n_2627)
);

AOI211xp5_ASAP7_75t_L g2628 ( 
.A1(n_2563),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_2628)
);

NOR4xp25_ASAP7_75t_L g2629 ( 
.A(n_2572),
.B(n_147),
.C(n_142),
.D(n_144),
.Y(n_2629)
);

AOI221xp5_ASAP7_75t_L g2630 ( 
.A1(n_2521),
.A2(n_884),
.B1(n_886),
.B2(n_877),
.C(n_874),
.Y(n_2630)
);

AOI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2562),
.A2(n_1698),
.B1(n_892),
.B2(n_902),
.Y(n_2631)
);

AOI211xp5_ASAP7_75t_L g2632 ( 
.A1(n_2520),
.A2(n_149),
.B(n_144),
.C(n_148),
.Y(n_2632)
);

OAI211xp5_ASAP7_75t_SL g2633 ( 
.A1(n_2567),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_2633)
);

NAND3xp33_ASAP7_75t_SL g2634 ( 
.A(n_2514),
.B(n_903),
.C(n_887),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2522),
.A2(n_1672),
.B1(n_1674),
.B2(n_1671),
.Y(n_2635)
);

AOI211xp5_ASAP7_75t_L g2636 ( 
.A1(n_2530),
.A2(n_154),
.B(n_151),
.C(n_153),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2501),
.B(n_153),
.Y(n_2637)
);

NAND3xp33_ASAP7_75t_SL g2638 ( 
.A(n_2601),
.B(n_2548),
.C(n_2492),
.Y(n_2638)
);

OAI21xp33_ASAP7_75t_SL g2639 ( 
.A1(n_2614),
.A2(n_2580),
.B(n_2621),
.Y(n_2639)
);

XNOR2xp5_ASAP7_75t_L g2640 ( 
.A(n_2615),
.B(n_2571),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2582),
.B(n_2492),
.Y(n_2641)
);

NAND4xp25_ASAP7_75t_L g2642 ( 
.A(n_2585),
.B(n_2499),
.C(n_2575),
.D(n_2553),
.Y(n_2642)
);

OAI21xp5_ASAP7_75t_SL g2643 ( 
.A1(n_2586),
.A2(n_2583),
.B(n_2604),
.Y(n_2643)
);

AOI211xp5_ASAP7_75t_L g2644 ( 
.A1(n_2594),
.A2(n_2524),
.B(n_159),
.C(n_156),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2602),
.B(n_156),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2581),
.B(n_158),
.Y(n_2646)
);

OAI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2605),
.A2(n_908),
.B1(n_909),
.B2(n_905),
.Y(n_2647)
);

A2O1A1Ixp33_ASAP7_75t_L g2648 ( 
.A1(n_2607),
.A2(n_161),
.B(n_158),
.C(n_159),
.Y(n_2648)
);

OAI21xp5_ASAP7_75t_SL g2649 ( 
.A1(n_2610),
.A2(n_161),
.B(n_162),
.Y(n_2649)
);

AOI221xp5_ASAP7_75t_L g2650 ( 
.A1(n_2587),
.A2(n_926),
.B1(n_935),
.B2(n_924),
.C(n_923),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2600),
.B(n_163),
.Y(n_2651)
);

AO21x1_ASAP7_75t_L g2652 ( 
.A1(n_2592),
.A2(n_164),
.B(n_166),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2626),
.Y(n_2653)
);

AOI221xp5_ASAP7_75t_L g2654 ( 
.A1(n_2603),
.A2(n_2591),
.B1(n_2593),
.B2(n_2599),
.C(n_2589),
.Y(n_2654)
);

AOI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2606),
.A2(n_166),
.B(n_167),
.Y(n_2655)
);

OA211x2_ASAP7_75t_L g2656 ( 
.A1(n_2584),
.A2(n_172),
.B(n_168),
.C(n_169),
.Y(n_2656)
);

OAI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_2609),
.A2(n_1671),
.B1(n_1674),
.B2(n_1672),
.Y(n_2657)
);

NOR3xp33_ASAP7_75t_L g2658 ( 
.A(n_2590),
.B(n_168),
.C(n_169),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2626),
.Y(n_2659)
);

INVxp67_ASAP7_75t_L g2660 ( 
.A(n_2624),
.Y(n_2660)
);

AOI211xp5_ASAP7_75t_L g2661 ( 
.A1(n_2596),
.A2(n_175),
.B(n_172),
.C(n_173),
.Y(n_2661)
);

A2O1A1Ixp33_ASAP7_75t_L g2662 ( 
.A1(n_2598),
.A2(n_176),
.B(n_173),
.C(n_175),
.Y(n_2662)
);

AOI221xp5_ASAP7_75t_L g2663 ( 
.A1(n_2629),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.C(n_182),
.Y(n_2663)
);

AOI21xp5_ASAP7_75t_SL g2664 ( 
.A1(n_2617),
.A2(n_178),
.B(n_179),
.Y(n_2664)
);

AOI222xp33_ASAP7_75t_L g2665 ( 
.A1(n_2620),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.C1(n_185),
.C2(n_186),
.Y(n_2665)
);

AOI221x1_ASAP7_75t_SL g2666 ( 
.A1(n_2597),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.C(n_187),
.Y(n_2666)
);

BUFx8_ASAP7_75t_SL g2667 ( 
.A(n_2626),
.Y(n_2667)
);

AOI221xp5_ASAP7_75t_L g2668 ( 
.A1(n_2608),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2637),
.Y(n_2669)
);

AOI322xp5_ASAP7_75t_L g2670 ( 
.A1(n_2634),
.A2(n_188),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.C1(n_193),
.C2(n_194),
.Y(n_2670)
);

OAI211xp5_ASAP7_75t_L g2671 ( 
.A1(n_2595),
.A2(n_196),
.B(n_192),
.C(n_195),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2588),
.B(n_195),
.Y(n_2672)
);

OA22x2_ASAP7_75t_L g2673 ( 
.A1(n_2612),
.A2(n_199),
.B1(n_196),
.B2(n_198),
.Y(n_2673)
);

OAI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_2672),
.A2(n_2631),
.B1(n_2613),
.B2(n_2627),
.Y(n_2674)
);

AOI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2643),
.A2(n_2633),
.B1(n_2622),
.B2(n_2611),
.Y(n_2675)
);

AOI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2639),
.A2(n_2616),
.B1(n_2619),
.B2(n_2623),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2646),
.B(n_2636),
.Y(n_2677)
);

AOI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2651),
.A2(n_2618),
.B(n_2632),
.Y(n_2678)
);

NOR3xp33_ASAP7_75t_L g2679 ( 
.A(n_2654),
.B(n_2630),
.C(n_2628),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2638),
.A2(n_2625),
.B1(n_2635),
.B2(n_1674),
.Y(n_2680)
);

OAI21xp5_ASAP7_75t_SL g2681 ( 
.A1(n_2649),
.A2(n_199),
.B(n_200),
.Y(n_2681)
);

OR2x2_ASAP7_75t_L g2682 ( 
.A(n_2645),
.B(n_202),
.Y(n_2682)
);

OAI221xp5_ASAP7_75t_L g2683 ( 
.A1(n_2666),
.A2(n_2662),
.B1(n_2641),
.B2(n_2663),
.C(n_2648),
.Y(n_2683)
);

OAI32xp33_ASAP7_75t_L g2684 ( 
.A1(n_2660),
.A2(n_204),
.A3(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2653),
.B(n_205),
.Y(n_2685)
);

OAI211xp5_ASAP7_75t_L g2686 ( 
.A1(n_2671),
.A2(n_2644),
.B(n_2664),
.C(n_2642),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2661),
.A2(n_1672),
.B1(n_1628),
.B2(n_1668),
.Y(n_2687)
);

AOI22x1_ASAP7_75t_L g2688 ( 
.A1(n_2653),
.A2(n_2659),
.B1(n_2655),
.B2(n_2640),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2659),
.B(n_208),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2667),
.A2(n_1067),
.B1(n_1069),
.B2(n_1066),
.Y(n_2690)
);

AOI221xp5_ASAP7_75t_L g2691 ( 
.A1(n_2652),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.C(n_212),
.Y(n_2691)
);

AOI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2658),
.A2(n_213),
.B1(n_210),
.B2(n_212),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2669),
.B(n_2647),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2685),
.Y(n_2694)
);

AOI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2686),
.A2(n_2656),
.B1(n_2673),
.B2(n_2668),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2677),
.B(n_2676),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_L g2697 ( 
.A(n_2683),
.B(n_2650),
.Y(n_2697)
);

AOI211xp5_ASAP7_75t_L g2698 ( 
.A1(n_2681),
.A2(n_2657),
.B(n_2670),
.C(n_2665),
.Y(n_2698)
);

NOR2x1_ASAP7_75t_L g2699 ( 
.A(n_2689),
.B(n_213),
.Y(n_2699)
);

NAND4xp75_ASAP7_75t_L g2700 ( 
.A(n_2675),
.B(n_217),
.C(n_214),
.D(n_216),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2685),
.Y(n_2701)
);

NAND3xp33_ASAP7_75t_L g2702 ( 
.A(n_2691),
.B(n_2688),
.C(n_2679),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2682),
.B(n_216),
.Y(n_2703)
);

NAND4xp25_ASAP7_75t_L g2704 ( 
.A(n_2678),
.B(n_220),
.C(n_217),
.D(n_219),
.Y(n_2704)
);

NAND3x1_ASAP7_75t_L g2705 ( 
.A(n_2692),
.B(n_2680),
.C(n_2684),
.Y(n_2705)
);

INVx2_ASAP7_75t_SL g2706 ( 
.A(n_2693),
.Y(n_2706)
);

INVx5_ASAP7_75t_L g2707 ( 
.A(n_2690),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2674),
.Y(n_2708)
);

A2O1A1Ixp33_ASAP7_75t_L g2709 ( 
.A1(n_2687),
.A2(n_222),
.B(n_219),
.C(n_221),
.Y(n_2709)
);

AOI211xp5_ASAP7_75t_L g2710 ( 
.A1(n_2683),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2700),
.Y(n_2711)
);

CKINVDCx20_ASAP7_75t_R g2712 ( 
.A(n_2696),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2706),
.Y(n_2713)
);

INVx1_ASAP7_75t_SL g2714 ( 
.A(n_2701),
.Y(n_2714)
);

BUFx2_ASAP7_75t_L g2715 ( 
.A(n_2699),
.Y(n_2715)
);

NAND2x1p5_ASAP7_75t_L g2716 ( 
.A(n_2694),
.B(n_1645),
.Y(n_2716)
);

CKINVDCx20_ASAP7_75t_R g2717 ( 
.A(n_2695),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_2708),
.Y(n_2718)
);

NOR2x1_ASAP7_75t_L g2719 ( 
.A(n_2704),
.B(n_223),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2703),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2702),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2710),
.B(n_224),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2705),
.Y(n_2723)
);

CKINVDCx16_ASAP7_75t_R g2724 ( 
.A(n_2697),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2698),
.Y(n_2725)
);

AOI211xp5_ASAP7_75t_L g2726 ( 
.A1(n_2709),
.A2(n_230),
.B(n_225),
.C(n_229),
.Y(n_2726)
);

INVx1_ASAP7_75t_SL g2727 ( 
.A(n_2707),
.Y(n_2727)
);

BUFx3_ASAP7_75t_L g2728 ( 
.A(n_2707),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2706),
.Y(n_2729)
);

AO22x2_ASAP7_75t_L g2730 ( 
.A1(n_2714),
.A2(n_232),
.B1(n_225),
.B2(n_231),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2718),
.B(n_231),
.Y(n_2731)
);

INVx5_ASAP7_75t_L g2732 ( 
.A(n_2718),
.Y(n_2732)
);

OAI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2713),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2729),
.Y(n_2734)
);

OAI22xp5_ASAP7_75t_SL g2735 ( 
.A1(n_2712),
.A2(n_237),
.B1(n_233),
.B2(n_235),
.Y(n_2735)
);

OAI22xp5_ASAP7_75t_SL g2736 ( 
.A1(n_2717),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2718),
.Y(n_2737)
);

XNOR2x1_ASAP7_75t_L g2738 ( 
.A(n_2719),
.B(n_238),
.Y(n_2738)
);

NAND3xp33_ASAP7_75t_SL g2739 ( 
.A(n_2726),
.B(n_239),
.C(n_241),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2723),
.B(n_241),
.Y(n_2740)
);

XNOR2x1_ASAP7_75t_L g2741 ( 
.A(n_2721),
.B(n_244),
.Y(n_2741)
);

NOR2x1_ASAP7_75t_L g2742 ( 
.A(n_2715),
.B(n_244),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_SL g2743 ( 
.A1(n_2728),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_2743)
);

XOR2x2_ASAP7_75t_L g2744 ( 
.A(n_2722),
.B(n_245),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_2727),
.Y(n_2745)
);

AOI22x1_ASAP7_75t_L g2746 ( 
.A1(n_2724),
.A2(n_251),
.B1(n_247),
.B2(n_249),
.Y(n_2746)
);

OAI22x1_ASAP7_75t_L g2747 ( 
.A1(n_2711),
.A2(n_252),
.B1(n_249),
.B2(n_251),
.Y(n_2747)
);

XNOR2x1_ASAP7_75t_L g2748 ( 
.A(n_2725),
.B(n_2720),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_SL g2749 ( 
.A1(n_2716),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2742),
.Y(n_2750)
);

INVxp67_ASAP7_75t_SL g2751 ( 
.A(n_2747),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2740),
.Y(n_2752)
);

AO21x2_ASAP7_75t_L g2753 ( 
.A1(n_2731),
.A2(n_255),
.B(n_256),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2730),
.Y(n_2754)
);

AO22x2_ASAP7_75t_L g2755 ( 
.A1(n_2741),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2755)
);

AOI22xp33_ASAP7_75t_L g2756 ( 
.A1(n_2737),
.A2(n_1067),
.B1(n_1069),
.B2(n_1066),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2745),
.B(n_258),
.Y(n_2757)
);

AOI21xp33_ASAP7_75t_L g2758 ( 
.A1(n_2734),
.A2(n_260),
.B(n_262),
.Y(n_2758)
);

XNOR2xp5_ASAP7_75t_L g2759 ( 
.A(n_2748),
.B(n_263),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2736),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2732),
.Y(n_2761)
);

NAND2x1_ASAP7_75t_L g2762 ( 
.A(n_2749),
.B(n_264),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2746),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_SL g2764 ( 
.A1(n_2738),
.A2(n_265),
.B(n_266),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2759),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2755),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2753),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2757),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2762),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2751),
.Y(n_2770)
);

CKINVDCx20_ASAP7_75t_R g2771 ( 
.A(n_2760),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2761),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2761),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2754),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2750),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2763),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2752),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2764),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2778),
.Y(n_2779)
);

INVxp67_ASAP7_75t_SL g2780 ( 
.A(n_2778),
.Y(n_2780)
);

OAI22x1_ASAP7_75t_SL g2781 ( 
.A1(n_2770),
.A2(n_2732),
.B1(n_2744),
.B2(n_2739),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2767),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2769),
.Y(n_2783)
);

OAI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2772),
.A2(n_2758),
.B(n_2743),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_SL g2785 ( 
.A1(n_2771),
.A2(n_2735),
.B1(n_2756),
.B2(n_2733),
.Y(n_2785)
);

BUFx2_ASAP7_75t_L g2786 ( 
.A(n_2766),
.Y(n_2786)
);

OAI22xp33_ASAP7_75t_L g2787 ( 
.A1(n_2773),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_SL g2788 ( 
.A1(n_2775),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_2788)
);

OAI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2774),
.A2(n_269),
.B(n_271),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2776),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2777),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2791)
);

OAI322xp33_ASAP7_75t_L g2792 ( 
.A1(n_2765),
.A2(n_272),
.A3(n_274),
.B1(n_276),
.B2(n_277),
.C1(n_278),
.C2(n_279),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2768),
.A2(n_277),
.B1(n_280),
.B2(n_282),
.Y(n_2793)
);

OAI21xp5_ASAP7_75t_SL g2794 ( 
.A1(n_2783),
.A2(n_280),
.B(n_282),
.Y(n_2794)
);

OAI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2790),
.A2(n_2786),
.B1(n_2780),
.B2(n_2779),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2788),
.Y(n_2796)
);

OAI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2782),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2785),
.A2(n_286),
.B1(n_288),
.B2(n_290),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2781),
.A2(n_286),
.B1(n_288),
.B2(n_292),
.Y(n_2799)
);

INVx1_ASAP7_75t_SL g2800 ( 
.A(n_2791),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2789),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_SL g2802 ( 
.A1(n_2784),
.A2(n_293),
.B(n_294),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2792),
.Y(n_2803)
);

NAND2xp33_ASAP7_75t_SL g2804 ( 
.A(n_2787),
.B(n_2793),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2790),
.Y(n_2805)
);

AOI211xp5_ASAP7_75t_L g2806 ( 
.A1(n_2795),
.A2(n_294),
.B(n_295),
.C(n_296),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2805),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_2807)
);

NOR2xp67_ASAP7_75t_L g2808 ( 
.A(n_2794),
.B(n_298),
.Y(n_2808)
);

NAND5xp2_ASAP7_75t_L g2809 ( 
.A(n_2803),
.B(n_299),
.C(n_300),
.D(n_301),
.E(n_302),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2799),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_2810)
);

OAI211xp5_ASAP7_75t_SL g2811 ( 
.A1(n_2800),
.A2(n_2796),
.B(n_2801),
.C(n_2802),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2798),
.A2(n_304),
.B1(n_307),
.B2(n_308),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2797),
.Y(n_2813)
);

OAI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2804),
.A2(n_307),
.B1(n_309),
.B2(n_311),
.Y(n_2814)
);

OAI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2805),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2805),
.Y(n_2816)
);

AOI22xp33_ASAP7_75t_L g2817 ( 
.A1(n_2816),
.A2(n_1066),
.B1(n_1073),
.B2(n_1077),
.Y(n_2817)
);

OAI33xp33_ASAP7_75t_R g2818 ( 
.A1(n_2809),
.A2(n_313),
.A3(n_314),
.B1(n_315),
.B2(n_317),
.B3(n_318),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_R g2819 ( 
.A(n_2813),
.B(n_314),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2808),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_2820)
);

AOI32xp33_ASAP7_75t_L g2821 ( 
.A1(n_2811),
.A2(n_2810),
.A3(n_2812),
.B1(n_2814),
.B2(n_2806),
.Y(n_2821)
);

AOI222xp33_ASAP7_75t_L g2822 ( 
.A1(n_2807),
.A2(n_2815),
.B1(n_321),
.B2(n_322),
.C1(n_323),
.C2(n_324),
.Y(n_2822)
);

OAI222xp33_ASAP7_75t_L g2823 ( 
.A1(n_2816),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.C1(n_323),
.C2(n_326),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2816),
.A2(n_320),
.B(n_327),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2808),
.Y(n_2825)
);

OAI32xp33_ASAP7_75t_L g2826 ( 
.A1(n_2816),
.A2(n_328),
.A3(n_330),
.B1(n_334),
.B2(n_337),
.Y(n_2826)
);

AOI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2820),
.A2(n_328),
.B1(n_330),
.B2(n_1078),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_R g2828 ( 
.A1(n_2819),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2825),
.A2(n_2822),
.B1(n_2824),
.B2(n_2818),
.Y(n_2829)
);

AOI22xp5_ASAP7_75t_SL g2830 ( 
.A1(n_2821),
.A2(n_343),
.B1(n_345),
.B2(n_350),
.Y(n_2830)
);

AO21x2_ASAP7_75t_L g2831 ( 
.A1(n_2829),
.A2(n_2823),
.B(n_2817),
.Y(n_2831)
);

AOI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2827),
.A2(n_2826),
.B1(n_1078),
.B2(n_1077),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2831),
.A2(n_2830),
.B(n_2828),
.Y(n_2833)
);

AOI211xp5_ASAP7_75t_L g2834 ( 
.A1(n_2833),
.A2(n_2832),
.B(n_1078),
.C(n_1077),
.Y(n_2834)
);


endmodule