module fake_jpeg_9105_n_53 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_15),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_12),
.B(n_20),
.C(n_19),
.D(n_18),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_25),
.A3(n_13),
.B1(n_8),
.B2(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_30),
.B1(n_5),
.B2(n_7),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_4),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_23),
.B1(n_25),
.B2(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_41),
.B1(n_42),
.B2(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_4),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_33),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B(n_47),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_35),
.A3(n_42),
.B1(n_39),
.B2(n_5),
.C1(n_7),
.C2(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_43),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_46),
.B(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_45),
.Y(n_53)
);


endmodule