module real_aes_17777_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_1395, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_1395;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1172 ( .A1(n_0), .A2(n_175), .B1(n_1142), .B2(n_1146), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_1), .A2(n_181), .B1(n_782), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_1), .A2(n_53), .B1(n_563), .B2(n_916), .Y(n_915) );
OAI211xp5_ASAP7_75t_L g502 ( .A1(n_2), .A2(n_503), .B(n_505), .C(n_520), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_2), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_3), .A2(n_105), .B1(n_921), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_SL g1114 ( .A1(n_3), .A2(n_112), .B1(n_828), .B2(n_1115), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_4), .A2(n_41), .B1(n_1142), .B2(n_1146), .Y(n_1180) );
INVx1_ASAP7_75t_L g904 ( .A(n_5), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g922 ( .A1(n_5), .A2(n_55), .B1(n_566), .B2(n_715), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_6), .A2(n_58), .B1(n_547), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_6), .A2(n_43), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_7), .A2(n_195), .B1(n_782), .B2(n_892), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_7), .A2(n_223), .B1(n_563), .B2(n_742), .Y(n_1369) );
INVx1_ASAP7_75t_L g603 ( .A(n_8), .Y(n_603) );
AO22x1_ASAP7_75t_L g629 ( .A1(n_8), .A2(n_130), .B1(n_515), .B2(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g248 ( .A(n_9), .Y(n_248) );
AND2x2_ASAP7_75t_L g301 ( .A(n_9), .B(n_204), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_9), .B(n_258), .Y(n_320) );
AND2x2_ASAP7_75t_L g334 ( .A(n_9), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g613 ( .A(n_10), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_10), .A2(n_81), .B1(n_474), .B2(n_510), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_11), .A2(n_140), .B1(n_577), .B2(n_1092), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1108 ( .A1(n_11), .A2(n_14), .B1(n_898), .B2(n_1109), .C(n_1110), .Y(n_1108) );
INVx2_ASAP7_75t_L g1145 ( .A(n_12), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_12), .B(n_85), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_12), .B(n_1151), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_13), .A2(n_74), .B1(n_538), .B2(n_909), .Y(n_1363) );
AOI22xp33_ASAP7_75t_SL g1098 ( .A1(n_14), .A2(n_25), .B1(n_702), .B2(n_755), .Y(n_1098) );
INVx1_ASAP7_75t_L g1089 ( .A(n_15), .Y(n_1089) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_16), .A2(n_187), .B1(n_715), .B2(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1118 ( .A(n_16), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_17), .A2(n_23), .B1(n_1149), .B2(n_1152), .Y(n_1166) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_18), .A2(n_108), .B1(n_1149), .B2(n_1152), .Y(n_1171) );
INVx1_ASAP7_75t_L g1048 ( .A(n_19), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1066 ( .A1(n_19), .A2(n_154), .B1(n_715), .B2(n_1067), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_20), .A2(n_46), .B1(n_803), .B2(n_884), .C(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1079 ( .A(n_20), .Y(n_1079) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_21), .A2(n_522), .B(n_524), .C(n_526), .Y(n_521) );
INVx1_ASAP7_75t_L g582 ( .A(n_21), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_22), .A2(n_79), .B1(n_538), .B2(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_24), .A2(n_226), .B1(n_987), .B2(n_991), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_24), .A2(n_226), .B1(n_1026), .B2(n_1029), .Y(n_1025) );
A2O1A1Ixp33_ASAP7_75t_L g1121 ( .A1(n_25), .A2(n_802), .B(n_1122), .C(n_1128), .Y(n_1121) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_26), .B(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_26), .A2(n_141), .B1(n_368), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_27), .A2(n_77), .B1(n_1142), .B2(n_1301), .Y(n_1300) );
XNOR2xp5_ASAP7_75t_L g1343 ( .A(n_27), .B(n_1344), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_27), .A2(n_1379), .B1(n_1384), .B2(n_1389), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_28), .A2(n_141), .B1(n_507), .B2(n_630), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_28), .A2(n_217), .B1(n_368), .B2(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g886 ( .A(n_29), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_30), .A2(n_72), .B1(n_1142), .B2(n_1160), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_31), .A2(n_48), .B1(n_538), .B2(n_757), .Y(n_1104) );
OAI211xp5_ASAP7_75t_L g1106 ( .A1(n_31), .A2(n_894), .B(n_1107), .C(n_1116), .Y(n_1106) );
XOR2x2_ASAP7_75t_L g816 ( .A(n_32), .B(n_817), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_33), .A2(n_149), .B1(n_782), .B2(n_900), .Y(n_1357) );
AOI22xp33_ASAP7_75t_SL g1371 ( .A1(n_33), .A2(n_109), .B1(n_391), .B2(n_763), .Y(n_1371) );
INVx1_ASAP7_75t_L g435 ( .A(n_34), .Y(n_435) );
XNOR2x2_ASAP7_75t_L g1083 ( .A(n_35), .B(n_1084), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_36), .A2(n_54), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_36), .A2(n_231), .B1(n_370), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_37), .A2(n_117), .B1(n_752), .B2(n_753), .Y(n_751) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_37), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g1385 ( .A1(n_38), .A2(n_1386), .B1(n_1387), .B2(n_1388), .Y(n_1385) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_38), .Y(n_1386) );
INVx1_ASAP7_75t_L g358 ( .A(n_39), .Y(n_358) );
INVx1_ASAP7_75t_L g366 ( .A(n_39), .Y(n_366) );
INVx1_ASAP7_75t_L g661 ( .A(n_40), .Y(n_661) );
INVxp67_ASAP7_75t_SL g1039 ( .A(n_41), .Y(n_1039) );
AND4x1_ASAP7_75t_L g1082 ( .A(n_41), .B(n_1041), .C(n_1044), .D(n_1064), .Y(n_1082) );
AOI22xp5_ASAP7_75t_L g1177 ( .A1(n_42), .A2(n_114), .B1(n_1142), .B2(n_1160), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_43), .A2(n_123), .B1(n_547), .B2(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_44), .A2(n_202), .B1(n_1149), .B2(n_1152), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_45), .A2(n_112), .B1(n_921), .B2(n_947), .Y(n_1096) );
AOI221xp5_ASAP7_75t_L g1123 ( .A1(n_45), .A2(n_105), .B1(n_838), .B2(n_1124), .C(n_1125), .Y(n_1123) );
INVx1_ASAP7_75t_L g1081 ( .A(n_46), .Y(n_1081) );
INVx1_ASAP7_75t_L g241 ( .A(n_47), .Y(n_241) );
INVx2_ASAP7_75t_L g378 ( .A(n_49), .Y(n_378) );
INVx1_ASAP7_75t_L g649 ( .A(n_50), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_51), .A2(n_103), .B1(n_777), .B2(n_823), .C(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g873 ( .A(n_51), .Y(n_873) );
INVx1_ASAP7_75t_L g759 ( .A(n_52), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_53), .A2(n_172), .B1(n_835), .B2(n_897), .C(n_898), .Y(n_896) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_54), .A2(n_80), .B1(n_370), .B2(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g903 ( .A(n_55), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_56), .A2(n_115), .B1(n_828), .B2(n_829), .Y(n_833) );
INVx1_ASAP7_75t_L g860 ( .A(n_56), .Y(n_860) );
INVx1_ASAP7_75t_L g713 ( .A(n_57), .Y(n_713) );
INVx1_ASAP7_75t_L g795 ( .A(n_58), .Y(n_795) );
INVx1_ASAP7_75t_L g464 ( .A(n_59), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_59), .A2(n_113), .B1(n_473), .B2(n_476), .C(n_483), .Y(n_482) );
AOI21xp33_ASAP7_75t_L g889 ( .A1(n_60), .A2(n_836), .B(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_60), .A2(n_155), .B1(n_391), .B2(n_568), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_61), .A2(n_183), .B1(n_646), .B2(n_757), .Y(n_1043) );
OAI211xp5_ASAP7_75t_L g1045 ( .A1(n_61), .A2(n_894), .B(n_1046), .C(n_1049), .Y(n_1045) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_62), .A2(n_182), .B1(n_407), .B2(n_411), .C1(n_620), .C2(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g633 ( .A(n_62), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g883 ( .A1(n_63), .A2(n_884), .B(n_885), .C(n_887), .Y(n_883) );
INVx1_ASAP7_75t_L g913 ( .A(n_63), .Y(n_913) );
INVx1_ASAP7_75t_L g734 ( .A(n_64), .Y(n_734) );
OAI222xp33_ASAP7_75t_L g786 ( .A1(n_64), .A2(n_106), .B1(n_787), .B2(n_790), .C1(n_796), .C2(n_803), .Y(n_786) );
OAI22xp5_ASAP7_75t_SL g671 ( .A1(n_65), .A2(n_83), .B1(n_672), .B2(n_673), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g687 ( .A1(n_65), .A2(n_566), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g839 ( .A(n_66), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_67), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_68), .A2(n_89), .B1(n_1142), .B2(n_1146), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_69), .A2(n_107), .B1(n_1149), .B2(n_1152), .Y(n_1157) );
INVx1_ASAP7_75t_L g1348 ( .A(n_70), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_71), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_73), .A2(n_229), .B1(n_515), .B2(n_1055), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_73), .A2(n_93), .B1(n_1072), .B2(n_1073), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1353 ( .A1(n_74), .A2(n_1354), .B(n_1355), .C(n_1358), .Y(n_1353) );
INVx1_ASAP7_75t_L g317 ( .A(n_75), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_75), .A2(n_192), .B1(n_380), .B2(n_382), .C(n_385), .Y(n_379) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_76), .Y(n_243) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_76), .B(n_241), .Y(n_1143) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_78), .Y(n_595) );
OAI211xp5_ASAP7_75t_SL g893 ( .A1(n_79), .A2(n_894), .B(n_895), .C(n_902), .Y(n_893) );
AOI221xp5_ASAP7_75t_SL g517 ( .A1(n_80), .A2(n_231), .B1(n_474), .B2(n_518), .C(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g609 ( .A(n_81), .Y(n_609) );
OAI211xp5_ASAP7_75t_L g665 ( .A1(n_82), .A2(n_666), .B(n_667), .C(n_668), .Y(n_665) );
INVxp33_ASAP7_75t_SL g689 ( .A(n_82), .Y(n_689) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_83), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_84), .Y(n_726) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_85), .B(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1151 ( .A(n_85), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_86), .A2(n_206), .B1(n_420), .B2(n_423), .Y(n_419) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_86), .Y(n_429) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_87), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g1076 ( .A1(n_87), .A2(n_185), .B1(n_389), .B2(n_1077), .Y(n_1076) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_88), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_90), .A2(n_150), .B1(n_1149), .B2(n_1152), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_91), .Y(n_1042) );
INVx1_ASAP7_75t_L g843 ( .A(n_92), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_93), .A2(n_194), .B1(n_510), .B2(n_825), .C(n_1062), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_94), .Y(n_956) );
INVx1_ASAP7_75t_L g376 ( .A(n_95), .Y(n_376) );
INVx2_ASAP7_75t_L g387 ( .A(n_95), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_95), .B(n_378), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_96), .A2(n_135), .B1(n_362), .B2(n_390), .Y(n_469) );
INVx1_ASAP7_75t_L g484 ( .A(n_96), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g1351 ( .A1(n_97), .A2(n_512), .B(n_776), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_97), .A2(n_149), .B1(n_391), .B2(n_568), .Y(n_1370) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_98), .A2(n_156), .B1(n_997), .B2(n_998), .Y(n_996) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_98), .A2(n_156), .B1(n_1005), .B2(n_1008), .Y(n_1004) );
INVx1_ASAP7_75t_L g339 ( .A(n_99), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_100), .A2(n_132), .B1(n_271), .B2(n_278), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_100), .A2(n_180), .B1(n_389), .B2(n_391), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_101), .A2(n_125), .B1(n_522), .B2(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g561 ( .A(n_101), .Y(n_561) );
INVx1_ASAP7_75t_L g617 ( .A(n_102), .Y(n_617) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_102), .B(n_474), .Y(n_642) );
INVx1_ASAP7_75t_L g861 ( .A(n_103), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_104), .B(n_728), .Y(n_879) );
INVx1_ASAP7_75t_L g732 ( .A(n_106), .Y(n_732) );
INVxp67_ASAP7_75t_SL g1350 ( .A(n_109), .Y(n_1350) );
INVx1_ASAP7_75t_L g1362 ( .A(n_110), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_111), .A2(n_212), .B1(n_1149), .B2(n_1152), .Y(n_1148) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_113), .A2(n_215), .B1(n_369), .B2(n_458), .C(n_459), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g436 ( .A(n_114), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g869 ( .A(n_115), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_116), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_117), .A2(n_227), .B1(n_772), .B2(n_775), .C(n_777), .Y(n_771) );
OAI211xp5_ASAP7_75t_SL g974 ( .A1(n_118), .A2(n_969), .B(n_975), .C(n_978), .Y(n_974) );
INVx1_ASAP7_75t_L g1024 ( .A(n_118), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_119), .A2(n_120), .B1(n_1142), .B2(n_1146), .Y(n_1156) );
INVx1_ASAP7_75t_L g1360 ( .A(n_121), .Y(n_1360) );
OAI22xp33_ASAP7_75t_L g1373 ( .A1(n_121), .A2(n_161), .B1(n_566), .B2(n_1374), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_122), .Y(n_951) );
INVx1_ASAP7_75t_L g791 ( .A(n_123), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_124), .A2(n_128), .B1(n_1149), .B2(n_1152), .Y(n_1179) );
INVx1_ASAP7_75t_L g579 ( .A(n_125), .Y(n_579) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_126), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_127), .A2(n_228), .B1(n_420), .B2(n_423), .Y(n_444) );
INVxp33_ASAP7_75t_SL g494 ( .A(n_127), .Y(n_494) );
NAND5xp2_ASAP7_75t_L g500 ( .A(n_129), .B(n_501), .C(n_540), .D(n_564), .E(n_573), .Y(n_500) );
INVx1_ASAP7_75t_L g586 ( .A(n_129), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_130), .A2(n_375), .B(n_390), .Y(n_618) );
INVx1_ASAP7_75t_L g644 ( .A(n_131), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_132), .A2(n_221), .B1(n_354), .B2(n_361), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_133), .Y(n_955) );
BUFx3_ASAP7_75t_L g360 ( .A(n_134), .Y(n_360) );
INVx1_ASAP7_75t_L g478 ( .A(n_135), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_136), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g1161 ( .A1(n_137), .A2(n_139), .B1(n_1149), .B2(n_1152), .Y(n_1161) );
INVx1_ASAP7_75t_L g451 ( .A(n_138), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_138), .A2(n_174), .B1(n_473), .B2(n_476), .C(n_477), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_140), .B(n_1127), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_142), .A2(n_205), .B1(n_1142), .B2(n_1146), .Y(n_1167) );
AOI221xp5_ASAP7_75t_L g1356 ( .A1(n_143), .A2(n_223), .B1(n_777), .B2(n_823), .C(n_835), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_143), .A2(n_195), .B1(n_752), .B2(n_755), .Y(n_1372) );
INVx1_ASAP7_75t_L g849 ( .A(n_144), .Y(n_849) );
OAI21xp33_ASAP7_75t_L g756 ( .A1(n_145), .A2(n_757), .B(n_758), .Y(n_756) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_146), .Y(n_255) );
INVx1_ASAP7_75t_L g439 ( .A(n_147), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_148), .A2(n_179), .B1(n_508), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_148), .A2(n_173), .B1(n_391), .B2(n_550), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_151), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_152), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_153), .A2(n_180), .B1(n_278), .B2(n_313), .C(n_315), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_153), .A2(n_186), .B1(n_368), .B2(n_370), .C(n_375), .Y(n_367) );
INVx1_ASAP7_75t_L g1047 ( .A(n_154), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_155), .A2(n_218), .B1(n_782), .B2(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g462 ( .A(n_157), .Y(n_462) );
INVx1_ASAP7_75t_L g761 ( .A(n_158), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g939 ( .A(n_159), .Y(n_939) );
INVx1_ASAP7_75t_L g596 ( .A(n_160), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_160), .B(n_420), .Y(n_598) );
INVx1_ASAP7_75t_L g1359 ( .A(n_161), .Y(n_1359) );
INVx1_ASAP7_75t_L g737 ( .A(n_162), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g684 ( .A1(n_163), .A2(n_476), .B(n_512), .Y(n_684) );
INVx1_ASAP7_75t_L g698 ( .A(n_163), .Y(n_698) );
INVx1_ASAP7_75t_L g983 ( .A(n_164), .Y(n_983) );
OAI211xp5_ASAP7_75t_L g1011 ( .A1(n_164), .A2(n_1012), .B(n_1014), .C(n_1016), .Y(n_1011) );
XOR2x2_ASAP7_75t_L g930 ( .A(n_165), .B(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g572 ( .A(n_166), .Y(n_572) );
OAI211xp5_ASAP7_75t_L g820 ( .A1(n_167), .A2(n_787), .B(n_821), .C(n_830), .Y(n_820) );
INVx1_ASAP7_75t_L g876 ( .A(n_167), .Y(n_876) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_168), .A2(n_220), .B1(n_835), .B2(n_836), .C(n_838), .Y(n_834) );
INVx1_ASAP7_75t_L g852 ( .A(n_168), .Y(n_852) );
INVxp67_ASAP7_75t_SL g1058 ( .A(n_169), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_169), .A2(n_193), .B1(n_702), .B2(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g845 ( .A(n_170), .Y(n_845) );
OAI332xp33_ASAP7_75t_SL g850 ( .A1(n_170), .A2(n_554), .A3(n_715), .B1(n_851), .B2(n_857), .B3(n_858), .C1(n_864), .C2(n_868), .Y(n_850) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_171), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_172), .A2(n_181), .B1(n_755), .B2(n_916), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_173), .A2(n_214), .B1(n_474), .B2(n_510), .C(n_512), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g468 ( .A1(n_174), .A2(n_384), .B(n_385), .Y(n_468) );
XOR2x2_ASAP7_75t_L g656 ( .A(n_175), .B(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_176), .A2(n_222), .B1(n_630), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g700 ( .A(n_176), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_177), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g888 ( .A(n_178), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_178), .A2(n_218), .B1(n_763), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_179), .A2(n_214), .B1(n_391), .B2(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_R g635 ( .A(n_182), .B(n_636), .Y(n_635) );
OA22x2_ASAP7_75t_L g880 ( .A1(n_184), .A2(n_881), .B1(n_923), .B2(n_924), .Y(n_880) );
CKINVDCx16_ASAP7_75t_R g923 ( .A(n_184), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_185), .A2(n_193), .B1(n_777), .B2(n_1051), .C(n_1052), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_186), .A2(n_192), .B1(n_282), .B2(n_286), .C(n_290), .Y(n_281) );
INVx1_ASAP7_75t_L g1117 ( .A(n_187), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_188), .Y(n_937) );
INVx1_ASAP7_75t_L g591 ( .A(n_189), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_190), .A2(n_209), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g867 ( .A(n_190), .Y(n_867) );
INVx1_ASAP7_75t_L g1088 ( .A(n_191), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_194), .A2(n_229), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_196), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_196), .A2(n_199), .B1(n_407), .B2(n_411), .C(n_414), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_197), .A2(n_227), .B1(n_380), .B2(n_742), .Y(n_741) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_197), .Y(n_797) );
OAI211xp5_ASAP7_75t_SL g445 ( .A1(n_198), .A2(n_401), .B(n_414), .C(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g489 ( .A(n_198), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_199), .A2(n_208), .B1(n_297), .B2(n_305), .C(n_310), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_200), .Y(n_670) );
INVx1_ASAP7_75t_L g842 ( .A(n_201), .Y(n_842) );
OAI211xp5_ASAP7_75t_L g1346 ( .A1(n_203), .A2(n_884), .B(n_1347), .C(n_1349), .Y(n_1346) );
INVx1_ASAP7_75t_L g1367 ( .A(n_203), .Y(n_1367) );
BUFx3_ASAP7_75t_L g258 ( .A(n_204), .Y(n_258) );
INVx1_ASAP7_75t_L g335 ( .A(n_204), .Y(n_335) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_206), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_207), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_208), .A2(n_210), .B1(n_393), .B2(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g854 ( .A(n_209), .Y(n_854) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_210), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_211), .Y(n_948) );
INVx1_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
INVx2_ASAP7_75t_L g300 ( .A(n_213), .Y(n_300) );
INVx1_ASAP7_75t_L g325 ( .A(n_213), .Y(n_325) );
INVx1_ASAP7_75t_L g479 ( .A(n_215), .Y(n_479) );
INVx1_ASAP7_75t_L g606 ( .A(n_216), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_216), .A2(n_233), .B1(n_508), .B2(n_515), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_217), .B(n_476), .Y(n_675) );
INVx1_ASAP7_75t_L g907 ( .A(n_219), .Y(n_907) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_220), .Y(n_865) );
INVx1_ASAP7_75t_L g316 ( .A(n_221), .Y(n_316) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_222), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_224), .Y(n_456) );
INVx1_ASAP7_75t_L g809 ( .A(n_225), .Y(n_809) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_228), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_230), .Y(n_669) );
INVx1_ASAP7_75t_L g681 ( .A(n_232), .Y(n_681) );
INVx1_ASAP7_75t_L g615 ( .A(n_233), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_259), .B(n_1133), .Y(n_234) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g1377 ( .A(n_238), .B(n_247), .Y(n_1377) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g1383 ( .A(n_240), .B(n_243), .Y(n_1383) );
INVx1_ASAP7_75t_L g1391 ( .A(n_240), .Y(n_1391) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g1393 ( .A(n_243), .B(n_1391), .Y(n_1393) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g1001 ( .A(n_247), .B(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g292 ( .A(n_248), .B(n_258), .Y(n_292) );
AND2x4_ASAP7_75t_L g513 ( .A(n_248), .B(n_257), .Y(n_513) );
INVx1_ASAP7_75t_L g997 ( .A(n_249), .Y(n_997) );
AND2x4_ASAP7_75t_SL g1376 ( .A(n_249), .B(n_1377), .Y(n_1376) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
OR2x6_ASAP7_75t_L g989 ( .A(n_251), .B(n_990), .Y(n_989) );
INVxp67_ASAP7_75t_L g1127 ( .A(n_251), .Y(n_1127) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
BUFx4f_ASAP7_75t_L g523 ( .A(n_252), .Y(n_523) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g277 ( .A(n_254), .Y(n_277) );
INVx2_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
NAND2x1_ASAP7_75t_L g289 ( .A(n_254), .B(n_255), .Y(n_289) );
INVx1_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
AND2x2_ASAP7_75t_L g433 ( .A(n_254), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g475 ( .A(n_254), .B(n_255), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_255), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g284 ( .A(n_255), .B(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g304 ( .A(n_255), .Y(n_304) );
INVx1_ASAP7_75t_L g329 ( .A(n_255), .Y(n_329) );
AND2x2_ASAP7_75t_L g338 ( .A(n_255), .B(n_277), .Y(n_338) );
INVx2_ASAP7_75t_L g434 ( .A(n_255), .Y(n_434) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g977 ( .A(n_257), .Y(n_977) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g981 ( .A(n_258), .Y(n_981) );
AND2x4_ASAP7_75t_L g985 ( .A(n_258), .B(n_307), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B1(n_812), .B2(n_1132), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
XNOR2x1_ASAP7_75t_L g262 ( .A(n_263), .B(n_496), .Y(n_262) );
BUFx2_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
XNOR2x1_ASAP7_75t_L g265 ( .A(n_266), .B(n_436), .Y(n_265) );
XNOR2x1_ASAP7_75t_L g266 ( .A(n_267), .B(n_435), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_351), .Y(n_267) );
NAND3xp33_ASAP7_75t_SL g268 ( .A(n_269), .B(n_321), .C(n_344), .Y(n_268) );
AOI211xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_281), .B(n_296), .C(n_312), .Y(n_269) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_272), .Y(n_1059) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g480 ( .A(n_274), .Y(n_480) );
INVx4_ASAP7_75t_L g673 ( .A(n_274), .Y(n_673) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_274), .Y(n_802) );
INVx8_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
OR2x2_ASAP7_75t_L g995 ( .A(n_275), .B(n_981), .Y(n_995) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_280), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
OAI22x1_ASAP7_75t_SL g483 ( .A1(n_280), .A2(n_456), .B1(n_480), .B2(n_484), .Y(n_483) );
INVx2_ASAP7_75t_SL g968 ( .A(n_280), .Y(n_968) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_287), .B1(n_316), .B2(n_317), .C(n_318), .Y(n_315) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g640 ( .A(n_284), .Y(n_640) );
BUFx2_ASAP7_75t_L g672 ( .A(n_284), .Y(n_672) );
BUFx2_ASAP7_75t_L g794 ( .A(n_284), .Y(n_794) );
AND2x2_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_285), .Y(n_530) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g790 ( .A1(n_287), .A2(n_513), .B1(n_791), .B2(n_792), .C(n_795), .Y(n_790) );
BUFx4f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x6_ASAP7_75t_L g310 ( .A(n_288), .B(n_311), .Y(n_310) );
INVx4_ASAP7_75t_L g525 ( .A(n_288), .Y(n_525) );
BUFx4f_ASAP7_75t_L g536 ( .A(n_288), .Y(n_536) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g342 ( .A(n_289), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_290), .A2(n_310), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x4_ASAP7_75t_L g485 ( .A(n_292), .B(n_486), .Y(n_485) );
INVx4_ASAP7_75t_L g519 ( .A(n_292), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_292), .B(n_675), .C(n_676), .D(n_678), .Y(n_674) );
INVx1_ASAP7_75t_SL g777 ( .A(n_292), .Y(n_777) );
INVx4_ASAP7_75t_L g898 ( .A(n_292), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_292), .B(n_486), .Y(n_972) );
INVx1_ASAP7_75t_L g487 ( .A(n_293), .Y(n_487) );
OR2x2_ASAP7_75t_L g570 ( .A(n_293), .B(n_396), .Y(n_570) );
OR2x2_ASAP7_75t_L g696 ( .A(n_293), .B(n_386), .Y(n_696) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_293), .Y(n_1036) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g309 ( .A(n_294), .Y(n_309) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g490 ( .A(n_297), .Y(n_490) );
INVx2_ASAP7_75t_SL g634 ( .A(n_297), .Y(n_634) );
NAND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_L g311 ( .A(n_298), .Y(n_311) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
BUFx2_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
INVx2_ASAP7_75t_L g427 ( .A(n_300), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_301), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_301), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g533 ( .A(n_301), .Y(n_533) );
AND2x6_ASAP7_75t_L g783 ( .A(n_301), .B(n_474), .Y(n_783) );
AND2x2_ASAP7_75t_L g840 ( .A(n_301), .B(n_527), .Y(n_840) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g527 ( .A(n_304), .Y(n_527) );
INVx1_ASAP7_75t_L g806 ( .A(n_304), .Y(n_806) );
AND2x4_ASAP7_75t_L g980 ( .A(n_304), .B(n_981), .Y(n_980) );
INVx1_ASAP7_75t_SL g632 ( .A(n_305), .Y(n_632) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
OR2x2_ASAP7_75t_L g492 ( .A(n_306), .B(n_309), .Y(n_492) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
INVxp67_ASAP7_75t_L g539 ( .A(n_309), .Y(n_539) );
INVx1_ASAP7_75t_L g1002 ( .A(n_309), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_310), .Y(n_495) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_318), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_318), .B(n_628), .Y(n_627) );
INVx4_ASAP7_75t_L g958 ( .A(n_318), .Y(n_958) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OR2x6_ASAP7_75t_L g554 ( .A(n_319), .B(n_375), .Y(n_554) );
INVx1_ASAP7_75t_L g653 ( .A(n_319), .Y(n_653) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_330), .B1(n_331), .B2(n_339), .C1(n_340), .C2(n_343), .Y(n_321) );
AOI21xp33_ASAP7_75t_SL g493 ( .A1(n_322), .A2(n_494), .B(n_495), .Y(n_493) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g557 ( .A(n_324), .B(n_404), .Y(n_557) );
OR2x2_ASAP7_75t_L g651 ( .A(n_324), .B(n_327), .Y(n_651) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_325), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g706 ( .A(n_325), .Y(n_706) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g350 ( .A(n_328), .B(n_334), .Y(n_350) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_328), .Y(n_507) );
INVx3_ASAP7_75t_L g516 ( .A(n_328), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g488 ( .A1(n_331), .A2(n_447), .B1(n_462), .B2(n_489), .C1(n_490), .C2(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g647 ( .A(n_331), .Y(n_647) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_336), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g341 ( .A(n_333), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g636 ( .A(n_333), .B(n_342), .Y(n_636) );
AND2x2_ASAP7_75t_L g431 ( .A(n_334), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g504 ( .A(n_334), .B(n_336), .Y(n_504) );
BUFx2_ASAP7_75t_L g534 ( .A(n_334), .Y(n_534) );
AND2x4_ASAP7_75t_SL g663 ( .A(n_334), .B(n_474), .Y(n_663) );
AND2x4_ASAP7_75t_L g769 ( .A(n_334), .B(n_432), .Y(n_769) );
AND2x4_ASAP7_75t_L g785 ( .A(n_334), .B(n_630), .Y(n_785) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_335), .Y(n_990) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g1055 ( .A(n_337), .Y(n_1055) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g508 ( .A(n_338), .Y(n_508) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_338), .Y(n_630) );
BUFx3_ASAP7_75t_L g782 ( .A(n_338), .Y(n_782) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_339), .A2(n_400), .B(n_406), .C(n_419), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g471 ( .A1(n_340), .A2(n_448), .B1(n_472), .B2(n_481), .C1(n_482), .C2(n_485), .Y(n_471) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g683 ( .A(n_342), .Y(n_683) );
BUFx2_ASAP7_75t_SL g969 ( .A(n_342), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_347), .B(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_348), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_348), .A2(n_430), .B1(n_595), .B2(n_596), .Y(n_594) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x4_ASAP7_75t_L g430 ( .A(n_349), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g768 ( .A(n_350), .Y(n_768) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_350), .Y(n_846) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_399), .B(n_425), .C(n_428), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_367), .B1(n_379), .B2(n_388), .C(n_392), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x6_ASAP7_75t_SL g420 ( .A(n_355), .B(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g568 ( .A(n_355), .Y(n_568) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_355), .Y(n_1095) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_356), .Y(n_548) );
BUFx8_ASAP7_75t_L g763 ( .A(n_356), .Y(n_763) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g374 ( .A(n_358), .Y(n_374) );
AND2x4_ASAP7_75t_L g372 ( .A(n_359), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_360), .Y(n_363) );
AND2x4_ASAP7_75t_L g369 ( .A(n_360), .B(n_365), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_360), .B(n_366), .Y(n_455) );
OR2x2_ASAP7_75t_L g602 ( .A(n_360), .B(n_374), .Y(n_602) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx12f_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
AND2x4_ASAP7_75t_L g424 ( .A(n_362), .B(n_422), .Y(n_424) );
INVx5_ASAP7_75t_L g746 ( .A(n_362), .Y(n_746) );
BUFx3_ASAP7_75t_L g921 ( .A(n_362), .Y(n_921) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_362), .Y(n_1073) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_363), .B(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_363), .Y(n_1020) );
INVx1_ASAP7_75t_L g413 ( .A(n_364), .Y(n_413) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g381 ( .A(n_369), .Y(n_381) );
AND2x2_ASAP7_75t_L g398 ( .A(n_369), .B(n_395), .Y(n_398) );
BUFx2_ASAP7_75t_L g545 ( .A(n_369), .Y(n_545) );
BUFx2_ASAP7_75t_L g563 ( .A(n_369), .Y(n_563) );
BUFx2_ASAP7_75t_L g755 ( .A(n_369), .Y(n_755) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_369), .B(n_377), .Y(n_1015) );
BUFx2_ASAP7_75t_L g1070 ( .A(n_369), .Y(n_1070) );
INVx8_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_371), .Y(n_458) );
INVx2_ASAP7_75t_L g577 ( .A(n_371), .Y(n_577) );
INVx3_ASAP7_75t_L g752 ( .A(n_371), .Y(n_752) );
INVx8_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
AND2x2_ASAP7_75t_L g394 ( .A(n_372), .B(n_395), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_372), .B(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g702 ( .A(n_372), .Y(n_702) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_372), .Y(n_711) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g460 ( .A(n_375), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND3x1_ASAP7_75t_L g705 ( .A(n_376), .B(n_377), .C(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g404 ( .A(n_377), .B(n_405), .Y(n_404) );
OR2x4_ASAP7_75t_L g1007 ( .A(n_377), .B(n_602), .Y(n_1007) );
INVx1_ASAP7_75t_L g1010 ( .A(n_377), .Y(n_1010) );
OR2x6_ASAP7_75t_L g1030 ( .A(n_377), .B(n_1031), .Y(n_1030) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp33_ASAP7_75t_SL g386 ( .A(n_378), .B(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g543 ( .A(n_378), .Y(n_543) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g552 ( .A(n_381), .Y(n_552) );
INVx1_ASAP7_75t_L g1077 ( .A(n_381), .Y(n_1077) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_383), .A2(n_451), .B1(n_452), .B2(n_456), .C(n_457), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_383), .A2(n_415), .B1(n_608), .B2(n_609), .C(n_610), .Y(n_607) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g612 ( .A(n_384), .Y(n_612) );
INVx5_ASAP7_75t_L g708 ( .A(n_384), .Y(n_708) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
AND3x4_ASAP7_75t_L g542 ( .A(n_387), .B(n_427), .C(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g610 ( .A(n_387), .B(n_543), .Y(n_610) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_387), .Y(n_1034) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g748 ( .A(n_391), .Y(n_748) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_394), .A2(n_398), .B1(n_439), .B2(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x6_ASAP7_75t_L g538 ( .A(n_403), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g646 ( .A(n_403), .B(n_539), .Y(n_646) );
AND2x6_ASAP7_75t_L g408 ( .A(n_404), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g412 ( .A(n_404), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g418 ( .A(n_404), .Y(n_418) );
INVx4_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_408), .A2(n_412), .B1(n_447), .B2(n_448), .Y(n_446) );
AND2x4_ASAP7_75t_SL g556 ( .A(n_409), .B(n_557), .Y(n_556) );
NAND2x1_ASAP7_75t_L g692 ( .A(n_409), .B(n_557), .Y(n_692) );
AND2x2_ASAP7_75t_L g733 ( .A(n_409), .B(n_557), .Y(n_733) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_409), .B(n_557), .Y(n_1080) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g560 ( .A(n_413), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_414), .A2(n_600), .B1(n_607), .B2(n_611), .C(n_616), .Y(n_599) );
OR2x6_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g872 ( .A(n_415), .Y(n_872) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
BUFx3_ASAP7_75t_L g950 ( .A(n_416), .Y(n_950) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_417), .Y(n_1023) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_422), .Y(n_623) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_424), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_425), .Y(n_686) );
INVx1_ASAP7_75t_L g1130 ( .A(n_425), .Y(n_1130) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21x1_ASAP7_75t_L g501 ( .A1(n_426), .A2(n_502), .B(n_537), .Y(n_501) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI31xp33_ASAP7_75t_SL g443 ( .A1(n_427), .A2(n_444), .A3(n_445), .B(n_449), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g597 ( .A1(n_427), .A2(n_598), .A3(n_599), .B(n_619), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_430), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g571 ( .A(n_430), .Y(n_571) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_432), .Y(n_776) );
INVx1_ASAP7_75t_L g837 ( .A(n_432), .Y(n_837) );
INVx2_ASAP7_75t_L g1113 ( .A(n_432), .Y(n_1113) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g476 ( .A(n_433), .Y(n_476) );
INVx2_ASAP7_75t_L g511 ( .A(n_433), .Y(n_511) );
AND2x4_ASAP7_75t_L g999 ( .A(n_433), .B(n_990), .Y(n_999) );
AOI211x1_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_440), .C(n_470), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_461), .C(n_463), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_452), .A2(n_681), .B1(n_708), .B2(n_709), .C(n_710), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_452), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g581 ( .A(n_453), .B(n_570), .Y(n_581) );
INVx1_ASAP7_75t_L g856 ( .A(n_453), .Y(n_856) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_454), .Y(n_605) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_455), .Y(n_1031) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_468), .C(n_469), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_465), .A2(n_617), .B(n_618), .Y(n_616) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g940 ( .A(n_466), .Y(n_940) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g575 ( .A(n_467), .B(n_570), .Y(n_575) );
INVx4_ASAP7_75t_L g863 ( .A(n_467), .Y(n_863) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_488), .C(n_493), .Y(n_470) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g679 ( .A(n_474), .Y(n_679) );
INVx1_ASAP7_75t_L g826 ( .A(n_474), .Y(n_826) );
BUFx6f_ASAP7_75t_L g835 ( .A(n_474), .Y(n_835) );
AND2x2_ASAP7_75t_L g976 ( .A(n_474), .B(n_977), .Y(n_976) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g774 ( .A(n_475), .Y(n_774) );
INVx1_ASAP7_75t_L g824 ( .A(n_476), .Y(n_824) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_476), .Y(n_897) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g757 ( .A(n_492), .B(n_575), .Y(n_757) );
AND2x4_ASAP7_75t_L g909 ( .A(n_492), .B(n_575), .Y(n_909) );
AO22x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_723), .B1(n_810), .B2(n_811), .Y(n_496) );
INVx1_ASAP7_75t_L g810 ( .A(n_497), .Y(n_810) );
XNOR2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_656), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_590), .B1(n_654), .B2(n_655), .Y(n_498) );
INVx1_ASAP7_75t_L g655 ( .A(n_499), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_583), .C(n_587), .Y(n_499) );
INVx1_ASAP7_75t_L g584 ( .A(n_501), .Y(n_584) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_504), .A2(n_769), .B1(n_842), .B2(n_843), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .B1(n_514), .B2(n_517), .Y(n_505) );
INVx3_ASAP7_75t_L g901 ( .A(n_507), .Y(n_901) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g518 ( .A(n_511), .Y(n_518) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g838 ( .A(n_513), .Y(n_838) );
INVx1_ASAP7_75t_L g890 ( .A(n_513), .Y(n_890) );
INVx2_ASAP7_75t_L g1062 ( .A(n_513), .Y(n_1062) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g677 ( .A(n_516), .Y(n_677) );
INVx2_ASAP7_75t_L g779 ( .A(n_516), .Y(n_779) );
INVx2_ASAP7_75t_L g828 ( .A(n_516), .Y(n_828) );
INVx1_ASAP7_75t_L g892 ( .A(n_516), .Y(n_892) );
INVx1_ASAP7_75t_L g1053 ( .A(n_518), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_518), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_532), .B1(n_534), .B2(n_535), .Y(n_520) );
INVx2_ASAP7_75t_SL g961 ( .A(n_522), .Y(n_961) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g666 ( .A(n_523), .Y(n_666) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_523), .Y(n_799) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g667 ( .A(n_525), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_529), .B2(n_531), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_527), .A2(n_529), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_528), .A2(n_556), .B1(n_558), .B2(n_561), .C(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_531), .A2(n_574), .B1(n_576), .B2(n_579), .C1(n_580), .C2(n_582), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_532), .A2(n_534), .B1(n_665), .B2(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NOR2x1_ASAP7_75t_L g805 ( .A(n_533), .B(n_806), .Y(n_805) );
OAI211xp5_ASAP7_75t_L g887 ( .A1(n_536), .A2(n_888), .B(n_889), .C(n_891), .Y(n_887) );
OAI211xp5_ASAP7_75t_L g1349 ( .A1(n_536), .A2(n_1350), .B(n_1351), .C(n_1352), .Y(n_1349) );
INVx5_ASAP7_75t_L g721 ( .A(n_538), .Y(n_721) );
INVx1_ASAP7_75t_L g585 ( .A(n_540), .Y(n_585) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_555), .Y(n_540) );
AOI33xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_544), .A3(n_546), .B1(n_549), .B2(n_551), .B3(n_553), .Y(n_541) );
BUFx3_ASAP7_75t_L g740 ( .A(n_542), .Y(n_740) );
AOI33xp33_ASAP7_75t_L g914 ( .A1(n_542), .A2(n_915), .A3(n_917), .B1(n_918), .B2(n_919), .B3(n_920), .Y(n_914) );
AOI33xp33_ASAP7_75t_L g1068 ( .A1(n_542), .A2(n_1069), .A3(n_1071), .B1(n_1074), .B2(n_1075), .B3(n_1076), .Y(n_1068) );
AOI33xp33_ASAP7_75t_L g1368 ( .A1(n_542), .A2(n_919), .A3(n_1369), .B1(n_1370), .B2(n_1371), .B3(n_1372), .Y(n_1368) );
INVx3_ASAP7_75t_L g1019 ( .A(n_543), .Y(n_1019) );
INVx2_ASAP7_75t_L g866 ( .A(n_547), .Y(n_866) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_548), .Y(n_550) );
INVx2_ASAP7_75t_L g943 ( .A(n_548), .Y(n_943) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_548), .B(n_1010), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_552), .A2(n_577), .B1(n_595), .B2(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_SL g919 ( .A(n_554), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_556), .A2(n_558), .B1(n_886), .B2(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_556), .A2(n_558), .B1(n_1348), .B2(n_1367), .Y(n_1366) );
AND2x4_ASAP7_75t_SL g558 ( .A(n_557), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g562 ( .A(n_557), .B(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g693 ( .A(n_557), .B(n_559), .Y(n_693) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g722 ( .A(n_562), .Y(n_722) );
INVx3_ASAP7_75t_L g738 ( .A(n_562), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_562), .B(n_911), .C(n_922), .Y(n_910) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_562), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_563), .Y(n_1092) );
INVx1_ASAP7_75t_L g589 ( .A(n_564), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_572), .Y(n_564) );
NAND2x1_ASAP7_75t_L g565 ( .A(n_566), .B(n_571), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVxp67_ASAP7_75t_L g718 ( .A(n_569), .Y(n_718) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g578 ( .A(n_570), .Y(n_578) );
INVx1_ASAP7_75t_L g588 ( .A(n_573), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_574), .A2(n_580), .B1(n_670), .B2(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x4_ASAP7_75t_L g760 ( .A(n_577), .B(n_578), .Y(n_760) );
AND2x4_ASAP7_75t_L g762 ( .A(n_578), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g728 ( .A(n_581), .B(n_651), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_586), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_586), .A2(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
XNOR2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_624), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B1(n_604), .B2(n_606), .Y(n_600) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_601), .Y(n_938) );
BUFx4f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g717 ( .A(n_602), .Y(n_717) );
BUFx3_ASAP7_75t_L g859 ( .A(n_602), .Y(n_859) );
BUFx3_ASAP7_75t_L g870 ( .A(n_602), .Y(n_870) );
OR2x4_ASAP7_75t_L g1028 ( .A(n_602), .B(n_1010), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_604), .A2(n_938), .B1(n_955), .B2(n_956), .Y(n_954) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g614 ( .A(n_605), .Y(n_614) );
INVx3_ASAP7_75t_L g699 ( .A(n_605), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_608), .A2(n_639), .B(n_641), .C(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_612), .A2(n_698), .B1(n_699), .B2(n_700), .C(n_701), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_614), .A2(n_942), .B1(n_943), .B2(n_944), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_621), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_643), .C(n_648), .Y(n_624) );
NOR3xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_635), .C(n_637), .Y(n_625) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_629), .B(n_631), .Y(n_626) );
BUFx2_ASAP7_75t_L g829 ( .A(n_630), .Y(n_829) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
BUFx2_ASAP7_75t_L g808 ( .A(n_653), .Y(n_808) );
INVx1_ASAP7_75t_L g1063 ( .A(n_653), .Y(n_1063) );
AND5x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_690), .C(n_712), .D(n_719), .E(n_722), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_686), .B(n_687), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .C(n_674), .D(n_680), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AOI221x1_ASAP7_75t_L g690 ( .A1(n_661), .A2(n_669), .B1(n_691), .B2(n_693), .C(n_694), .Y(n_690) );
BUFx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g789 ( .A(n_663), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_672), .A2(n_682), .B1(n_942), .B2(n_948), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_672), .A2(n_939), .B1(n_956), .B2(n_962), .Y(n_965) );
INVx2_ASAP7_75t_L g963 ( .A(n_673), .Y(n_963) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B(n_684), .C(n_685), .Y(n_680) );
INVx5_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_691), .A2(n_693), .B1(n_839), .B2(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AO22x1_ASAP7_75t_L g731 ( .A1(n_693), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_693), .A2(n_1079), .B1(n_1080), .B2(n_1081), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_693), .A2(n_733), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_697), .B1(n_703), .B2(n_707), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx8_ASAP7_75t_L g857 ( .A(n_696), .Y(n_857) );
BUFx4f_ASAP7_75t_L g935 ( .A(n_696), .Y(n_935) );
INVx2_ASAP7_75t_SL g743 ( .A(n_702), .Y(n_743) );
BUFx3_ASAP7_75t_L g916 ( .A(n_702), .Y(n_916) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g750 ( .A(n_705), .Y(n_750) );
INVx8_ASAP7_75t_L g947 ( .A(n_708), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
OR2x6_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_716), .B(n_718), .Y(n_1374) );
INVx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_721), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_721), .B(n_843), .Y(n_877) );
AND4x1_ASAP7_75t_L g1064 ( .A(n_722), .B(n_1065), .C(n_1068), .D(n_1078), .Y(n_1064) );
INVx2_ASAP7_75t_L g811 ( .A(n_723), .Y(n_811) );
XOR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_809), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_725), .B(n_764), .Y(n_724) );
AOI211x1_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_729), .C(n_756), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g906 ( .A1(n_727), .A2(n_907), .B(n_908), .Y(n_906) );
AOI21xp33_ASAP7_75t_L g1041 ( .A1(n_727), .A2(n_1042), .B(n_1043), .Y(n_1041) );
AOI21xp5_ASAP7_75t_L g1102 ( .A1(n_727), .A2(n_1103), .B(n_1104), .Y(n_1102) );
AOI21xp33_ASAP7_75t_L g1361 ( .A1(n_727), .A2(n_1362), .B(n_1363), .Y(n_1361) );
INVx8_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_739), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_736), .B(n_738), .Y(n_735) );
NAND2xp5_ASAP7_75t_R g784 ( .A(n_737), .B(n_785), .Y(n_784) );
NAND4xp25_ASAP7_75t_L g874 ( .A(n_738), .B(n_875), .C(n_877), .D(n_878), .Y(n_874) );
AOI33xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .A3(n_744), .B1(n_747), .B2(n_749), .B3(n_751), .Y(n_739) );
AOI33xp33_ASAP7_75t_L g1090 ( .A1(n_740), .A2(n_1091), .A3(n_1093), .B1(n_1096), .B2(n_1097), .B3(n_1098), .Y(n_1090) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
BUFx2_ASAP7_75t_L g953 ( .A(n_750), .Y(n_953) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_750), .Y(n_1075) );
BUFx2_ASAP7_75t_L g1097 ( .A(n_750), .Y(n_1097) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g848 ( .A(n_757), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_759), .A2(n_761), .B1(n_767), .B2(n_769), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_762), .B(n_842), .Y(n_878) );
INVx2_ASAP7_75t_L g1067 ( .A(n_762), .Y(n_1067) );
INVx2_ASAP7_75t_L g1100 ( .A(n_762), .Y(n_1100) );
INVx3_ASAP7_75t_L g853 ( .A(n_763), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_786), .B(n_807), .Y(n_764) );
NAND3xp33_ASAP7_75t_SL g765 ( .A(n_766), .B(n_770), .C(n_784), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_767), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_767), .A2(n_1117), .B1(n_1118), .B2(n_1119), .Y(n_1116) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_769), .Y(n_905) );
INVx1_ASAP7_75t_L g1120 ( .A(n_769), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_778), .B(n_783), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g1124 ( .A(n_773), .Y(n_1124) );
BUFx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
BUFx3_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
BUFx3_ASAP7_75t_L g1115 ( .A(n_782), .Y(n_1115) );
INVx1_ASAP7_75t_L g830 ( .A(n_783), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_783), .A2(n_896), .B(n_899), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g1049 ( .A1(n_783), .A2(n_1050), .B(n_1054), .Y(n_1049) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_783), .A2(n_1108), .B(n_1114), .Y(n_1107) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_783), .A2(n_1356), .B(n_1357), .Y(n_1355) );
INVx3_ASAP7_75t_L g894 ( .A(n_785), .Y(n_894) );
INVx2_ASAP7_75t_SL g1354 ( .A(n_785), .Y(n_1354) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g884 ( .A(n_788), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_788), .A2(n_805), .B1(n_1088), .B2(n_1089), .Y(n_1128) );
INVx4_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx4_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_800), .B2(n_801), .Y(n_796) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx5_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_807), .A2(n_820), .B(n_831), .Y(n_819) );
OAI21xp5_ASAP7_75t_SL g882 ( .A1(n_807), .A2(n_883), .B(n_893), .Y(n_882) );
OAI21xp5_ASAP7_75t_SL g1345 ( .A1(n_807), .A2(n_1346), .B(n_1353), .Y(n_1345) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_SL g1132 ( .A(n_812), .Y(n_1132) );
XNOR2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_926), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_880), .B2(n_925), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_874), .C(n_879), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_847), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_827), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1051 ( .A(n_826), .Y(n_1051) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_841), .C(n_844), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_839), .B2(n_840), .Y(n_832) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_835), .Y(n_1109) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_840), .B(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_840), .B(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_846), .A2(n_905), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_846), .A2(n_905), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B(n_850), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B1(n_854), .B2(n_855), .Y(n_851) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_861), .B2(n_862), .Y(n_858) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B1(n_871), .B2(n_873), .Y(n_868) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g925 ( .A(n_880), .Y(n_925) );
INVx1_ASAP7_75t_L g924 ( .A(n_881), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_906), .C(n_910), .Y(n_881) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_912), .B(n_914), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B1(n_1083), .B2(n_1131), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OA22x2_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_1037), .B2(n_1038), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_932), .B(n_973), .C(n_1003), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_957), .Y(n_932) );
OAI33xp33_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_936), .A3(n_941), .B1(n_945), .B2(n_952), .B3(n_954), .Y(n_933) );
BUFx3_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_937), .A2(n_955), .B1(n_960), .B2(n_962), .Y(n_959) );
INVx1_ASAP7_75t_L g1072 ( .A(n_943), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_944), .A2(n_951), .B1(n_967), .B2(n_969), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_948), .B1(n_949), .B2(n_951), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g1013 ( .A(n_950), .Y(n_1013) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
OAI33xp33_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_959), .A3(n_964), .B1(n_965), .B2(n_966), .B3(n_970), .Y(n_957) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_967), .A2(n_1058), .B1(n_1059), .B2(n_1060), .C(n_1061), .Y(n_1057) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
OAI31xp33_ASAP7_75t_SL g973 ( .A1(n_974), .A2(n_986), .A3(n_996), .B(n_1000), .Y(n_973) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_978) );
BUFx3_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_982), .A2(n_1017), .B1(n_1021), .B2(n_1024), .Y(n_1016) );
BUFx3_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx3_ASAP7_75t_SL g998 ( .A(n_999), .Y(n_998) );
BUFx3_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI31xp33_ASAP7_75t_SL g1003 ( .A1(n_1004), .A2(n_1011), .A3(n_1025), .B(n_1032), .Y(n_1003) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
CKINVDCx8_ASAP7_75t_R g1014 ( .A(n_1015), .Y(n_1014) );
BUFx3_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_1019), .B(n_1023), .Y(n_1022) );
BUFx6f_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1035), .Y(n_1032) );
INVx1_ASAP7_75t_SL g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
AO21x2_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1040), .B(n_1082), .Y(n_1038) );
NAND3xp33_ASAP7_75t_SL g1040 ( .A(n_1041), .B(n_1044), .C(n_1064), .Y(n_1040) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1056), .B(n_1063), .Y(n_1044) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_1083), .Y(n_1131) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1102), .C(n_1105), .Y(n_1084) );
NOR3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1099), .C(n_1101), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1090), .Y(n_1086) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
NOR3xp33_ASAP7_75t_L g1364 ( .A(n_1101), .B(n_1365), .C(n_1373), .Y(n_1364) );
OAI21xp5_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1121), .B(n_1129), .Y(n_1105) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1126), .Y(n_1122) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1338), .B1(n_1341), .B2(n_1375), .C(n_1378), .Y(n_1133) );
AND4x1_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1267), .C(n_1303), .D(n_1327), .Y(n_1134) );
NOR4xp25_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1208), .C(n_1230), .D(n_1244), .Y(n_1135) );
OAI211xp5_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1162), .B(n_1181), .C(n_1201), .Y(n_1136) );
OAI211xp5_ASAP7_75t_SL g1304 ( .A1(n_1137), .A2(n_1305), .B(n_1306), .C(n_1316), .Y(n_1304) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1154), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1139), .B(n_1158), .Y(n_1249) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1139), .Y(n_1262) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1140), .B(n_1190), .Y(n_1189) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1140), .B(n_1158), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1140), .B(n_1164), .Y(n_1237) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_1140), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1148), .Y(n_1140) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1142), .Y(n_1340) );
AND2x6_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1143), .B(n_1147), .Y(n_1146) );
AND2x4_ASAP7_75t_L g1149 ( .A(n_1143), .B(n_1150), .Y(n_1149) );
AND2x6_ASAP7_75t_L g1152 ( .A(n_1143), .B(n_1153), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1143), .B(n_1147), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1143), .B(n_1147), .Y(n_1301) );
OAI21xp5_ASAP7_75t_L g1390 ( .A1(n_1144), .A2(n_1391), .B(n_1392), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1145), .B(n_1151), .Y(n_1150) );
A2O1A1Ixp33_ASAP7_75t_L g1236 ( .A1(n_1154), .A2(n_1237), .B(n_1238), .C(n_1239), .Y(n_1236) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1154), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1158), .Y(n_1154) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1155), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1155), .B(n_1190), .Y(n_1212) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1155), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1155), .B(n_1237), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1155), .B(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1155), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_1158), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1158), .B(n_1192), .Y(n_1235) );
HB1xp67_ASAP7_75t_SL g1278 ( .A(n_1158), .Y(n_1278) );
OAI322xp33_ASAP7_75t_L g1332 ( .A1(n_1158), .A2(n_1163), .A3(n_1174), .B1(n_1194), .B2(n_1305), .C1(n_1319), .C2(n_1333), .Y(n_1332) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1161), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1168), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1163), .B(n_1216), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1163), .B(n_1308), .Y(n_1307) );
CKINVDCx14_ASAP7_75t_R g1163 ( .A(n_1164), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1164), .B(n_1194), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1164), .B(n_1216), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1164), .B(n_1186), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1164), .B(n_1243), .Y(n_1294) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1164), .B(n_1312), .Y(n_1320) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1164), .B(n_1242), .Y(n_1324) );
INVx3_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
CKINVDCx5p33_ASAP7_75t_R g1184 ( .A(n_1165), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1165), .B(n_1229), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1165), .B(n_1242), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1165), .B(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1165), .B(n_1170), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1331 ( .A(n_1165), .B(n_1218), .Y(n_1331) );
AND2x4_ASAP7_75t_SL g1165 ( .A(n_1166), .B(n_1167), .Y(n_1165) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1173), .Y(n_1169) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1170), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1170), .B(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1170), .B(n_1175), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1170), .B(n_1174), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1170), .B(n_1175), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1170), .B(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1173), .B(n_1186), .Y(n_1214) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1173), .Y(n_1246) );
OAI322xp33_ASAP7_75t_L g1272 ( .A1(n_1173), .A2(n_1223), .A3(n_1261), .B1(n_1273), .B2(n_1274), .C1(n_1275), .C2(n_1278), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1178), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1174), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1175), .B(n_1178), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1175), .B(n_1219), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1175), .B(n_1186), .Y(n_1225) );
NOR3xp33_ASAP7_75t_SL g1325 ( .A(n_1175), .B(n_1183), .C(n_1299), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1178), .Y(n_1197) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1178), .Y(n_1219) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1178), .Y(n_1298) );
NAND2x1_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
AOI221xp5_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1188), .B1(n_1191), .B2(n_1195), .C(n_1198), .Y(n_1181) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1182), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1185), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1183), .B(n_1214), .Y(n_1213) );
A2O1A1Ixp33_ASAP7_75t_L g1296 ( .A1(n_1183), .A2(n_1212), .B(n_1220), .C(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1184), .B(n_1188), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1184), .B(n_1254), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1184), .B(n_1196), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1184), .B(n_1249), .Y(n_1291) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1185), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1186), .B(n_1207), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1186), .B(n_1217), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1186), .B(n_1218), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1186), .B(n_1196), .Y(n_1269) );
NAND3xp33_ASAP7_75t_L g1284 ( .A(n_1186), .B(n_1285), .C(n_1287), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1186), .B(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1187), .Y(n_1207) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1188), .Y(n_1226) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1189), .B(n_1204), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1190), .B(n_1256), .Y(n_1255) );
HB1xp67_ASAP7_75t_SL g1274 ( .A(n_1190), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1190), .B(n_1243), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1193), .Y(n_1191) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1192), .Y(n_1204) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1192), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1192), .B(n_1271), .Y(n_1270) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OAI221xp5_ASAP7_75t_SL g1244 ( .A1(n_1194), .A2(n_1245), .B1(n_1249), .B2(n_1250), .C(n_1252), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1196), .B(n_1247), .Y(n_1251) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1196), .Y(n_1333) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1200), .Y(n_1198) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1199), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_1199), .A2(n_1211), .B1(n_1319), .B2(n_1321), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1205), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1204), .B(n_1299), .Y(n_1337) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
AOI21xp33_ASAP7_75t_L g1239 ( .A1(n_1206), .A2(n_1240), .B(n_1241), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1215), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1213), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1212), .B(n_1242), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1336 ( .A(n_1213), .Y(n_1336) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1214), .Y(n_1220) );
O2A1O1Ixp33_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1220), .B(n_1221), .C(n_1222), .Y(n_1215) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1216), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1217), .B(n_1266), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1286 ( .A(n_1217), .B(n_1246), .Y(n_1286) );
OAI21xp5_ASAP7_75t_SL g1313 ( .A1(n_1217), .A2(n_1294), .B(n_1297), .Y(n_1313) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AOI211xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1224), .B(n_1226), .C(n_1227), .Y(n_1222) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1223), .Y(n_1238) );
NOR2xp33_ASAP7_75t_L g1314 ( .A(n_1223), .B(n_1315), .Y(n_1314) );
CKINVDCx14_ASAP7_75t_R g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1229), .B(n_1262), .Y(n_1261) );
A2O1A1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1229), .A2(n_1281), .B(n_1282), .C(n_1283), .Y(n_1280) );
A2O1A1Ixp33_ASAP7_75t_L g1230 ( .A1(n_1231), .A2(n_1233), .B(n_1234), .C(n_1236), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
NAND3xp33_ASAP7_75t_L g1264 ( .A(n_1235), .B(n_1262), .C(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1238), .B(n_1262), .Y(n_1316) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_1240), .A2(n_1242), .B1(n_1298), .B2(n_1329), .C(n_1330), .Y(n_1328) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1241), .Y(n_1281) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1249), .Y(n_1271) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1249), .Y(n_1326) );
CKINVDCx14_ASAP7_75t_R g1250 ( .A(n_1251), .Y(n_1250) );
AOI221xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1255), .B1(n_1257), .B2(n_1260), .C(n_1263), .Y(n_1252) );
OAI31xp33_ASAP7_75t_L g1310 ( .A1(n_1256), .A2(n_1311), .A3(n_1312), .B(n_1313), .Y(n_1310) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1259), .Y(n_1282) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1262), .B(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI31xp33_ASAP7_75t_SL g1267 ( .A1(n_1268), .A2(n_1272), .A3(n_1279), .B(n_1299), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1269), .Y(n_1309) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
NAND4xp25_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1284), .C(n_1289), .D(n_1296), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
OAI21xp5_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1292), .B(n_1295), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVxp67_ASAP7_75t_SL g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1294), .Y(n_1329) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1297), .Y(n_1305) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1298), .B(n_1323), .Y(n_1322) );
INVx3_ASAP7_75t_L g1317 ( .A(n_1299), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1302), .Y(n_1299) );
AOI222xp33_ASAP7_75t_L g1303 ( .A1(n_1304), .A2(n_1317), .B1(n_1318), .B2(n_1325), .C1(n_1326), .C2(n_1395), .Y(n_1303) );
AOI211xp5_ASAP7_75t_L g1306 ( .A1(n_1307), .A2(n_1309), .B(n_1310), .C(n_1314), .Y(n_1306) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVxp67_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
OAI31xp33_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1332), .A3(n_1334), .B(n_1337), .Y(n_1327) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVxp67_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
CKINVDCx20_ASAP7_75t_R g1338 ( .A(n_1339), .Y(n_1338) );
CKINVDCx20_ASAP7_75t_R g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
HB1xp67_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1344), .Y(n_1388) );
NAND3xp33_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1361), .C(n_1364), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1368), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
BUFx3_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVxp33_ASAP7_75t_SL g1384 ( .A(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
endmodule