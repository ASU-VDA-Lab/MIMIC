module fake_jpeg_26929_n_323 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_22),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_32),
.B1(n_20),
.B2(n_36),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_60),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_31),
.C(n_34),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_76),
.C(n_34),
.Y(n_113)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_32),
.B1(n_20),
.B2(n_36),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_26),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_44),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_49),
.B1(n_48),
.B2(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_28),
.B1(n_26),
.B2(n_18),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_19),
.B1(n_27),
.B2(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_82),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_18),
.B(n_19),
.C(n_27),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_34),
.C(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_44),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_47),
.B1(n_29),
.B2(n_38),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_94),
.B1(n_95),
.B2(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_85),
.B(n_97),
.Y(n_145)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_90),
.Y(n_126)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_93),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_21),
.B1(n_22),
.B2(n_35),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_103),
.B(n_118),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_76),
.A3(n_81),
.B1(n_78),
.B2(n_47),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_105),
.B(n_74),
.C(n_63),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_35),
.A3(n_45),
.B1(n_57),
.B2(n_72),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_21),
.B1(n_23),
.B2(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_111),
.B1(n_54),
.B2(n_52),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_23),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_67),
.Y(n_129)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_9),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_137),
.C(n_100),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_122),
.A2(n_129),
.B(n_132),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_98),
.B1(n_96),
.B2(n_90),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_33),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_1),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_119),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_153),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_0),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_62),
.B1(n_33),
.B2(n_2),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_142),
.B1(n_150),
.B2(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_86),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_88),
.B(n_11),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_83),
.A2(n_62),
.B1(n_33),
.B2(n_11),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_101),
.Y(n_147)
);

OR2x2_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_16),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_85),
.B(n_7),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_62),
.B1(n_6),
.B2(n_12),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_0),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_6),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_167),
.B(n_123),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_151),
.B1(n_124),
.B2(n_152),
.Y(n_208)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_168),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_113),
.B(n_100),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_93),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_184),
.Y(n_203)
);

INVxp33_ASAP7_75t_SL g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

BUFx16f_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_147),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_181),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_121),
.A2(n_117),
.B1(n_89),
.B2(n_92),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_142),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_121),
.A2(n_117),
.B1(n_87),
.B2(n_13),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_5),
.B1(n_15),
.B2(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_180),
.A2(n_182),
.B1(n_188),
.B2(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_5),
.B1(n_15),
.B2(n_14),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_12),
.C(n_16),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_150),
.C(n_141),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_2),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_16),
.Y(n_199)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_145),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_199),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_200),
.B(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_197),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_129),
.C(n_146),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_184),
.C(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_157),
.A2(n_128),
.B(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_209),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_153),
.B1(n_135),
.B2(n_139),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_139),
.B1(n_155),
.B2(n_120),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_164),
.B(n_124),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_143),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_217),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_209),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_161),
.A2(n_3),
.B1(n_4),
.B2(n_188),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_172),
.B1(n_204),
.B2(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_3),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_3),
.B1(n_4),
.B2(n_156),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_179),
.B1(n_183),
.B2(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_213),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_235),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_167),
.B(n_174),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_239),
.B(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_225),
.B1(n_202),
.B2(n_207),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_173),
.B1(n_165),
.B2(n_166),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_229),
.C(n_233),
.Y(n_246)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_160),
.A3(n_185),
.B1(n_187),
.B2(n_169),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_159),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_213),
.B1(n_199),
.B2(n_210),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_196),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_190),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_205),
.B1(n_192),
.B2(n_214),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_213),
.B1(n_232),
.B2(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_194),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_243),
.B(n_259),
.Y(n_275)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_201),
.C(n_210),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_225),
.C(n_227),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_208),
.B1(n_207),
.B2(n_194),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_256),
.B1(n_260),
.B2(n_221),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_255),
.B(n_239),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_242),
.Y(n_267)
);

NAND2x1p5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_191),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_213),
.B(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_262),
.B(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_265),
.C(n_249),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_229),
.C(n_219),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_260),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_228),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_232),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_248),
.B1(n_247),
.B2(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_265),
.C(n_262),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_248),
.B1(n_243),
.B2(n_221),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_276),
.B(n_244),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_284),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_236),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_268),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_257),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_275),
.B1(n_271),
.B2(n_254),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_298),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_282),
.B(n_274),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_282),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_269),
.C(n_264),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_280),
.C(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_252),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_252),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_291),
.B1(n_286),
.B2(n_223),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_295),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_292),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_290),
.B(n_267),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_297),
.C(n_290),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_314),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_309),
.C(n_304),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

OAI21x1_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_311),
.B(n_250),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_321),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_319),
.Y(n_323)
);


endmodule