module fake_jpeg_15097_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_26),
.B1(n_18),
.B2(n_19),
.Y(n_66)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_17),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_16),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_61),
.B1(n_66),
.B2(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_57),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_66),
.Y(n_71)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_19),
.B1(n_16),
.B2(n_3),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_19),
.A3(n_18),
.B1(n_16),
.B2(n_42),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_66),
.B1(n_62),
.B2(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_48),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_19),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_88),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_80),
.B1(n_73),
.B2(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_66),
.B(n_25),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_16),
.B(n_59),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_106),
.B1(n_103),
.B2(n_97),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_93),
.A3(n_84),
.B1(n_83),
.B2(n_89),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_94),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_79),
.A3(n_41),
.B1(n_70),
.B2(n_82),
.C1(n_78),
.C2(n_47),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_82),
.B(n_2),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_115),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_1),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_90),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_44),
.C(n_4),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_88),
.B(n_85),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_55),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_11),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_10),
.B1(n_11),
.B2(n_5),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_100),
.B1(n_51),
.B2(n_3),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_124),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_113),
.B1(n_116),
.B2(n_114),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_124),
.B(n_123),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_140),
.B(n_6),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_SL g140 ( 
.A(n_137),
.B(n_127),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_139),
.A2(n_136),
.B(n_112),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_142),
.B(n_6),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_6),
.Y(n_145)
);


endmodule