module fake_jpeg_119_n_600 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_600);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_600;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_1),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_57),
.B(n_68),
.Y(n_139)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g180 ( 
.A(n_61),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_64),
.Y(n_127)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_16),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_85),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_15),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_86),
.B(n_87),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_26),
.B(n_15),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_12),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_92),
.B(n_113),
.Y(n_178)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_12),
.C(n_10),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_41),
.C(n_46),
.Y(n_156)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_52),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_35),
.B(n_12),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_18),
.Y(n_114)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_10),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_9),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_18),
.B1(n_33),
.B2(n_50),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_120),
.A2(n_132),
.B1(n_147),
.B2(n_164),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_44),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_122),
.B(n_153),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_64),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_125),
.B(n_136),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_18),
.B1(n_33),
.B2(n_50),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_97),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_59),
.A2(n_52),
.B1(n_46),
.B2(n_41),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_176),
.B1(n_179),
.B2(n_192),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_17),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_155),
.B(n_165),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_159),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_42),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_61),
.B(n_30),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_90),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_167),
.B(n_185),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_69),
.A2(n_17),
.B1(n_53),
.B2(n_42),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_91),
.A2(n_53),
.B1(n_38),
.B2(n_52),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_177),
.A2(n_38),
.B1(n_36),
.B2(n_28),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_60),
.A2(n_38),
.B1(n_40),
.B2(n_56),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_65),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_62),
.A2(n_38),
.B1(n_40),
.B2(n_56),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_94),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_193),
.B(n_206),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_144),
.A2(n_112),
.B1(n_74),
.B2(n_111),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_194),
.Y(n_273)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_197),
.Y(n_302)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_199),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_139),
.A2(n_85),
.B1(n_66),
.B2(n_70),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_204),
.A2(n_222),
.B1(n_230),
.B2(n_121),
.Y(n_271)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_106),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_100),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_213),
.Y(n_269)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_211),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_103),
.C(n_101),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_212),
.B(n_258),
.C(n_120),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_0),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_214),
.B(n_235),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_172),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_245),
.Y(n_275)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_218),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_164),
.A2(n_84),
.B1(n_63),
.B2(n_104),
.Y(n_222)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_172),
.A2(n_76),
.B1(n_61),
.B2(n_72),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g303 ( 
.A(n_228),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_132),
.A2(n_72),
.B1(n_38),
.B2(n_36),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_232),
.A2(n_255),
.B1(n_257),
.B2(n_261),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_233),
.A2(n_147),
.B1(n_259),
.B2(n_230),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_161),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_177),
.A2(n_28),
.B1(n_45),
.B2(n_10),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_238),
.A2(n_150),
.B1(n_142),
.B2(n_149),
.Y(n_288)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_118),
.Y(n_240)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_118),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_244),
.B(n_250),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_166),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_246),
.Y(n_284)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_247),
.B(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_248),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_190),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_251),
.Y(n_305)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_148),
.A2(n_81),
.B1(n_79),
.B2(n_45),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_131),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_259),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_152),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_123),
.B(n_0),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_180),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_129),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_271),
.A2(n_308),
.B1(n_202),
.B2(n_224),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_286),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_195),
.A2(n_142),
.B1(n_130),
.B2(n_128),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_278),
.A2(n_309),
.B1(n_197),
.B2(n_219),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_135),
.C(n_133),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_319),
.C(n_244),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_217),
.A2(n_9),
.B(n_149),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_296),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_288),
.A2(n_8),
.B1(n_272),
.B2(n_273),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_190),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_293),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_173),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_252),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_254),
.A2(n_150),
.B(n_134),
.C(n_173),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_320),
.B(n_266),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_217),
.B(n_2),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_206),
.A2(n_145),
.B1(n_141),
.B2(n_137),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_210),
.A2(n_183),
.B1(n_134),
.B2(n_141),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_213),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_209),
.B(n_183),
.C(n_145),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_253),
.A2(n_137),
.B1(n_4),
.B2(n_5),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_196),
.B(n_3),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_3),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_263),
.B(n_198),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_323),
.B(n_328),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_324),
.Y(n_386)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_327),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_263),
.B(n_212),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_312),
.A2(n_254),
.B(n_225),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_329),
.A2(n_321),
.B(n_295),
.Y(n_374)
);

AO22x1_ASAP7_75t_SL g330 ( 
.A1(n_301),
.A2(n_254),
.B1(n_258),
.B2(n_205),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_351),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_281),
.A2(n_254),
.B1(n_199),
.B2(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_332),
.Y(n_380)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_335),
.A2(n_338),
.B1(n_340),
.B2(n_346),
.Y(n_376)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_337),
.A2(n_358),
.B1(n_279),
.B2(n_297),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_271),
.A2(n_234),
.B1(n_200),
.B2(n_231),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_269),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_342),
.C(n_368),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_278),
.A2(n_247),
.B1(n_220),
.B2(n_241),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_305),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_344),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_290),
.A2(n_250),
.B1(n_240),
.B2(n_239),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_345),
.A2(n_356),
.B1(n_285),
.B2(n_268),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_301),
.A2(n_216),
.B1(n_201),
.B2(n_203),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_281),
.A2(n_232),
.B1(n_243),
.B2(n_246),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_347),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_273),
.A2(n_228),
.B1(n_211),
.B2(n_218),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_348),
.A2(n_363),
.B(n_321),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_269),
.B(n_4),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_368),
.Y(n_412)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_293),
.A2(n_223),
.B1(n_5),
.B2(n_6),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_366),
.B1(n_370),
.B2(n_311),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_274),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g381 ( 
.A1(n_354),
.A2(n_359),
.B1(n_310),
.B2(n_295),
.Y(n_381)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_356)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_286),
.A2(n_8),
.B1(n_319),
.B2(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_364),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_315),
.A2(n_275),
.B(n_306),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_300),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_367),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_286),
.A2(n_309),
.B1(n_320),
.B2(n_280),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_276),
.B(n_299),
.C(n_313),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_294),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_362),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_286),
.A2(n_268),
.B1(n_297),
.B2(n_265),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_374),
.A2(n_406),
.B(n_341),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_334),
.A2(n_294),
.B(n_292),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_395),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_285),
.B(n_264),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_292),
.C(n_291),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_342),
.C(n_369),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_392),
.A2(n_393),
.B1(n_340),
.B2(n_338),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_359),
.A2(n_302),
.B1(n_304),
.B2(n_270),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_302),
.B1(n_270),
.B2(n_300),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_394),
.A2(n_399),
.B1(n_401),
.B2(n_356),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_324),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_334),
.A2(n_279),
.B1(n_311),
.B2(n_291),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_404),
.B1(n_408),
.B2(n_345),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_298),
.B1(n_289),
.B2(n_318),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_357),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_410),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_346),
.A2(n_298),
.B1(n_289),
.B2(n_318),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_370),
.A2(n_303),
.B1(n_310),
.B2(n_328),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_329),
.A2(n_363),
.B(n_325),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_337),
.A2(n_344),
.B1(n_364),
.B2(n_360),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_352),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_323),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_412),
.B(n_325),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_413),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_391),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_414),
.B(n_416),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_391),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_418),
.A2(n_421),
.B1(n_424),
.B2(n_427),
.Y(n_465)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_382),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_425),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_330),
.B1(n_335),
.B2(n_331),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_423),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_383),
.A2(n_330),
.B1(n_331),
.B2(n_349),
.Y(n_424)
);

INVx5_ASAP7_75t_SL g425 ( 
.A(n_400),
.Y(n_425)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_383),
.A2(n_330),
.B1(n_354),
.B2(n_348),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_429),
.A2(n_438),
.B1(n_440),
.B2(n_377),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_373),
.B(n_326),
.Y(n_431)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_373),
.B(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_433),
.A2(n_434),
.B(n_372),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_383),
.A2(n_333),
.B(n_336),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_412),
.Y(n_435)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_382),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_439),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_376),
.A2(n_355),
.B1(n_343),
.B2(n_350),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_405),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_376),
.A2(n_327),
.B1(n_357),
.B2(n_353),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_385),
.B(n_367),
.C(n_361),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_446),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_385),
.B(n_390),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_446),
.B(n_422),
.Y(n_456)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_393),
.A2(n_365),
.B1(n_396),
.B2(n_387),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_449),
.A2(n_394),
.B1(n_399),
.B2(n_374),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_476),
.B(n_479),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_456),
.C(n_444),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_455),
.A2(n_474),
.B1(n_480),
.B2(n_415),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_443),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_459),
.B(n_457),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_379),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_473),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_470),
.B1(n_448),
.B2(n_449),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_423),
.B(n_432),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_467),
.B(n_472),
.Y(n_496)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_417),
.A2(n_380),
.B1(n_406),
.B2(n_410),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_445),
.B(n_377),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_424),
.B(n_375),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_421),
.A2(n_380),
.B1(n_401),
.B2(n_381),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_434),
.A2(n_380),
.B(n_378),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_441),
.A2(n_384),
.B(n_395),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_417),
.A2(n_381),
.B1(n_378),
.B2(n_384),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_483),
.A2(n_494),
.B1(n_499),
.B2(n_500),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_458),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_484),
.B(n_505),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_486),
.A2(n_474),
.B1(n_480),
.B2(n_466),
.Y(n_511)
);

AND3x1_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_415),
.C(n_416),
.Y(n_487)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

MAJx2_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_498),
.C(n_501),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_460),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_495),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_414),
.Y(n_491)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_491),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_420),
.C(n_437),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_493),
.C(n_508),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_433),
.C(n_386),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_465),
.A2(n_429),
.B1(n_419),
.B2(n_427),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_477),
.B(n_375),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_438),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_469),
.A2(n_440),
.B1(n_426),
.B2(n_418),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_469),
.A2(n_384),
.B1(n_425),
.B2(n_439),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_451),
.B(n_447),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_503),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_472),
.B(n_381),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_504),
.B(n_485),
.Y(n_512)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_478),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_453),
.B(n_398),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_507),
.Y(n_521)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_452),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_461),
.B(n_386),
.C(n_405),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_518),
.B1(n_528),
.B2(n_502),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_520),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_494),
.A2(n_470),
.B1(n_462),
.B2(n_476),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_513),
.A2(n_519),
.B1(n_504),
.B2(n_505),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_517),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_492),
.B(n_467),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_483),
.A2(n_464),
.B1(n_473),
.B2(n_436),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_496),
.B(n_450),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_463),
.Y(n_523)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_523),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_479),
.C(n_455),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_524),
.B(n_529),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_488),
.A2(n_487),
.B(n_484),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_488),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_491),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_493),
.B(n_407),
.C(n_398),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_407),
.C(n_402),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_496),
.C(n_508),
.Y(n_537)
);

XNOR2x1_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_548),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_536),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_509),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_539),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_540),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_485),
.C(n_500),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_499),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_525),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_544),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_482),
.C(n_471),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_542),
.B(n_549),
.C(n_514),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_464),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_507),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_514),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_518),
.B(n_497),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_547),
.B(n_521),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_513),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_481),
.C(n_471),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_522),
.A2(n_497),
.B1(n_481),
.B2(n_381),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_550),
.A2(n_519),
.B1(n_526),
.B2(n_528),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_552),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_561),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_526),
.Y(n_556)
);

OAI21x1_ASAP7_75t_SL g578 ( 
.A1(n_556),
.A2(n_538),
.B(n_402),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_559),
.B(n_564),
.Y(n_569)
);

XNOR2x1_ASAP7_75t_L g560 ( 
.A(n_538),
.B(n_520),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_565),
.Y(n_574)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_562),
.B(n_563),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_545),
.A2(n_522),
.B1(n_515),
.B2(n_531),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_511),
.C(n_531),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_517),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_542),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_546),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_532),
.C(n_539),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_568),
.B(n_571),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_554),
.A2(n_510),
.B1(n_548),
.B2(n_425),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_570),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_555),
.A2(n_510),
.B(n_537),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_572),
.A2(n_578),
.B(n_556),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_551),
.B(n_541),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_577),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_549),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_568),
.B(n_557),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_579),
.B(n_586),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_SL g588 ( 
.A(n_580),
.B(n_567),
.C(n_573),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_557),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_584),
.B(n_585),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_576),
.B(n_564),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_569),
.B(n_554),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_588),
.A2(n_589),
.B(n_591),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_582),
.A2(n_576),
.B(n_558),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_581),
.A2(n_570),
.B(n_558),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_590),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_592),
.B(n_594),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_587),
.A2(n_583),
.B(n_560),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_593),
.B(n_583),
.C(n_430),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_596),
.A2(n_595),
.B(n_403),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_597),
.A2(n_403),
.B(n_430),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_L g599 ( 
.A(n_598),
.B(n_442),
.C(n_389),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_442),
.Y(n_600)
);


endmodule