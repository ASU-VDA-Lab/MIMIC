module fake_jpeg_4578_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_16),
.B1(n_20),
.B2(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_17),
.B(n_13),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_13),
.B1(n_17),
.B2(n_10),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_41),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_35),
.B1(n_40),
.B2(n_22),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_58),
.B1(n_35),
.B2(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_48),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_29),
.B1(n_34),
.B2(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_59),
.C(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_55),
.C(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_56),
.B(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_68),
.B1(n_58),
.B2(n_36),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_83),
.B1(n_73),
.B2(n_70),
.Y(n_87)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_27),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_25),
.A3(n_24),
.B1(n_18),
.B2(n_11),
.C(n_13),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_72),
.B1(n_10),
.B2(n_8),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_2),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_8),
.C(n_4),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_93),
.C(n_84),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_7),
.Y(n_93)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_93),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_82),
.C(n_4),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_3),
.C(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_92),
.B1(n_82),
.B2(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_101),
.B(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

NAND2x1p5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_101),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_3),
.B(n_5),
.Y(n_108)
);

OA21x2_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_5),
.B(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_106),
.Y(n_110)
);


endmodule