module real_aes_6162_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_87), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g439 ( .A(n_0), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_1), .A2(n_144), .B(n_149), .C(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_2), .A2(n_139), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g457 ( .A(n_3), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_4), .B(n_163), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_5), .A2(n_104), .B1(n_112), .B2(n_732), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_6), .A2(n_16), .B1(n_720), .B2(n_721), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_6), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_7), .A2(n_139), .B(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_L g144 ( .A(n_8), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g173 ( .A(n_9), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_10), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_10), .B(n_44), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_11), .A2(n_251), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_12), .B(n_154), .Y(n_190) );
INVx1_ASAP7_75t_L g479 ( .A(n_13), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_14), .B(n_153), .Y(n_527) );
INVx1_ASAP7_75t_L g137 ( .A(n_15), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_16), .Y(n_720) );
INVx1_ASAP7_75t_L g539 ( .A(n_17), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_18), .A2(n_174), .B(n_199), .C(n_201), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_19), .B(n_163), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_20), .B(n_468), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_21), .B(n_139), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_22), .B(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_23), .A2(n_153), .B(n_155), .C(n_159), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_24), .B(n_163), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_25), .B(n_154), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_26), .A2(n_157), .B(n_201), .C(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_27), .B(n_154), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_28), .Y(n_219) );
INVx1_ASAP7_75t_L g233 ( .A(n_29), .Y(n_233) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_30), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_31), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_32), .B(n_154), .Y(n_458) );
INVx1_ASAP7_75t_L g256 ( .A(n_33), .Y(n_256) );
INVx1_ASAP7_75t_L g492 ( .A(n_34), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_35), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g142 ( .A(n_36), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_37), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_38), .A2(n_153), .B(n_212), .C(n_214), .Y(n_211) );
INVxp67_ASAP7_75t_L g257 ( .A(n_39), .Y(n_257) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_40), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_41), .A2(n_149), .B(n_232), .C(n_238), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_42), .A2(n_144), .B(n_149), .C(n_507), .Y(n_506) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_43), .A2(n_92), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_43), .Y(n_123) );
INVx1_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
INVx1_ASAP7_75t_L g491 ( .A(n_45), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_46), .A2(n_171), .B(n_172), .C(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_47), .B(n_154), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_48), .A2(n_120), .B1(n_432), .B2(n_433), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_48), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_49), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_50), .Y(n_253) );
INVx1_ASAP7_75t_L g147 ( .A(n_51), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_52), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_53), .B(n_139), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_54), .A2(n_149), .B1(n_159), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_55), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_56), .Y(n_454) );
CKINVDCx14_ASAP7_75t_R g169 ( .A(n_57), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_58), .A2(n_171), .B(n_214), .C(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_59), .Y(n_520) );
INVx1_ASAP7_75t_L g476 ( .A(n_60), .Y(n_476) );
INVx1_ASAP7_75t_L g145 ( .A(n_61), .Y(n_145) );
INVx1_ASAP7_75t_L g136 ( .A(n_62), .Y(n_136) );
INVx1_ASAP7_75t_SL g213 ( .A(n_63), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_65), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g222 ( .A(n_66), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_SL g467 ( .A1(n_67), .A2(n_214), .B(n_468), .C(n_469), .Y(n_467) );
INVxp67_ASAP7_75t_L g470 ( .A(n_68), .Y(n_470) );
INVx1_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_70), .A2(n_139), .B(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_71), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_72), .A2(n_139), .B(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_73), .Y(n_495) );
INVx1_ASAP7_75t_L g514 ( .A(n_74), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_75), .A2(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g197 ( .A(n_76), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_77), .Y(n_230) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_78), .A2(n_445), .B1(n_717), .B2(n_723), .C1(n_727), .C2(n_728), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_79), .A2(n_144), .B(n_149), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_80), .A2(n_139), .B(n_146), .Y(n_138) );
INVx1_ASAP7_75t_L g200 ( .A(n_81), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_82), .B(n_234), .Y(n_508) );
INVx2_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g187 ( .A(n_84), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_85), .B(n_468), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_86), .A2(n_144), .B(n_149), .C(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g436 ( .A(n_87), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g715 ( .A(n_87), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_87), .B(n_438), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_88), .A2(n_149), .B(n_221), .C(n_224), .Y(n_220) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_89), .A2(n_718), .B1(n_719), .B2(n_722), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_89), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_90), .B(n_166), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_91), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_92), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_93), .A2(n_144), .B(n_149), .C(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_94), .Y(n_531) );
INVx1_ASAP7_75t_L g466 ( .A(n_95), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_96), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_97), .B(n_234), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_98), .B(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_99), .B(n_132), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_100), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g156 ( .A(n_101), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_102), .A2(n_139), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g732 ( .A(n_104), .Y(n_732) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO21x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_443), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g731 ( .A(n_115), .Y(n_731) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_434), .B(n_441), .Y(n_118) );
INVx1_ASAP7_75t_L g433 ( .A(n_120), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B1(n_430), .B2(n_431), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_121), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_124), .A2(n_714), .B1(n_724), .B2(n_725), .Y(n_723) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g431 ( .A(n_125), .Y(n_431) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_356), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_298), .C(n_328), .D(n_338), .Y(n_126) );
OAI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_203), .B(n_261), .C(n_288), .Y(n_127) );
OAI222xp33_ASAP7_75t_L g383 ( .A1(n_128), .A2(n_303), .B1(n_384), .B2(n_385), .C1(n_386), .C2(n_387), .Y(n_383) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_178), .Y(n_128) );
AOI33xp33_ASAP7_75t_L g309 ( .A1(n_129), .A2(n_296), .A3(n_297), .B1(n_310), .B2(n_315), .B3(n_317), .Y(n_309) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_129), .A2(n_367), .B(n_369), .C(n_371), .Y(n_366) );
OR2x2_ASAP7_75t_L g382 ( .A(n_129), .B(n_368), .Y(n_382) );
INVx1_ASAP7_75t_L g415 ( .A(n_129), .Y(n_415) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
INVx2_ASAP7_75t_L g292 ( .A(n_130), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_130), .B(n_194), .Y(n_308) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_130), .Y(n_343) );
AND2x2_ASAP7_75t_L g372 ( .A(n_130), .B(n_165), .Y(n_372) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_162), .Y(n_130) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_131), .A2(n_195), .B(n_202), .Y(n_194) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_131), .A2(n_208), .B(n_216), .Y(n_207) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_132), .A2(n_464), .B(n_471), .Y(n_463) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g249 ( .A(n_133), .Y(n_249) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_134), .B(n_135), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx2_ASAP7_75t_L g251 ( .A(n_139), .Y(n_251) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_140), .B(n_144), .Y(n_184) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g237 ( .A(n_141), .Y(n_237) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
INVx1_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
INVx1_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
INVx3_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVx1_ASAP7_75t_L g468 ( .A(n_143), .Y(n_468) );
INVx4_ASAP7_75t_SL g161 ( .A(n_144), .Y(n_161) );
BUFx3_ASAP7_75t_L g238 ( .A(n_144), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_148), .B(n_152), .C(n_161), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_148), .A2(n_161), .B(n_169), .C(n_170), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g196 ( .A1(n_148), .A2(n_161), .B(n_197), .C(n_198), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_148), .A2(n_161), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_148), .A2(n_161), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_148), .A2(n_161), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_148), .A2(n_161), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_148), .A2(n_161), .B(n_536), .C(n_537), .Y(n_535) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx3_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_153), .B(n_213), .Y(n_212) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_157), .B(n_200), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_157), .A2(n_234), .B1(n_256), .B2(n_257), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_157), .B(n_539), .Y(n_538) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_158), .A2(n_189), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g459 ( .A(n_159), .Y(n_459) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_161), .A2(n_184), .B1(n_489), .B2(n_493), .Y(n_488) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_163), .A2(n_474), .B(n_480), .Y(n_473) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_164), .B(n_193), .Y(n_192) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_164), .A2(n_218), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_164), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_164), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g272 ( .A(n_165), .Y(n_272) );
BUFx3_ASAP7_75t_L g280 ( .A(n_165), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_165), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g291 ( .A(n_165), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_165), .B(n_179), .Y(n_320) );
AND2x2_ASAP7_75t_L g389 ( .A(n_165), .B(n_323), .Y(n_389) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_177), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx2_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_166), .A2(n_184), .B(n_230), .C(n_231), .Y(n_229) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_166), .A2(n_534), .B(n_540), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx5_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_174), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_174), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
INVx2_ASAP7_75t_SL g283 ( .A(n_178), .Y(n_283) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_194), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_179), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g325 ( .A(n_179), .Y(n_325) );
AND2x2_ASAP7_75t_L g336 ( .A(n_179), .B(n_292), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_179), .B(n_321), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_179), .B(n_323), .Y(n_368) );
AND2x2_ASAP7_75t_L g427 ( .A(n_179), .B(n_372), .Y(n_427) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g297 ( .A(n_180), .B(n_194), .Y(n_297) );
AND2x2_ASAP7_75t_L g307 ( .A(n_180), .B(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g329 ( .A(n_180), .Y(n_329) );
AND3x2_ASAP7_75t_L g388 ( .A(n_180), .B(n_389), .C(n_390), .Y(n_388) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_192), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_181), .B(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_181), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_181), .B(n_531), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_184), .A2(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_184), .A2(n_454), .B(n_455), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_184), .A2(n_514), .B(n_515), .Y(n_513) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_190), .C(n_191), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_188), .A2(n_191), .B(n_222), .C(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_191), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_191), .A2(n_517), .B(n_518), .Y(n_516) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_194), .Y(n_279) );
INVx1_ASAP7_75t_SL g323 ( .A(n_194), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_194), .B(n_272), .C(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_241), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_204), .A2(n_307), .B(n_359), .C(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_206), .B(n_228), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_206), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g375 ( .A(n_206), .Y(n_375) );
AND2x2_ASAP7_75t_L g396 ( .A(n_206), .B(n_243), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_206), .B(n_305), .Y(n_424) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AND2x2_ASAP7_75t_L g269 ( .A(n_207), .B(n_260), .Y(n_269) );
INVx2_ASAP7_75t_L g276 ( .A(n_207), .Y(n_276) );
AND2x2_ASAP7_75t_L g296 ( .A(n_207), .B(n_243), .Y(n_296) );
AND2x2_ASAP7_75t_L g346 ( .A(n_207), .B(n_228), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_207), .Y(n_350) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_215), .Y(n_528) );
INVx2_ASAP7_75t_SL g260 ( .A(n_217), .Y(n_260) );
BUFx2_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
AND2x2_ASAP7_75t_L g413 ( .A(n_217), .B(n_228), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g259 ( .A(n_227), .Y(n_259) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_227), .A2(n_523), .B(n_530), .Y(n_522) );
INVx3_ASAP7_75t_SL g243 ( .A(n_228), .Y(n_243) );
AND2x2_ASAP7_75t_L g268 ( .A(n_228), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g275 ( .A(n_228), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g305 ( .A(n_228), .B(n_265), .Y(n_305) );
OR2x2_ASAP7_75t_L g314 ( .A(n_228), .B(n_260), .Y(n_314) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_228), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_228), .B(n_290), .Y(n_337) );
AND2x2_ASAP7_75t_L g365 ( .A(n_228), .B(n_245), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_228), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g403 ( .A(n_228), .B(n_244), .Y(n_403) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_239), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .C(n_236), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_234), .A2(n_457), .B(n_458), .C(n_459), .Y(n_456) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_237), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g327 ( .A(n_243), .B(n_276), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_243), .B(n_269), .Y(n_355) );
AND2x2_ASAP7_75t_L g373 ( .A(n_243), .B(n_290), .Y(n_373) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_260), .Y(n_244) );
AND2x2_ASAP7_75t_L g274 ( .A(n_245), .B(n_260), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_245), .B(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g312 ( .A(n_245), .Y(n_312) );
OR2x2_ASAP7_75t_L g360 ( .A(n_245), .B(n_280), .Y(n_360) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_250), .B(n_258), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_247), .A2(n_266), .B(n_267), .Y(n_265) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_247), .A2(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AOI21xp5_ASAP7_75t_SL g504 ( .A1(n_248), .A2(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_249), .A2(n_453), .B(n_460), .Y(n_452) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_249), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_249), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_258), .Y(n_267) );
AND2x2_ASAP7_75t_L g295 ( .A(n_260), .B(n_265), .Y(n_295) );
INVx1_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
AND2x2_ASAP7_75t_L g398 ( .A(n_260), .B(n_276), .Y(n_398) );
AOI222xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_270), .B1(n_273), .B2(n_277), .C1(n_281), .C2(n_284), .Y(n_261) );
INVx1_ASAP7_75t_L g393 ( .A(n_262), .Y(n_393) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_268), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_263), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g300 ( .A(n_263), .B(n_269), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_263), .B(n_291), .Y(n_316) );
OAI222xp33_ASAP7_75t_L g338 ( .A1(n_263), .A2(n_339), .B1(n_344), .B2(n_345), .C1(n_353), .C2(n_355), .Y(n_338) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g326 ( .A(n_265), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_265), .B(n_346), .Y(n_386) );
AND2x2_ASAP7_75t_L g397 ( .A(n_265), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g405 ( .A(n_268), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_270), .B(n_321), .Y(n_384) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_272), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g342 ( .A(n_272), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx3_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_275), .A2(n_378), .B(n_381), .C(n_383), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_275), .B(n_312), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_275), .B(n_295), .Y(n_417) );
AND2x2_ASAP7_75t_L g290 ( .A(n_276), .B(n_286), .Y(n_290) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_280), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g369 ( .A(n_280), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g408 ( .A(n_280), .B(n_308), .Y(n_408) );
INVx1_ASAP7_75t_L g420 ( .A(n_280), .Y(n_420) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_283), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g401 ( .A(n_286), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_291), .B(n_293), .C(n_297), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_289), .A2(n_319), .B1(n_334), .B2(n_337), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_290), .B(n_304), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_290), .B(n_312), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_291), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g354 ( .A(n_291), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_291), .B(n_341), .Y(n_361) );
INVx2_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NOR4xp25_ASAP7_75t_L g299 ( .A(n_296), .B(n_300), .C(n_301), .D(n_304), .Y(n_299) );
INVx1_ASAP7_75t_SL g370 ( .A(n_297), .Y(n_370) );
AND2x2_ASAP7_75t_L g414 ( .A(n_297), .B(n_415), .Y(n_414) );
OAI211xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_306), .B(n_309), .C(n_318), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_305), .B(n_375), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_307), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_425) );
INVx1_ASAP7_75t_SL g380 ( .A(n_308), .Y(n_380) );
AND2x2_ASAP7_75t_L g419 ( .A(n_308), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_312), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_316), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_317), .B(n_342), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_324), .B(n_326), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g394 ( .A(n_321), .Y(n_394) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g422 ( .A(n_322), .Y(n_422) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B(n_333), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_329), .Y(n_341) );
OR2x2_ASAP7_75t_L g379 ( .A(n_329), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI21xp33_ASAP7_75t_SL g374 ( .A1(n_332), .A2(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_336), .A2(n_363), .B1(n_366), .B2(n_373), .C(n_374), .Y(n_362) );
INVx1_ASAP7_75t_SL g406 ( .A(n_337), .Y(n_406) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g353 ( .A(n_341), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_350), .B2(n_351), .Y(n_345) );
INVx1_ASAP7_75t_L g385 ( .A(n_346), .Y(n_385) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_349), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_391), .C(n_404), .D(n_416), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g357 ( .A(n_358), .B(n_362), .C(n_377), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_360), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_367), .B(n_372), .Y(n_376) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_379), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_409), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_381), .A2(n_396), .B(n_397), .C(n_399), .Y(n_395) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_382), .A2(n_400), .B1(n_402), .B2(n_403), .Y(n_399) );
INVx2_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_394), .C(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g410 ( .A(n_403), .Y(n_410) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_411), .B(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B1(n_421), .B2(n_423), .C(n_425), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_431), .A2(n_446), .B1(n_714), .B2(n_716), .Y(n_445) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g442 ( .A(n_436), .Y(n_442) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_437), .B(n_715), .Y(n_730) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g714 ( .A(n_438), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AOI21xp33_ASAP7_75t_SL g443 ( .A1(n_441), .A2(n_444), .B(n_731), .Y(n_443) );
INVx1_ASAP7_75t_L g724 ( .A(n_446), .Y(n_724) );
NAND2x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_630), .Y(n_446) );
NOR5xp2_ASAP7_75t_L g447 ( .A(n_448), .B(n_553), .C(n_585), .D(n_600), .E(n_617), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_481), .B(n_500), .C(n_541), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_462), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_450), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_450), .B(n_605), .Y(n_668) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_451), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_451), .B(n_497), .Y(n_554) );
AND2x2_ASAP7_75t_L g595 ( .A(n_451), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_451), .B(n_564), .Y(n_599) );
OR2x2_ASAP7_75t_L g636 ( .A(n_451), .B(n_487), .Y(n_636) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g486 ( .A(n_452), .B(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g544 ( .A(n_452), .Y(n_544) );
OR2x2_ASAP7_75t_L g707 ( .A(n_452), .B(n_547), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_462), .A2(n_610), .B1(n_611), .B2(n_614), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_462), .B(n_544), .Y(n_693) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_472), .Y(n_462) );
AND2x2_ASAP7_75t_L g499 ( .A(n_463), .B(n_487), .Y(n_499) );
AND2x2_ASAP7_75t_L g546 ( .A(n_463), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g551 ( .A(n_463), .Y(n_551) );
INVx3_ASAP7_75t_L g564 ( .A(n_463), .Y(n_564) );
OR2x2_ASAP7_75t_L g584 ( .A(n_463), .B(n_547), .Y(n_584) );
AND2x2_ASAP7_75t_L g603 ( .A(n_463), .B(n_473), .Y(n_603) );
BUFx2_ASAP7_75t_L g635 ( .A(n_463), .Y(n_635) );
AND2x4_ASAP7_75t_L g550 ( .A(n_472), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g485 ( .A(n_473), .Y(n_485) );
INVx2_ASAP7_75t_L g498 ( .A(n_473), .Y(n_498) );
OR2x2_ASAP7_75t_L g566 ( .A(n_473), .B(n_547), .Y(n_566) );
AND2x2_ASAP7_75t_L g596 ( .A(n_473), .B(n_487), .Y(n_596) );
AND2x2_ASAP7_75t_L g613 ( .A(n_473), .B(n_544), .Y(n_613) );
AND2x2_ASAP7_75t_L g653 ( .A(n_473), .B(n_564), .Y(n_653) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_473), .B(n_499), .Y(n_689) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_483), .B(n_496), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_484), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g627 ( .A1(n_485), .A2(n_499), .B(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_485), .B(n_487), .Y(n_683) );
AND2x2_ASAP7_75t_L g619 ( .A(n_486), .B(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_487), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_496), .B(n_544), .Y(n_712) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_497), .A2(n_655), .B1(n_656), .B2(n_661), .Y(n_654) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
AND2x2_ASAP7_75t_L g545 ( .A(n_498), .B(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g583 ( .A(n_498), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g620 ( .A(n_498), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_499), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g674 ( .A(n_499), .Y(n_674) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_521), .Y(n_501) );
INVx4_ASAP7_75t_L g560 ( .A(n_502), .Y(n_560) );
AND2x2_ASAP7_75t_L g638 ( .A(n_502), .B(n_605), .Y(n_638) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx3_ASAP7_75t_L g557 ( .A(n_503), .Y(n_557) );
AND2x2_ASAP7_75t_L g571 ( .A(n_503), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
INVx2_ASAP7_75t_L g589 ( .A(n_503), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_503), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g646 ( .A(n_503), .B(n_641), .Y(n_646) );
AND2x2_ASAP7_75t_L g711 ( .A(n_503), .B(n_681), .Y(n_711) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
AND2x2_ASAP7_75t_L g552 ( .A(n_512), .B(n_533), .Y(n_552) );
INVx2_ASAP7_75t_L g572 ( .A(n_512), .Y(n_572) );
INVx1_ASAP7_75t_L g577 ( .A(n_521), .Y(n_577) );
AND2x2_ASAP7_75t_L g623 ( .A(n_521), .B(n_571), .Y(n_623) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_532), .Y(n_521) );
INVx2_ASAP7_75t_L g562 ( .A(n_522), .Y(n_562) );
INVx1_ASAP7_75t_L g570 ( .A(n_522), .Y(n_570) );
AND2x2_ASAP7_75t_L g588 ( .A(n_522), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_522), .B(n_572), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .Y(n_525) );
AND2x2_ASAP7_75t_L g605 ( .A(n_532), .B(n_562), .Y(n_605) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g558 ( .A(n_533), .Y(n_558) );
AND2x2_ASAP7_75t_L g641 ( .A(n_533), .B(n_572), .Y(n_641) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_548), .B(n_552), .Y(n_541) );
INVx1_ASAP7_75t_SL g586 ( .A(n_542), .Y(n_586) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_543), .B(n_550), .Y(n_643) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g592 ( .A(n_544), .B(n_547), .Y(n_592) );
AND2x2_ASAP7_75t_L g621 ( .A(n_544), .B(n_565), .Y(n_621) );
OR2x2_ASAP7_75t_L g624 ( .A(n_544), .B(n_584), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_545), .A2(n_637), .B1(n_689), .B2(n_690), .C1(n_692), .C2(n_694), .Y(n_688) );
BUFx2_ASAP7_75t_L g602 ( .A(n_547), .Y(n_602) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g591 ( .A(n_550), .B(n_592), .Y(n_591) );
INVx3_ASAP7_75t_SL g608 ( .A(n_550), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_550), .B(n_602), .Y(n_662) );
AND2x2_ASAP7_75t_L g597 ( .A(n_552), .B(n_557), .Y(n_597) );
INVx1_ASAP7_75t_L g616 ( .A(n_552), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_555), .B1(n_559), .B2(n_563), .C(n_567), .Y(n_553) );
OR2x2_ASAP7_75t_L g625 ( .A(n_555), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g610 ( .A(n_557), .B(n_580), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_557), .B(n_570), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_557), .B(n_605), .Y(n_655) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_557), .Y(n_665) );
NAND2x1_ASAP7_75t_SL g676 ( .A(n_557), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g561 ( .A(n_558), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g581 ( .A(n_558), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_558), .B(n_576), .Y(n_607) );
INVx1_ASAP7_75t_L g673 ( .A(n_558), .Y(n_673) );
INVx1_ASAP7_75t_L g648 ( .A(n_559), .Y(n_648) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g660 ( .A(n_560), .Y(n_660) );
NOR2xp67_ASAP7_75t_L g672 ( .A(n_560), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g677 ( .A(n_561), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_561), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g580 ( .A(n_562), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_562), .B(n_572), .Y(n_593) );
INVx1_ASAP7_75t_L g659 ( .A(n_562), .Y(n_659) );
INVx1_ASAP7_75t_L g680 ( .A(n_563), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_573), .B(n_582), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g713 ( .A(n_569), .B(n_646), .Y(n_713) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g681 ( .A(n_570), .B(n_641), .Y(n_681) );
AOI32xp33_ASAP7_75t_L g594 ( .A1(n_571), .A2(n_577), .A3(n_595), .B1(n_597), .B2(n_598), .Y(n_594) );
AOI322xp5_ASAP7_75t_L g696 ( .A1(n_571), .A2(n_603), .A3(n_686), .B1(n_697), .B2(n_698), .C1(n_699), .C2(n_701), .Y(n_696) );
INVx2_ASAP7_75t_L g576 ( .A(n_572), .Y(n_576) );
INVx1_ASAP7_75t_L g686 ( .A(n_572), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_574), .B(n_580), .Y(n_629) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_575), .B(n_641), .Y(n_691) );
INVx1_ASAP7_75t_L g578 ( .A(n_576), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_576), .B(n_605), .Y(n_695) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_584), .B(n_679), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_587), .B1(n_590), .B2(n_593), .C(n_594), .Y(n_585) );
OR2x2_ASAP7_75t_L g606 ( .A(n_587), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g615 ( .A(n_587), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g640 ( .A(n_588), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g644 ( .A(n_598), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_604), .B1(n_606), .B2(n_608), .C(n_609), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_602), .A2(n_633), .B1(n_637), .B2(n_638), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_603), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_603), .Y(n_708) );
INVx1_ASAP7_75t_L g702 ( .A(n_605), .Y(n_702) );
INVx1_ASAP7_75t_SL g637 ( .A(n_606), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_608), .B(n_636), .Y(n_698) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_613), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g679 ( .A(n_613), .Y(n_679) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_622), .B1(n_624), .B2(n_625), .C(n_627), .Y(n_617) );
NOR2xp33_ASAP7_75t_SL g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_619), .A2(n_637), .B1(n_683), .B2(n_684), .Y(n_682) );
CKINVDCx14_ASAP7_75t_R g622 ( .A(n_623), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_624), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR3xp33_ASAP7_75t_SL g630 ( .A(n_631), .B(n_663), .C(n_687), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_639), .C(n_647), .D(n_654), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g710 ( .A(n_635), .Y(n_710) );
INVx3_ASAP7_75t_SL g704 ( .A(n_636), .Y(n_704) );
OR2x2_ASAP7_75t_L g709 ( .A(n_636), .B(n_710), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_644), .B2(n_646), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_641), .B(n_659), .Y(n_700) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B(n_651), .Y(n_647) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_666), .B(n_669), .C(n_682), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g697 ( .A(n_668), .Y(n_697) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_674), .B1(n_675), .B2(n_678), .C1(n_680), .C2(n_681), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND4xp25_ASAP7_75t_SL g706 ( .A(n_679), .B(n_707), .C(n_708), .D(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND3xp33_ASAP7_75t_SL g687 ( .A(n_688), .B(n_696), .C(n_705), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_705) );
INVx1_ASAP7_75t_L g726 ( .A(n_716), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_717), .Y(n_727) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
endmodule