module fake_jpeg_1676_n_553 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_553);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_49),
.Y(n_106)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_50),
.Y(n_164)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_51),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_53),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_14),
.C(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_15),
.B(n_14),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_32),
.B(n_14),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_72),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_15),
.B(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_83),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_35),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_27),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_76),
.B(n_82),
.Y(n_139)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_12),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_0),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_102),
.Y(n_125)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_25),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_40),
.Y(n_135)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_49),
.A2(n_51),
.B1(n_100),
.B2(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_115),
.B1(n_122),
.B2(n_143),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_45),
.B1(n_25),
.B2(n_30),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_114),
.A2(n_131),
.B1(n_44),
.B2(n_85),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_52),
.A2(n_45),
.B1(n_30),
.B2(n_37),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_55),
.A2(n_40),
.B1(n_37),
.B2(n_17),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_58),
.B(n_17),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_128),
.B(n_130),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_39),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_72),
.A2(n_21),
.B1(n_31),
.B2(n_39),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_31),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_50),
.A2(n_94),
.B1(n_84),
.B2(n_97),
.Y(n_143)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_24),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_150),
.B(n_166),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_73),
.A2(n_24),
.B1(n_23),
.B2(n_44),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_163),
.B1(n_81),
.B2(n_104),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_77),
.A2(n_23),
.B1(n_44),
.B2(n_18),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_78),
.B(n_21),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_122),
.A2(n_62),
.B1(n_59),
.B2(n_71),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_171),
.A2(n_196),
.B1(n_203),
.B2(n_209),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_109),
.A2(n_101),
.B1(n_57),
.B2(n_86),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_174),
.A2(n_194),
.B1(n_208),
.B2(n_165),
.Y(n_250)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_75),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_183),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_118),
.A2(n_106),
.B1(n_165),
.B2(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_179),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_184),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_66),
.B(n_98),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_206),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_113),
.A2(n_44),
.B1(n_91),
.B2(n_87),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_93),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_164),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_185),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_117),
.B(n_126),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_193),
.Y(n_237)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_192),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_80),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_195),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_74),
.B1(n_48),
.B2(n_18),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_105),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_106),
.B(n_2),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_202),
.B(n_146),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_144),
.A2(n_48),
.B1(n_18),
.B2(n_66),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_2),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_216),
.Y(n_239)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_121),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_144),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.Y(n_231)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_215),
.Y(n_233)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_110),
.B(n_5),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_139),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_164),
.B1(n_141),
.B2(n_145),
.Y(n_222)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_5),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_249),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_170),
.A2(n_143),
.B1(n_148),
.B2(n_155),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_223),
.A2(n_244),
.B(n_251),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_120),
.B1(n_151),
.B2(n_145),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_202),
.B1(n_206),
.B2(n_190),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_178),
.B(n_120),
.CI(n_163),
.CON(n_228),
.SN(n_228)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_228),
.B(n_159),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_SL g240 ( 
.A(n_172),
.B(n_121),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_156),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_180),
.A2(n_132),
.B1(n_160),
.B2(n_133),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_193),
.A2(n_148),
.B1(n_141),
.B2(n_133),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_181),
.A2(n_108),
.B1(n_161),
.B2(n_157),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_179),
.B(n_210),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_278),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_179),
.B(n_207),
.C(n_183),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_258),
.A2(n_260),
.B(n_252),
.Y(n_304)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

AO22x1_ASAP7_75t_SL g260 ( 
.A1(n_223),
.A2(n_202),
.B1(n_218),
.B2(n_205),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_275),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_220),
.A2(n_184),
.B(n_191),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_263),
.B(n_274),
.Y(n_294)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_175),
.C(n_204),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_269),
.C(n_273),
.Y(n_289)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_220),
.B(n_216),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_268),
.B(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_214),
.C(n_187),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_282),
.B1(n_235),
.B2(n_247),
.Y(n_288)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_237),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_221),
.A2(n_228),
.B(n_250),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_227),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_167),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_277),
.B(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_249),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_221),
.A2(n_119),
.B(n_215),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_286),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_239),
.B(n_213),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_284),
.A2(n_224),
.B1(n_249),
.B2(n_240),
.Y(n_310)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_285),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_168),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_288),
.A2(n_292),
.B1(n_295),
.B2(n_302),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_242),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_293),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_221),
.B1(n_244),
.B2(n_235),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_280),
.A2(n_235),
.B1(n_249),
.B2(n_252),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_280),
.B1(n_266),
.B2(n_257),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_235),
.B1(n_238),
.B2(n_252),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_308),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_309),
.B(n_310),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_285),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_231),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_311),
.B(n_315),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_286),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_232),
.Y(n_316)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_271),
.A2(n_251),
.B1(n_222),
.B2(n_232),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_248),
.B1(n_254),
.B2(n_226),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_280),
.A2(n_189),
.B1(n_160),
.B2(n_197),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_318),
.A2(n_234),
.B1(n_236),
.B2(n_254),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_273),
.B(n_256),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_319),
.B(n_291),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_258),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_320),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_267),
.C(n_269),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_337),
.C(n_294),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_336),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_295),
.A2(n_277),
.B(n_274),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_324),
.A2(n_325),
.B(n_335),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_297),
.A2(n_284),
.B(n_263),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_302),
.A2(n_280),
.B1(n_266),
.B2(n_260),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_334),
.B1(n_339),
.B2(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

AO22x1_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_266),
.B1(n_278),
.B2(n_265),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_338),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_309),
.A2(n_260),
.B1(n_268),
.B2(n_281),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_279),
.B(n_259),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_264),
.C(n_255),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

OAI22x1_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_276),
.B1(n_272),
.B2(n_261),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_347),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_343),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_310),
.A2(n_224),
.B(n_255),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_348),
.B(n_354),
.Y(n_360)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_297),
.A2(n_201),
.B(n_247),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_307),
.B1(n_243),
.B2(n_246),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_256),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_290),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_317),
.A2(n_236),
.B1(n_243),
.B2(n_234),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_353),
.A2(n_318),
.B1(n_292),
.B2(n_315),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_293),
.A2(n_173),
.B(n_219),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_352),
.Y(n_357)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_344),
.A2(n_303),
.B1(n_304),
.B2(n_299),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_359),
.A2(n_236),
.B1(n_230),
.B2(n_226),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_345),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_361),
.B(n_230),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_325),
.B(n_294),
.CI(n_301),
.CON(n_362),
.SN(n_362)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_376),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_345),
.Y(n_363)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_363),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_365),
.C(n_372),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_319),
.C(n_313),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_324),
.A2(n_304),
.B(n_299),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_366),
.A2(n_360),
.B(n_326),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_377),
.B1(n_382),
.B2(n_385),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_313),
.C(n_291),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_350),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_308),
.Y(n_374)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_301),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_375),
.B(n_331),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_344),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_328),
.A2(n_300),
.B1(n_312),
.B2(n_314),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_300),
.Y(n_380)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_314),
.B1(n_307),
.B2(n_298),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_119),
.C(n_153),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_323),
.C(n_321),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_334),
.Y(n_384)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

NOR3xp33_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_346),
.C(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_393),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_357),
.A2(n_327),
.B1(n_349),
.B2(n_347),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

AOI21xp33_ASAP7_75t_L g423 ( 
.A1(n_395),
.A2(n_418),
.B(n_378),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_348),
.Y(n_396)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_396),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_387),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_408),
.Y(n_439)
);

BUFx5_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

BUFx12_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_404),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_364),
.B(n_372),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_410),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_409),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_369),
.A2(n_354),
.B1(n_335),
.B2(n_341),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_321),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_340),
.C(n_339),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_413),
.C(n_415),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_355),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_342),
.C(n_332),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_332),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_371),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_353),
.C(n_188),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_417),
.A2(n_370),
.B1(n_379),
.B2(n_358),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_402),
.A2(n_359),
.B1(n_369),
.B2(n_366),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_422),
.A2(n_431),
.B1(n_435),
.B2(n_417),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_424),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_377),
.C(n_380),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_382),
.C(n_356),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_427),
.C(n_432),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_379),
.C(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_430),
.B(n_153),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_385),
.B1(n_368),
.B2(n_387),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_368),
.C(n_386),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_414),
.C(n_411),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_444),
.C(n_391),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_386),
.B1(n_358),
.B2(n_355),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_246),
.Y(n_437)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_392),
.A2(n_362),
.B1(n_185),
.B2(n_192),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_440),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_395),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_397),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_415),
.C(n_389),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_416),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_453),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_442),
.A2(n_403),
.B(n_392),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_447),
.A2(n_454),
.B(n_459),
.Y(n_477)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_388),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_451),
.B(n_466),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_422),
.A2(n_403),
.B(n_398),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_420),
.A2(n_391),
.B1(n_362),
.B2(n_397),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_456),
.A2(n_219),
.B1(n_245),
.B2(n_211),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_430),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_404),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_462),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_434),
.A2(n_404),
.B(n_407),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_407),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_461),
.B1(n_447),
.B2(n_443),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_412),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_412),
.C(n_212),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_426),
.C(n_432),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_412),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_245),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_444),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_465),
.A2(n_438),
.B1(n_429),
.B2(n_439),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_195),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_428),
.C(n_431),
.Y(n_483)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_471),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_480),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_425),
.C(n_426),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_473),
.B(n_485),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_476),
.A2(n_454),
.B(n_457),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_440),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_245),
.B(n_112),
.Y(n_499)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_481),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_439),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_483),
.B(n_137),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_435),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_487),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_173),
.C(n_186),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_448),
.A2(n_157),
.B1(n_200),
.B2(n_199),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_488),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_219),
.B1(n_245),
.B2(n_112),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_137),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_452),
.C(n_449),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_490),
.B(n_497),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_491),
.A2(n_492),
.B(n_5),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_469),
.A2(n_452),
.B(n_463),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_478),
.A2(n_450),
.B1(n_468),
.B2(n_467),
.Y(n_497)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_499),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g501 ( 
.A(n_483),
.B(n_112),
.CI(n_199),
.CON(n_501),
.SN(n_501)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_503),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_504),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_200),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_484),
.Y(n_505)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_505),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_473),
.B(n_5),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_506),
.B(n_6),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_471),
.C(n_477),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_508),
.A2(n_500),
.B(n_499),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_495),
.A2(n_474),
.B1(n_480),
.B2(n_472),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_511),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_482),
.C(n_489),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_485),
.C(n_6),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_516),
.Y(n_528)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_514),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_494),
.A2(n_6),
.B(n_7),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_515),
.A2(n_514),
.B(n_522),
.Y(n_531)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_521),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_7),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_520),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_496),
.B(n_7),
.C(n_8),
.Y(n_521)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_500),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_530),
.B(n_532),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_533),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_519),
.A2(n_501),
.B(n_498),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_502),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_513),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_535),
.B(n_540),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_528),
.A2(n_517),
.B(n_509),
.Y(n_539)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_539),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_521),
.Y(n_540)
);

NOR2x1_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_525),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_541),
.A2(n_538),
.B(n_504),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_525),
.C(n_520),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g546 ( 
.A1(n_542),
.A2(n_543),
.B(n_539),
.Y(n_546)
);

A2O1A1Ixp33_ASAP7_75t_SL g543 ( 
.A1(n_534),
.A2(n_529),
.B(n_501),
.C(n_517),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_546),
.A2(n_547),
.B(n_548),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_545),
.A2(n_7),
.B(n_8),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_544),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_8),
.C(n_9),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_8),
.C(n_9),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_10),
.Y(n_553)
);


endmodule