module fake_jpeg_29146_n_180 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_0),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_1),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_26),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_2),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_59),
.B(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_65),
.B1(n_70),
.B2(n_72),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_92),
.B(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_70),
.B1(n_65),
.B2(n_72),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_89),
.B1(n_91),
.B2(n_69),
.Y(n_102)
);

OR2x2_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_54),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_66),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_67),
.B1(n_52),
.B2(n_56),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_67),
.B1(n_52),
.B2(n_56),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_54),
.B1(n_51),
.B2(n_57),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_95),
.B(n_59),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_38),
.B(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_105),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_93),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_34),
.B1(n_48),
.B2(n_47),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_111),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_108),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_51),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_114),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_112),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_61),
.B1(n_68),
.B2(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_110),
.B1(n_9),
.B2(n_11),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_53),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_3),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_22),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_126),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_29),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_24),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_129),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_33),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_15),
.C(n_19),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_8),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_131),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_121),
.B(n_129),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_49),
.B1(n_27),
.B2(n_32),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_12),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_40),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_36),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_146),
.B(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_37),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_42),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_135),
.C(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_43),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_45),
.C(n_46),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_125),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_127),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_127),
.B(n_135),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_147),
.B(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_147),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_169),
.B(n_170),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_149),
.B(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_160),
.B1(n_159),
.B2(n_163),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_162),
.C(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_157),
.Y(n_180)
);


endmodule