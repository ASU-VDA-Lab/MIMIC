module fake_jpeg_24809_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_36),
.B1(n_34),
.B2(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_18),
.Y(n_99)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_65),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_49),
.B1(n_48),
.B2(n_41),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_37),
.B1(n_39),
.B2(n_28),
.Y(n_104)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_69),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_31),
.B1(n_35),
.B2(n_17),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_70),
.B1(n_37),
.B2(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_31),
.B1(n_35),
.B2(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_18),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_41),
.B1(n_48),
.B2(n_17),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_72),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_43),
.B1(n_32),
.B2(n_37),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_80),
.B1(n_99),
.B2(n_28),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_45),
.CI(n_23),
.CON(n_76),
.SN(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_40),
.B1(n_44),
.B2(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_85),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_101),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_25),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_88),
.B(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_25),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_38),
.B(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_39),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_47),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_36),
.B1(n_34),
.B2(n_25),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_50),
.B1(n_46),
.B2(n_26),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_74),
.B1(n_91),
.B2(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_120),
.B1(n_121),
.B2(n_135),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_50),
.B1(n_46),
.B2(n_26),
.Y(n_120)
);

AO22x1_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_22),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_82),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_24),
.B1(n_19),
.B2(n_33),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_50),
.B1(n_46),
.B2(n_33),
.Y(n_130)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_151),
.Y(n_186)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_150),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_76),
.B(n_88),
.C(n_84),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_155),
.B(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_81),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_153),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_84),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_163),
.B(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_117),
.B(n_76),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_165),
.B(n_123),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_80),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_123),
.C(n_122),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_103),
.B(n_102),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_88),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_169),
.B(n_143),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_130),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_138),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_113),
.B(n_134),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_172),
.A2(n_196),
.B(n_180),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_176),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_183),
.C(n_185),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_121),
.B(n_131),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_187),
.B(n_138),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_121),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_184),
.B(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_98),
.C(n_101),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_121),
.B(n_79),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_92),
.B1(n_87),
.B2(n_116),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_144),
.B1(n_158),
.B2(n_139),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_116),
.B1(n_114),
.B2(n_118),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_197),
.B1(n_201),
.B2(n_191),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_159),
.C(n_137),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_199),
.C(n_29),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_198),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_133),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_114),
.B1(n_118),
.B2(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_132),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_14),
.C(n_2),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_12),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_125),
.B1(n_126),
.B2(n_24),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_204),
.B1(n_201),
.B2(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_171),
.A2(n_149),
.B1(n_137),
.B2(n_157),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_165),
.B1(n_144),
.B2(n_125),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_224),
.B1(n_178),
.B2(n_184),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_21),
.B(n_2),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_214),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_222),
.C(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_139),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_218),
.A2(n_221),
.B(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_139),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_106),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_143),
.B1(n_29),
.B2(n_27),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_1),
.B(n_2),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_225),
.A2(n_227),
.B(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_27),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_21),
.B(n_1),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_232),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_170),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_251),
.C(n_231),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_250),
.B1(n_252),
.B2(n_257),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_199),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_189),
.B1(n_181),
.B2(n_183),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_185),
.C(n_189),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_187),
.B1(n_172),
.B2(n_174),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_217),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_1),
.B(n_4),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_230),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_229),
.B1(n_228),
.B2(n_218),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_215),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_268),
.C(n_275),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_214),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_232),
.C(n_210),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_213),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_207),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_205),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_216),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_219),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_218),
.C(n_206),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_276),
.B(n_279),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_211),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_252),
.C(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_257),
.B(n_248),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_244),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_233),
.B1(n_239),
.B2(n_247),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_284),
.B1(n_202),
.B2(n_248),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_237),
.B1(n_204),
.B2(n_243),
.Y(n_284)
);

BUFx12_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_7),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_273),
.B(n_264),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_290),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_237),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_241),
.B(n_266),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_255),
.C(n_234),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_100),
.C(n_1),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_300),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_295),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_305),
.B(n_309),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_271),
.B1(n_258),
.B2(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_313),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_310),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_311),
.B(n_8),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_287),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_307),
.B(n_308),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_5),
.B(n_6),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_6),
.C(n_7),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_293),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_7),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_8),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_286),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_316),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_318),
.B(n_302),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_294),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_323),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_324),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_306),
.B(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_322),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_303),
.B(n_285),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_332),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_288),
.B(n_285),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_330),
.A2(n_334),
.B(n_317),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_288),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_320),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_9),
.C(n_10),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_337),
.B(n_338),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_315),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_340),
.C(n_329),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_12),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_12),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_341),
.A2(n_329),
.B(n_15),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_343),
.C(n_338),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_345),
.Y(n_346)
);

AOI321xp33_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_344),
.A3(n_335),
.B1(n_336),
.B2(n_15),
.C(n_16),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_13),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_13),
.Y(n_349)
);


endmodule