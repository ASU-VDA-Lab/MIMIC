module fake_jpeg_31965_n_418 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_418);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_418;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_11),
.B(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_74),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_14),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_14),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_14),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_13),
.Y(n_84)
);

OR2x4_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_40),
.B1(n_25),
.B2(n_28),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_89),
.A2(n_36),
.B1(n_19),
.B2(n_43),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_17),
.Y(n_156)
);

CKINVDCx6p67_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_103),
.Y(n_159)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_28),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_51),
.Y(n_142)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_54),
.B1(n_86),
.B2(n_80),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_162),
.B1(n_167),
.B2(n_43),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_36),
.B(n_19),
.C(n_43),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_141),
.A2(n_165),
.B(n_175),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_156),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_28),
.B1(n_88),
.B2(n_53),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_151),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_60),
.C(n_75),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_46),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_169),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_105),
.A2(n_61),
.B1(n_67),
.B2(n_64),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_101),
.B(n_33),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_59),
.B1(n_56),
.B2(n_79),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_176),
.B1(n_114),
.B2(n_127),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_23),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_177),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_92),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_63),
.B1(n_50),
.B2(n_33),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_89),
.B1(n_127),
.B2(n_110),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_186),
.A2(n_188),
.B1(n_198),
.B2(n_152),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_130),
.B(n_103),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_190),
.A2(n_20),
.B(n_38),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_101),
.B(n_120),
.C(n_39),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_159),
.B(n_165),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_176),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_17),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_110),
.B1(n_119),
.B2(n_99),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_112),
.B1(n_119),
.B2(n_111),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_137),
.A2(n_112),
.B1(n_118),
.B2(n_95),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_141),
.A2(n_94),
.B1(n_113),
.B2(n_45),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_94),
.B1(n_45),
.B2(n_42),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_153),
.A2(n_126),
.B1(n_24),
.B2(n_19),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_159),
.B1(n_160),
.B2(n_166),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_140),
.B(n_44),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_0),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_143),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_228),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_147),
.C(n_139),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_220),
.C(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_143),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_231),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_216),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_174),
.B1(n_145),
.B2(n_150),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_229),
.B1(n_240),
.B2(n_242),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_148),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_163),
.B1(n_159),
.B2(n_168),
.Y(n_229)
);

AO22x1_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_200),
.B1(n_186),
.B2(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_170),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_169),
.C(n_177),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_244),
.B1(n_210),
.B2(n_212),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_16),
.CI(n_44),
.CON(n_234),
.SN(n_234)
);

OAI21xp33_ASAP7_75t_L g277 ( 
.A1(n_234),
.A2(n_238),
.B(n_243),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_235),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_39),
.B(n_38),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_239),
.B(n_194),
.Y(n_259)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_237),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_23),
.B(n_22),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_178),
.B1(n_24),
.B2(n_22),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_193),
.B(n_13),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_188),
.A2(n_183),
.B1(n_198),
.B2(n_192),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_16),
.B1(n_20),
.B2(n_3),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_242),
.B1(n_224),
.B2(n_225),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_20),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_247),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_248),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_182),
.B(n_20),
.C(n_2),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_235),
.A2(n_212),
.B1(n_215),
.B2(n_189),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_256),
.A2(n_245),
.B(n_208),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_257),
.A2(n_272),
.B1(n_253),
.B2(n_244),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_261),
.B1(n_227),
.B2(n_229),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_259),
.B(n_243),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_212),
.B1(n_181),
.B2(n_187),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_217),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_225),
.A2(n_213),
.B1(n_181),
.B2(n_187),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_215),
.B1(n_209),
.B2(n_189),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_276),
.B(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_208),
.B(n_184),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_280),
.A2(n_254),
.B(n_277),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_281),
.A2(n_271),
.B1(n_279),
.B2(n_275),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_218),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_284),
.C(n_306),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_255),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_299),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_220),
.C(n_232),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_228),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_274),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_290),
.B1(n_292),
.B2(n_302),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_250),
.B(n_234),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_289),
.B(n_259),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_230),
.B1(n_221),
.B2(n_226),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_297),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_230),
.B1(n_241),
.B2(n_240),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_293),
.A2(n_294),
.B(n_303),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_263),
.B(n_268),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_234),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_276),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_300),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_257),
.A2(n_230),
.B1(n_238),
.B2(n_235),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_254),
.A2(n_249),
.B(n_184),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_272),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_253),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_191),
.C(n_185),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_310),
.B(n_320),
.Y(n_347)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_313),
.B(n_314),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_279),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_316),
.B(n_330),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_268),
.B(n_269),
.C(n_265),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_318),
.A2(n_297),
.B(n_280),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_258),
.B1(n_261),
.B2(n_271),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_206),
.B1(n_20),
.B2(n_5),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_295),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_321),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_329),
.B1(n_292),
.B2(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

NAND2x1p5_ASAP7_75t_R g326 ( 
.A(n_300),
.B(n_260),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_303),
.B(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_327),
.A2(n_301),
.B1(n_283),
.B2(n_286),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_281),
.A2(n_262),
.B1(n_270),
.B2(n_267),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_267),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_331),
.A2(n_333),
.B1(n_342),
.B2(n_348),
.Y(n_358)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_322),
.A2(n_287),
.B1(n_294),
.B2(n_293),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_284),
.C(n_282),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_335),
.B(n_337),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_285),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_338),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_306),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_323),
.A2(n_301),
.B1(n_286),
.B2(n_262),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_191),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_349),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_203),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_349),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_323),
.A2(n_278),
.B1(n_185),
.B2(n_202),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_278),
.Y(n_349)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

AOI22x1_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_312),
.B1(n_326),
.B2(n_308),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_315),
.B1(n_329),
.B2(n_346),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_318),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_362),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_355),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_307),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_361),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_347),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_317),
.B1(n_308),
.B2(n_319),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_363),
.A2(n_365),
.B(n_331),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_317),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_339),
.C(n_348),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_314),
.Y(n_365)
);

AOI211xp5_ASAP7_75t_SL g366 ( 
.A1(n_345),
.A2(n_315),
.B(n_321),
.C(n_330),
.Y(n_366)
);

AOI211xp5_ASAP7_75t_L g375 ( 
.A1(n_366),
.A2(n_336),
.B(n_327),
.C(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_3),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_356),
.A2(n_336),
.B(n_341),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_369),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_372),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_371),
.A2(n_367),
.B1(n_357),
.B2(n_352),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_342),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_379),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_375),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_389)
);

OA21x2_ASAP7_75t_L g377 ( 
.A1(n_353),
.A2(n_309),
.B(n_325),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_8),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_325),
.C(n_309),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_351),
.C(n_352),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_206),
.Y(n_379)
);

AOI21xp33_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_358),
.B(n_359),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_380),
.B(n_351),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_384),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_382),
.B(n_377),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g385 ( 
.A(n_371),
.B(n_0),
.CI(n_3),
.CON(n_385),
.SN(n_385)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_386),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_389),
.A2(n_9),
.B(n_10),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_372),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_391),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_8),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_8),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_388),
.B(n_376),
.Y(n_394)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_394),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_397),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_385),
.A2(n_374),
.B1(n_378),
.B2(n_379),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_SL g402 ( 
.A(n_399),
.B(n_401),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_396),
.A2(n_393),
.B(n_400),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_403),
.A2(n_405),
.B(n_407),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_400),
.A2(n_399),
.B(n_390),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_398),
.A2(n_381),
.B(n_387),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_404),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_409),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_387),
.Y(n_409)
);

AO21x2_ASAP7_75t_L g410 ( 
.A1(n_402),
.A2(n_389),
.B(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_410),
.B(n_373),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_413),
.B(n_411),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_412),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_415),
.A2(n_381),
.B(n_370),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_9),
.C(n_10),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_417),
.B(n_9),
.Y(n_418)
);


endmodule