module real_jpeg_13259_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_320, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_320;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_62),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_62),
.B1(n_67),
.B2(n_72),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_4),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_165),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_4),
.A2(n_67),
.B1(n_72),
.B2(n_165),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_120),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_120),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_6),
.A2(n_67),
.B1(n_72),
.B2(n_120),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_186),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_7),
.A2(n_24),
.B1(n_26),
.B2(n_186),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_7),
.A2(n_67),
.B1(n_72),
.B2(n_186),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_11),
.A2(n_24),
.B1(n_26),
.B2(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_11),
.A2(n_47),
.B1(n_67),
.B2(n_72),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_51),
.B1(n_67),
.B2(n_72),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_51),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_13),
.A2(n_38),
.B(n_39),
.C(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_13),
.B(n_49),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_13),
.A2(n_24),
.B1(n_26),
.B2(n_179),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_13),
.A2(n_136),
.B1(n_137),
.B2(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_13),
.B(n_31),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_14),
.A2(n_24),
.B1(n_26),
.B2(n_33),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_33),
.B1(n_67),
.B2(n_72),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_14),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_122)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_93),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_77),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_77),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_19),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_34),
.CI(n_52),
.CON(n_19),
.SN(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_31),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_21),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_21),
.A2(n_31),
.B1(n_87),
.B2(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_21),
.A2(n_32),
.B(n_90),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_21),
.A2(n_31),
.B1(n_182),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_21),
.A2(n_31),
.B1(n_215),
.B2(n_228),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_58),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_22),
.A2(n_56),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_22),
.A2(n_88),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OA22x2_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_23),
.A2(n_26),
.B(n_227),
.C(n_229),
.Y(n_226)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_24),
.A2(n_26),
.B1(n_70),
.B2(n_73),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g229 ( 
.A(n_24),
.B(n_27),
.C(n_29),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_26),
.B(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_38),
.B2(n_43),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_29),
.A2(n_43),
.B(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g228 ( 
.A(n_30),
.B(n_179),
.CON(n_228),
.SN(n_228)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_32),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_45),
.B(n_48),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_35),
.A2(n_118),
.B(n_121),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_35),
.A2(n_48),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_35),
.A2(n_44),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_46),
.B1(n_49),
.B2(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_36),
.B(n_50),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_36),
.A2(n_49),
.B1(n_119),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_36),
.A2(n_49),
.B1(n_185),
.B2(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_37)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_61),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_49),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.C(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_55),
.A2(n_88),
.B(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_63),
.A2(n_64),
.B1(n_84),
.B2(n_85),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_81),
.C(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_74),
.B(n_76),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_74),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_76),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_65),
.A2(n_74),
.B1(n_234),
.B2(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_65),
.A2(n_74),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_65),
.A2(n_74),
.B1(n_242),
.B2(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_66),
.B(n_131),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_66),
.A2(n_113),
.B(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_66),
.B(n_179),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_SL g73 ( 
.A(n_70),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_70),
.B(n_72),
.C(n_179),
.Y(n_249)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_72),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_74),
.A2(n_114),
.B(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_74),
.A2(n_76),
.B(n_141),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_83),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_81),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_81),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_83),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B(n_89),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_301),
.B(n_314),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_166),
.B(n_300),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_148),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_96),
.B(n_148),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_123),
.B2(n_147),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_97),
.B(n_124),
.C(n_133),
.Y(n_312)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_115),
.C(n_117),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_99),
.A2(n_100),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_101),
.A2(n_102),
.B1(n_110),
.B2(n_111),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_103),
.A2(n_136),
.B(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_104),
.A2(n_109),
.B1(n_158),
.B2(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_104),
.A2(n_109),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_105),
.A2(n_109),
.B(n_160),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_106),
.A2(n_137),
.B(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_117),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_133),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B(n_132),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_127),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_128),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_132),
.B(n_304),
.C(n_308),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_132),
.B(n_304),
.CI(n_308),
.CON(n_313),
.SN(n_313)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_142),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_134),
.A2(n_135),
.B(n_144),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_157),
.B(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_136),
.A2(n_137),
.B1(n_257),
.B2(n_265),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_137),
.B(n_179),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_153),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_154),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.C(n_163),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_161),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_294),
.B(n_299),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_203),
.B1(n_219),
.B2(n_293),
.C(n_320),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_192),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_169),
.B(n_192),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_188),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_170),
.B(n_189),
.C(n_190),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_180),
.C(n_183),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_172),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_202),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_217),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_204),
.B(n_217),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_209),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_205),
.B(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_207),
.B(n_209),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_292),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_287),
.B(n_291),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_243),
.B(n_286),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_238),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_238),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_225),
.B(n_231),
.C(n_235),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_230),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_241),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_281),
.B(n_285),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_271),
.B(n_280),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_260),
.B(n_270),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_255),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_253),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_266),
.B(n_269),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_276),
.C(n_279),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_311),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_313),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_313),
.Y(n_319)
);


endmodule