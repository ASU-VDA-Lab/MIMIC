module real_jpeg_17537_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_2),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_65),
.B1(n_154),
.B2(n_160),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_2),
.A2(n_65),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_2),
.A2(n_65),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_576),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_3),
.B(n_577),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_4),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_5),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_5),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_6),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_7),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_7),
.A2(n_236),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_7),
.A2(n_236),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_7),
.A2(n_236),
.B1(n_504),
.B2(n_509),
.Y(n_503)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_8),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_8),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_8),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_9),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_9),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_9),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_9),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_10),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_114),
.B1(n_138),
.B2(n_142),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_10),
.A2(n_114),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_10),
.A2(n_114),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_11),
.A2(n_27),
.B1(n_278),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_11),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_11),
.A2(n_308),
.B1(n_357),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_11),
.A2(n_308),
.B1(n_437),
.B2(n_442),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_11),
.A2(n_308),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_13),
.A2(n_273),
.A3(n_277),
.B1(n_279),
.B2(n_284),
.Y(n_272)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_13),
.A2(n_67),
.B1(n_283),
.B2(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_13),
.B(n_45),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_13),
.B(n_98),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_13),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_13),
.B(n_118),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_13),
.A2(n_156),
.B1(n_283),
.B2(n_512),
.Y(n_511)
);

OAI32xp33_ASAP7_75t_L g515 ( 
.A1(n_13),
.A2(n_516),
.A3(n_518),
.B1(n_519),
.B2(n_523),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_32),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_14),
.A2(n_35),
.B1(n_216),
.B2(n_220),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_14),
.A2(n_35),
.B1(n_291),
.B2(n_297),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_14),
.A2(n_35),
.B1(n_325),
.B2(n_329),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_15),
.Y(n_190)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_15),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_16),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_16),
.A2(n_33),
.B1(n_78),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_16),
.A2(n_78),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_16),
.A2(n_78),
.B1(n_218),
.B2(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g335 ( 
.A(n_17),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_175),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_173),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_22),
.B(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_146),
.C(n_151),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_24),
.A2(n_146),
.B1(n_557),
.B2(n_558),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_24),
.Y(n_557)
);

XNOR2x1_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_69),
.Y(n_24)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_25),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g146 ( 
.A1(n_26),
.A2(n_58),
.B(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_29),
.Y(n_286)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_30),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_33),
.Y(n_149)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_36),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_36),
.A2(n_59),
.B(n_168),
.Y(n_167)
);

OAI22x1_ASAP7_75t_SL g227 ( 
.A1(n_36),
.A2(n_58),
.B1(n_228),
.B2(n_235),
.Y(n_227)
);

OAI21x1_ASAP7_75t_SL g330 ( 
.A1(n_36),
.A2(n_235),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_36),
.A2(n_58),
.B1(n_307),
.B2(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_36),
.A2(n_168),
.B(n_400),
.Y(n_399)
);

OR2x6_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_41),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_41),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_41),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_43),
.Y(n_230)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_45),
.B(n_148),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_45),
.A2(n_150),
.B1(n_306),
.B2(n_309),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_45),
.B(n_332),
.Y(n_331)
);

AO22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_55),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_50),
.Y(n_159)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_50),
.Y(n_370)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_53),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_54),
.Y(n_163)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_54),
.Y(n_270)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_117),
.B2(n_145),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_145),
.C(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_82),
.B(n_109),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_72),
.B(n_98),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_72),
.Y(n_323)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_77),
.Y(n_328)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

AOI21x1_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_153),
.B(n_164),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_82),
.A2(n_98),
.B(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_82),
.A2(n_109),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_82),
.A2(n_98),
.B1(n_153),
.B2(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_83),
.A2(n_111),
.B(n_165),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_83),
.A2(n_110),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_83),
.A2(n_110),
.B1(n_264),
.B2(n_353),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_L g366 ( 
.A1(n_83),
.A2(n_110),
.B1(n_353),
.B2(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_83),
.A2(n_110),
.B1(n_367),
.B2(n_511),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_98),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B1(n_92),
.B2(n_95),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_90),
.Y(n_265)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_105),
.Y(n_98)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_100),
.Y(n_435)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_101),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_102),
.Y(n_456)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_103),
.Y(n_255)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_107),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_113),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_146),
.C(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_117),
.B(n_152),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_127),
.B(n_136),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_118),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_118),
.B(n_223),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_118),
.A2(n_127),
.B1(n_434),
.B2(n_436),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_118),
.A2(n_127),
.B1(n_436),
.B2(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_119),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_119),
.B(n_137),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_119),
.A2(n_252),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_119)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_120),
.Y(n_448)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_120),
.Y(n_486)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_121),
.Y(n_423)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_124),
.Y(n_248)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_124),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_127),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_127),
.A2(n_394),
.B(n_539),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_131),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_135),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_137),
.A2(n_252),
.B(n_318),
.Y(n_347)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_146),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_146),
.A2(n_558),
.B1(n_561),
.B2(n_562),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_151),
.B(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_159),
.Y(n_329)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_160),
.Y(n_357)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_163),
.Y(n_517)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g578 ( 
.A(n_166),
.Y(n_578)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.CI(n_171),
.CON(n_166),
.SN(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_553),
.B(n_573),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_405),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_340),
.B(n_381),
.C(n_382),
.D(n_404),
.Y(n_178)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_179),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_310),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_180),
.B(n_310),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_239),
.C(n_260),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_181),
.A2(n_182),
.B1(n_239),
.B2(n_240),
.Y(n_342)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_226),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_183),
.B(n_227),
.C(n_238),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_213),
.Y(n_183)
);

XOR2x2_ASAP7_75t_L g358 ( 
.A(n_184),
.B(n_213),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_193),
.B(n_200),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_185),
.A2(n_193),
.B1(n_290),
.B2(n_301),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_185),
.A2(n_464),
.B1(n_469),
.B2(n_470),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_185),
.A2(n_200),
.B(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_186),
.B(n_206),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_186),
.A2(n_246),
.B(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_186),
.A2(n_446),
.B(n_452),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_186),
.A2(n_283),
.B1(n_477),
.B2(n_478),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_186),
.A2(n_465),
.B1(n_478),
.B2(n_492),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_188),
.Y(n_480)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_189),
.Y(n_451)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_190),
.Y(n_421)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_205),
.Y(n_489)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_222),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_225),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_228),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_234),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_230),
.Y(n_351)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_231),
.A2(n_234),
.B1(n_354),
.B2(n_357),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_231),
.A2(n_234),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_231),
.A2(n_234),
.B1(n_430),
.B2(n_466),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_250),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_241),
.B(n_250),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_242),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_246),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_249),
.A2(n_290),
.B(n_375),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_252),
.A2(n_253),
.B(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_259),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_260),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_271),
.C(n_305),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_262),
.B(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_268),
.Y(n_513)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_271),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_289),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_272),
.B(n_289),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_283),
.B(n_425),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_283),
.A2(n_424),
.B(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_283),
.B(n_520),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_304),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_320),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_320),
.C(n_337),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g397 ( 
.A(n_313),
.B(n_317),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_313),
.A2(n_319),
.B1(n_399),
.B2(n_401),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g565 ( 
.A1(n_319),
.A2(n_401),
.B(n_566),
.Y(n_565)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_336),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_330),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_336),
.C(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.C(n_359),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_341),
.B(n_343),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.C(n_358),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_358),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.C(n_352),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_352),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx2_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_379),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_360),
.B(n_379),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.C(n_365),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_361),
.B(n_550),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_365),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.C(n_373),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_366),
.B(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_371),
.A2(n_372),
.B1(n_374),
.B2(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_374),
.Y(n_543)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_375),
.Y(n_492)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_407),
.C(n_410),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_385),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_386),
.B(n_396),
.C(n_402),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_396),
.B1(n_402),
.B2(n_403),
.Y(n_388)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_389),
.Y(n_402)
);

OAI21xp33_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_392),
.B(n_395),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_392),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_395),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_395),
.A2(n_560),
.B1(n_563),
.B2(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_396),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_397),
.Y(n_566)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_546),
.B(n_552),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_533),
.B(n_545),
.Y(n_412)
);

OAI21x1_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_497),
.B(n_532),
.Y(n_413)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_461),
.B(n_496),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_444),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_416),
.B(n_444),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_432),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_417),
.A2(n_432),
.B1(n_433),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.A3(n_422),
.B1(n_424),
.B2(n_427),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_453),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_454),
.C(n_460),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_460),
.Y(n_453)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_474),
.B(n_495),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_472),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_472),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_490),
.B(n_494),
.Y(n_474)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_481),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_487),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_491),
.B(n_493),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_498),
.B(n_499),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_514),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_510),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_510),
.C(n_514),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_503),
.Y(n_539)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_530),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_530),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_527),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_535),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_534),
.B(n_535),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_540),
.B1(n_541),
.B2(n_544),
.Y(n_535)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_536),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_537),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_540),
.C(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_549),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_567),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_554),
.A2(n_574),
.B(n_575),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_559),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_555),
.B(n_559),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_563),
.C(n_564),
.Y(n_559)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_560),
.Y(n_572)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_561),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_564),
.A2(n_565),
.B1(n_570),
.B2(n_571),
.Y(n_569)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_SL g567 ( 
.A(n_568),
.B(n_569),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_569),
.Y(n_574)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);


endmodule