module fake_jpeg_31783_n_261 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_17),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_0),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_68),
.Y(n_89)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_63),
.Y(n_87)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_66),
.Y(n_91)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_0),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_25),
.B1(n_32),
.B2(n_24),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_25),
.B1(n_32),
.B2(n_39),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_74)
);

AND2x4_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_0),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_88),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_81),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_34),
.B1(n_35),
.B2(n_21),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_95),
.B1(n_105),
.B2(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_92),
.Y(n_111)
);

HAxp5_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_33),
.CON(n_88),
.SN(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_23),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_26),
.B1(n_22),
.B2(n_4),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_26),
.B1(n_22),
.B2(n_4),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_101),
.B(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_15),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_13),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_5),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_11),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_125),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_11),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_72),
.B1(n_104),
.B2(n_119),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_128),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_119),
.Y(n_141)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_55),
.B1(n_3),
.B2(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_2),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_75),
.B1(n_101),
.B2(n_83),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_137),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_77),
.B1(n_96),
.B2(n_99),
.Y(n_147)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_89),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_73),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_100),
.C(n_87),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_149),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_117),
.B(n_126),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_77),
.C(n_96),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_72),
.B1(n_76),
.B2(n_104),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_159),
.B1(n_110),
.B2(n_123),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_76),
.B(n_104),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_169),
.B(n_171),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_154),
.B(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_116),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_178),
.B1(n_145),
.B2(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_110),
.C(n_113),
.Y(n_175)
);

OAI211xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_184),
.B(n_185),
.C(n_144),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_120),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_124),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_188),
.B(n_146),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_153),
.B1(n_147),
.B2(n_143),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_194),
.B1(n_196),
.B2(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_190),
.A2(n_201),
.B(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_159),
.B1(n_141),
.B2(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_172),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_159),
.B1(n_162),
.B2(n_142),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_198),
.C(n_186),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_159),
.B1(n_142),
.B2(n_156),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_166),
.C(n_181),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_107),
.B1(n_155),
.B2(n_150),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_192),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_176),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_200),
.C(n_199),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_168),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_179),
.A3(n_173),
.B1(n_182),
.B2(n_174),
.C1(n_185),
.C2(n_177),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_217),
.A3(n_197),
.B1(n_214),
.B2(n_201),
.C1(n_192),
.C2(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_188),
.B(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_161),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

AO221x1_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_132),
.B1(n_133),
.B2(n_137),
.C(n_206),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_222),
.B(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_195),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_198),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_191),
.B1(n_196),
.B2(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_240),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_209),
.B1(n_216),
.B2(n_215),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_221),
.B1(n_232),
.B2(n_238),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_229),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_208),
.B(n_218),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_231),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_213),
.B1(n_220),
.B2(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_245),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_223),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_246),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_249),
.B(n_237),
.CI(n_235),
.CON(n_251),
.SN(n_251)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_254),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_247),
.B(n_244),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_251),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_259),
.C(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_256),
.Y(n_261)
);


endmodule