module fake_jpeg_12301_n_312 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_14),
.B(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_9),
.B1(n_3),
.B2(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_23),
.B1(n_52),
.B2(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_27),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_47),
.B(n_51),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_49),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_55),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_17),
.A2(n_26),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_60),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_62),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_10),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_88),
.Y(n_97)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_3),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_80),
.Y(n_101)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_27),
.B(n_1),
.Y(n_73)
);

OR2x4_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_25),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_5),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_81),
.Y(n_130)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_33),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_90),
.A2(n_117),
.B1(n_122),
.B2(n_64),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_28),
.B1(n_34),
.B2(n_32),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_108),
.B1(n_115),
.B2(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_37),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_112),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_76),
.B1(n_74),
.B2(n_45),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_42),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_28),
.B1(n_34),
.B2(n_32),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_126),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_42),
.B1(n_40),
.B2(n_34),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_32),
.B1(n_31),
.B2(n_35),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_115),
.B1(n_106),
.B2(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_6),
.Y(n_126)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_81),
.B(n_25),
.CON(n_128),
.SN(n_128)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_138),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_47),
.B(n_25),
.C(n_11),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_12),
.C(n_16),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_67),
.B(n_12),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_95),
.A2(n_78),
.B1(n_50),
.B2(n_48),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_153),
.B1(n_159),
.B2(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_130),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_48),
.B1(n_50),
.B2(n_58),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_145),
.A2(n_179),
.B(n_167),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_157),
.Y(n_192)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_58),
.B1(n_64),
.B2(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_167),
.B1(n_165),
.B2(n_181),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_1),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_16),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_101),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_180),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_111),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_152),
.C(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_168),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_94),
.B1(n_102),
.B2(n_131),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_91),
.A2(n_129),
.B1(n_133),
.B2(n_127),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_176),
.B1(n_162),
.B2(n_142),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_102),
.B1(n_131),
.B2(n_137),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_174),
.B1(n_180),
.B2(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_98),
.B(n_129),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_91),
.A2(n_100),
.B1(n_132),
.B2(n_114),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_104),
.B1(n_135),
.B2(n_90),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_104),
.B(n_97),
.Y(n_180)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_104),
.A2(n_118),
.B1(n_73),
.B2(n_117),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_163),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_89),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_173),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_145),
.B1(n_179),
.B2(n_143),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_191),
.B1(n_193),
.B2(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_153),
.B1(n_181),
.B2(n_148),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_211),
.B1(n_189),
.B2(n_210),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_206),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_163),
.A2(n_160),
.B1(n_144),
.B2(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_210),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_140),
.A2(n_149),
.B1(n_151),
.B2(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_215),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_178),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_146),
.C(n_155),
.Y(n_217)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_227),
.C(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_195),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_238),
.C(n_190),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_196),
.C(n_214),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_196),
.B(n_198),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_185),
.B(n_197),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_184),
.B(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_185),
.B(n_197),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_241),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_194),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_247),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_205),
.B(n_188),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_254),
.B(n_255),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_205),
.C(n_202),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_256),
.B(n_223),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_221),
.A3(n_228),
.B1(n_224),
.B2(n_225),
.C1(n_219),
.C2(n_232),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_230),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_233),
.B(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_266),
.B(n_268),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_241),
.C(n_253),
.Y(n_274)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_229),
.B1(n_218),
.B2(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_251),
.A2(n_220),
.B1(n_216),
.B2(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_234),
.B1(n_250),
.B2(n_248),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_255),
.B1(n_248),
.B2(n_243),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_278),
.B1(n_262),
.B2(n_270),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_253),
.CI(n_240),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_256),
.C(n_247),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_280),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_254),
.B1(n_245),
.B2(n_244),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_242),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_244),
.C(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_283),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_279),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_278),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_271),
.Y(n_294)
);

A2O1A1O1Ixp25_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_257),
.B(n_258),
.C(n_263),
.D(n_266),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_252),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_293),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_271),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_286),
.B(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_287),
.Y(n_301)
);

OAI21x1_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_272),
.B(n_290),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_307),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_298),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_305),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_309),
.C(n_272),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_291),
.Y(n_312)
);


endmodule