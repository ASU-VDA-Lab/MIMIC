module fake_jpeg_29713_n_120 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_2),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_37),
.Y(n_43)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_18),
.B1(n_14),
.B2(n_24),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_45),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_18),
.B1(n_14),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_55),
.B1(n_11),
.B2(n_7),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_68),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_32),
.B(n_30),
.C(n_38),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_65),
.B(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_42),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_29),
.B1(n_34),
.B2(n_30),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_24),
.Y(n_69)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_43),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_59),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_84),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_59),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_95),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_65),
.C(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_96),
.C(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_60),
.C(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_94),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_79),
.C(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

AO221x1_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_103),
.B1(n_85),
.B2(n_102),
.C(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_64),
.C(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_81),
.B1(n_88),
.B2(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_108),
.A3(n_74),
.B1(n_68),
.B2(n_53),
.C1(n_54),
.C2(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_71),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_61),
.B1(n_42),
.B2(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_111),
.C(n_112),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_110),
.C(n_42),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_116),
.B(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_10),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_10),
.Y(n_120)
);


endmodule