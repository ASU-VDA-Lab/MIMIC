module fake_jpeg_13987_n_550 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_550);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_10),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_59),
.B(n_103),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_18),
.B1(n_10),
.B2(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_64),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_34),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_68),
.B(n_49),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_23),
.A2(n_10),
.B(n_17),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_95),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_97),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_22),
.B(n_11),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_45),
.Y(n_141)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_29),
.B(n_11),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_26),
.B1(n_28),
.B2(n_21),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_109),
.A2(n_112),
.B1(n_119),
.B2(n_122),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_40),
.B1(n_28),
.B2(n_45),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_110),
.A2(n_121),
.B(n_144),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_28),
.B1(n_50),
.B2(n_48),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_51),
.B1(n_50),
.B2(n_48),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_40),
.B1(n_33),
.B2(n_45),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_51),
.B1(n_38),
.B2(n_36),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g196 ( 
.A(n_132),
.B(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_66),
.A2(n_33),
.B1(n_45),
.B2(n_43),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_52),
.A2(n_42),
.B1(n_45),
.B2(n_43),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_162),
.B1(n_166),
.B2(n_54),
.Y(n_206)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_82),
.Y(n_155)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_42),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_21),
.B1(n_25),
.B2(n_27),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_52),
.A2(n_42),
.B1(n_43),
.B2(n_20),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_104),
.A2(n_35),
.B1(n_49),
.B2(n_30),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_25),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_168),
.B(n_173),
.Y(n_231)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_171),
.Y(n_238)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_30),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_95),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_174),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_221),
.Y(n_276)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_178),
.Y(n_270)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_117),
.Y(n_179)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_110),
.A2(n_70),
.B1(n_96),
.B2(n_91),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_180),
.A2(n_206),
.B1(n_222),
.B2(n_62),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_116),
.B(n_100),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_182),
.B(n_194),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_27),
.B1(n_37),
.B2(n_41),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_120),
.B(n_105),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_186),
.B(n_212),
.C(n_217),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_37),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_195),
.Y(n_234)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

BUFx4f_ASAP7_75t_SL g246 ( 
.A(n_188),
.Y(n_246)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_109),
.A2(n_69),
.B1(n_57),
.B2(n_87),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_191),
.A2(n_192),
.B1(n_226),
.B2(n_160),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_162),
.B1(n_121),
.B2(n_153),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_41),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_106),
.B(n_90),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_113),
.Y(n_197)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_199),
.B(n_208),
.Y(n_275)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_73),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_209),
.Y(n_251)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_123),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_214),
.Y(n_265)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_131),
.B(n_100),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_164),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_218),
.Y(n_239)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_114),
.B(n_42),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_114),
.B(n_78),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_219),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_154),
.A2(n_42),
.B1(n_43),
.B2(n_78),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_225),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_85),
.B1(n_81),
.B2(n_74),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_228),
.B1(n_161),
.B2(n_145),
.Y(n_233)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_107),
.A2(n_72),
.B1(n_67),
.B2(n_65),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_149),
.A2(n_63),
.B1(n_61),
.B2(n_43),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_237),
.A2(n_242),
.B1(n_250),
.B2(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_186),
.B(n_145),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_240),
.B(n_252),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_142),
.B1(n_107),
.B2(n_126),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_241),
.A2(n_245),
.B1(n_248),
.B2(n_255),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_186),
.A2(n_148),
.B(n_62),
.C(n_129),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_207),
.B(n_212),
.C(n_209),
.D(n_215),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_142),
.B1(n_126),
.B2(n_163),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_169),
.A2(n_151),
.B1(n_115),
.B2(n_147),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_181),
.A2(n_147),
.B1(n_11),
.B2(n_3),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_169),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_0),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_0),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_12),
.C(n_17),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_212),
.C(n_178),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_191),
.A2(n_12),
.B1(n_17),
.B2(n_5),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_174),
.A2(n_12),
.B(n_16),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_273),
.A2(n_13),
.B(n_6),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_183),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_233),
.B1(n_245),
.B2(n_248),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_281),
.A2(n_324),
.B(n_326),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_271),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_283),
.A2(n_280),
.B1(n_238),
.B2(n_256),
.Y(n_340)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_286),
.B(n_287),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_175),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_247),
.C(n_269),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_234),
.B(n_203),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_290),
.B(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_197),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_239),
.B(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_300),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_255),
.A2(n_207),
.B(n_179),
.C(n_223),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_296),
.A2(n_279),
.B(n_246),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_189),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_297),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_199),
.B(n_201),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_232),
.B(n_244),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_177),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_226),
.B1(n_205),
.B2(n_188),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_301),
.A2(n_304),
.B1(n_311),
.B2(n_312),
.Y(n_361)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_250),
.B1(n_237),
.B2(n_267),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_303),
.A2(n_306),
.B1(n_314),
.B2(n_232),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_231),
.B(n_198),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_310),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_267),
.A2(n_172),
.B1(n_193),
.B2(n_200),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_231),
.B(n_170),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_323),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_251),
.B(n_216),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_171),
.B1(n_214),
.B2(n_210),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_259),
.A2(n_230),
.B1(n_240),
.B2(n_276),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_317),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_185),
.B1(n_190),
.B2(n_204),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_275),
.B(n_221),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_220),
.B1(n_6),
.B2(n_8),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_238),
.B1(n_280),
.B2(n_261),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_13),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_270),
.Y(n_354)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_236),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_321),
.Y(n_357)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_325),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_273),
.B(n_13),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_1),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_18),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_247),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_330),
.A2(n_337),
.B1(n_314),
.B2(n_309),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_331),
.B(n_338),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_332),
.A2(n_351),
.B(n_326),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_335),
.A2(n_345),
.B1(n_355),
.B2(n_304),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_289),
.A2(n_268),
.B1(n_258),
.B2(n_253),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_340),
.A2(n_292),
.B1(n_309),
.B2(n_298),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_356),
.C(n_297),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_295),
.A2(n_278),
.B1(n_258),
.B2(n_256),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_347),
.B(n_302),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_263),
.B(n_269),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_367),
.B(n_281),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_295),
.A2(n_238),
.B1(n_263),
.B2(n_262),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_359),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_303),
.A2(n_243),
.B1(n_262),
.B2(n_235),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_277),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_294),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_297),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_364),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_282),
.B(n_279),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_362),
.B(n_363),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_266),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_235),
.Y(n_364)
);

AOI22x1_ASAP7_75t_SL g367 ( 
.A1(n_284),
.A2(n_246),
.B1(n_266),
.B2(n_270),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_246),
.C(n_243),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_246),
.C(n_8),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_353),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_371),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_353),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_357),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_372),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_313),
.B1(n_292),
.B2(n_306),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_374),
.A2(n_376),
.B(n_379),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_394),
.C(n_403),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_378),
.A2(n_382),
.B(n_384),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_289),
.B(n_296),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_380),
.A2(n_388),
.B1(n_393),
.B2(n_398),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_326),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_316),
.Y(n_383)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_349),
.A2(n_324),
.B(n_287),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_357),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_387),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_335),
.A2(n_312),
.B1(n_318),
.B2(n_286),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_328),
.B(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_345),
.A2(n_351),
.B1(n_355),
.B2(n_333),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_325),
.C(n_307),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_296),
.B1(n_322),
.B2(n_321),
.Y(n_396)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_334),
.A2(n_296),
.B(n_323),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_329),
.A2(n_296),
.B1(n_243),
.B2(n_291),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_399),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_392),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_365),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_401),
.B(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_402),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_18),
.B1(n_8),
.B2(n_9),
.Y(n_404)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_358),
.A2(n_6),
.B1(n_14),
.B2(n_15),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_330),
.B1(n_366),
.B2(n_369),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_406),
.B(n_409),
.Y(n_442)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_412),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_334),
.Y(n_416)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_386),
.B(n_343),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_386),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_341),
.C(n_339),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_423),
.C(n_430),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_362),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_433),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_363),
.C(n_360),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_427),
.A2(n_378),
.B1(n_379),
.B2(n_382),
.Y(n_461)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_428),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_342),
.C(n_344),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_397),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_400),
.C(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_389),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_347),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_368),
.C(n_369),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_403),
.C(n_381),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_377),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_441),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_377),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_348),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_444),
.B(n_449),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_380),
.B1(n_393),
.B2(n_373),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_445),
.A2(n_456),
.B1(n_373),
.B2(n_407),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_406),
.B(n_381),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_448),
.B(n_450),
.Y(n_470)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_348),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_376),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_452),
.C(n_458),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_381),
.C(n_387),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_425),
.A2(n_374),
.B1(n_391),
.B2(n_401),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_453),
.A2(n_455),
.B1(n_459),
.B2(n_461),
.Y(n_482)
);

CKINVDCx14_ASAP7_75t_R g486 ( 
.A(n_454),
.Y(n_486)
);

XNOR2x1_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_396),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_419),
.A2(n_373),
.B1(n_398),
.B2(n_371),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_460),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_372),
.C(n_370),
.Y(n_458)
);

XNOR2x1_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_403),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_402),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g463 ( 
.A(n_410),
.B(n_384),
.CI(n_367),
.CON(n_463),
.SN(n_463)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_431),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_404),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_414),
.C(n_417),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_466),
.B(n_479),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_440),
.A2(n_434),
.B1(n_425),
.B2(n_427),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_467),
.B(n_468),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_424),
.C(n_417),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_469),
.A2(n_477),
.B1(n_480),
.B2(n_464),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_424),
.C(n_429),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_481),
.C(n_484),
.Y(n_495)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_446),
.Y(n_474)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_474),
.Y(n_488)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_475),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_445),
.A2(n_407),
.B1(n_435),
.B2(n_415),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_456),
.A2(n_418),
.B1(n_411),
.B2(n_434),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_424),
.C(n_418),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_443),
.A2(n_409),
.B1(n_453),
.B2(n_437),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_483),
.A2(n_405),
.B1(n_458),
.B2(n_463),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_438),
.B(n_411),
.C(n_431),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_426),
.C(n_350),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_459),
.C(n_448),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_491),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_439),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_493),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_469),
.A2(n_450),
.B1(n_441),
.B2(n_442),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_484),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_463),
.B1(n_455),
.B2(n_451),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_477),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_497),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_482),
.A2(n_457),
.B1(n_350),
.B2(n_336),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_501),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_350),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_499),
.B(n_503),
.Y(n_510)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_480),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_475),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_336),
.B1(n_346),
.B2(n_16),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_500),
.A2(n_472),
.B(n_465),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_515),
.B(n_497),
.Y(n_520)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_500),
.B(n_495),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_511),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_517),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_487),
.A2(n_501),
.B(n_496),
.C(n_471),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_491),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_516),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_495),
.A2(n_465),
.B(n_468),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_504),
.B(n_478),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_481),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_470),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_476),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_509),
.B(n_517),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_476),
.C(n_466),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_522),
.Y(n_531)
);

AO21x1_ASAP7_75t_L g522 ( 
.A1(n_518),
.A2(n_487),
.B(n_489),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_505),
.A2(n_488),
.B1(n_502),
.B2(n_494),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_529),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_505),
.A2(n_493),
.B(n_503),
.Y(n_525)
);

AOI21xp33_ASAP7_75t_L g537 ( 
.A1(n_525),
.A2(n_514),
.B(n_470),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_512),
.B(n_488),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_526),
.B(n_494),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_532),
.B(n_527),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_535),
.Y(n_539)
);

AO21x1_ASAP7_75t_L g534 ( 
.A1(n_523),
.A2(n_511),
.B(n_510),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_534),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_528),
.B(n_514),
.C(n_519),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_525),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_538),
.A2(n_530),
.B(n_536),
.Y(n_542)
);

OAI21x1_ASAP7_75t_SL g543 ( 
.A1(n_541),
.A2(n_534),
.B(n_531),
.Y(n_543)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_542),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_544),
.C(n_522),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_528),
.C(n_535),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_545),
.B(n_540),
.C(n_521),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_546),
.B(n_346),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_14),
.B(n_15),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_14),
.C(n_15),
.Y(n_550)
);


endmodule