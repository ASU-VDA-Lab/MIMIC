module fake_jpeg_12637_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_11),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_7),
.B(n_2),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_57),
.C(n_33),
.Y(n_86)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_6),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_17),
.B(n_5),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_66),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_10),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_69),
.Y(n_89)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_10),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_24),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_21),
.B1(n_34),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_81),
.B1(n_98),
.B2(n_49),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_77),
.B1(n_65),
.B2(n_64),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_21),
.B1(n_34),
.B2(n_30),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_78),
.A2(n_99),
.B(n_23),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_92),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_4),
.Y(n_128)
);

HAxp5_ASAP7_75t_SL g87 ( 
.A(n_41),
.B(n_26),
.CON(n_87),
.SN(n_87)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_0),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_102),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_27),
.B1(n_26),
.B2(n_0),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_26),
.B1(n_39),
.B2(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_11),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_26),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_112),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_80),
.B1(n_100),
.B2(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_114),
.B(n_123),
.Y(n_160)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_116),
.A2(n_133),
.B1(n_138),
.B2(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_142),
.B1(n_145),
.B2(n_87),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_3),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_136),
.C(n_139),
.Y(n_154)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_3),
.B(n_4),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_44),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_11),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_13),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_46),
.B1(n_61),
.B2(n_23),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_23),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_143),
.Y(n_149)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_73),
.A2(n_23),
.B1(n_90),
.B2(n_104),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_81),
.B1(n_98),
.B2(n_101),
.Y(n_156)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_72),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_171),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_82),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_91),
.B1(n_101),
.B2(n_110),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_164),
.B1(n_166),
.B2(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_97),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_165),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_91),
.B1(n_107),
.B2(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_80),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_161),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_134),
.C(n_142),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_121),
.C(n_125),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_181),
.B1(n_188),
.B2(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_166),
.B1(n_170),
.B2(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_145),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_127),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_113),
.B1(n_115),
.B2(n_124),
.Y(n_188)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_130),
.B1(n_139),
.B2(n_140),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_155),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_201),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_197),
.B1(n_183),
.B2(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_196),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_164),
.B1(n_158),
.B2(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_182),
.B1(n_172),
.B2(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_200),
.B1(n_181),
.B2(n_175),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_202),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_149),
.B1(n_151),
.B2(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_167),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_152),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

OA21x2_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_176),
.B(n_177),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_193),
.C(n_199),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_210),
.C(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_193),
.C(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_216),
.C(n_221),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_202),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_195),
.B(n_185),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_192),
.B(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_178),
.C(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_213),
.B1(n_209),
.B2(n_211),
.Y(n_222)
);

AOI22x1_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_217),
.B1(n_207),
.B2(n_206),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_224),
.B(n_192),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_227),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_213),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_230),
.B(n_232),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_186),
.B(n_184),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_226),
.A2(n_189),
.B(n_154),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_160),
.C(n_189),
.Y(n_231)
);

AOI31xp67_ASAP7_75t_SL g236 ( 
.A1(n_231),
.A2(n_188),
.A3(n_179),
.B(n_152),
.Y(n_236)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_234),
.B(n_235),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_226),
.B(n_225),
.C(n_160),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_147),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_237),
.B(n_147),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_240),
.B(n_162),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_146),
.C(n_162),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_146),
.Y(n_242)
);


endmodule