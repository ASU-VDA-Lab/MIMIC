module fake_jpeg_7052_n_277 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_277);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_39),
.B1(n_43),
.B2(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_13),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_13),
.B1(n_22),
.B2(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_27),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_44),
.C(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_59),
.Y(n_63)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_30),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_36),
.B1(n_40),
.B2(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_36),
.B1(n_40),
.B2(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_38),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_38),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.C(n_53),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_64),
.B1(n_71),
.B2(n_57),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_59),
.B(n_50),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_73),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_86),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_58),
.B1(n_49),
.B2(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_90),
.B1(n_96),
.B2(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_60),
.B1(n_36),
.B2(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_93),
.Y(n_105)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_53),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_36),
.B1(n_40),
.B2(n_37),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_91),
.B1(n_88),
.B2(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_104),
.B(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_111),
.B1(n_95),
.B2(n_39),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_76),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_70),
.A3(n_76),
.B1(n_53),
.B2(n_68),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_66),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_82),
.C(n_45),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_70),
.B1(n_68),
.B2(n_62),
.Y(n_111)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_53),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_115),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_27),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_133),
.B1(n_101),
.B2(n_51),
.Y(n_154)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_125),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_136),
.B1(n_23),
.B2(n_13),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.C(n_106),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_45),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_45),
.C(n_21),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_109),
.C(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_134),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_54),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_51),
.B1(n_57),
.B2(n_41),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_21),
.B(n_19),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_116),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_155),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_77),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_149),
.C(n_157),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_161),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_146),
.B(n_41),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_104),
.C(n_98),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_66),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_51),
.B1(n_41),
.B2(n_92),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_104),
.C(n_100),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_30),
.C(n_42),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_61),
.C(n_56),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_131),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_66),
.B(n_29),
.Y(n_171)
);

XOR2x2_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_43),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_170),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_119),
.B(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_47),
.B1(n_77),
.B2(n_16),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_153),
.B1(n_151),
.B2(n_148),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_171),
.B1(n_18),
.B2(n_16),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_61),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_157),
.B1(n_41),
.B2(n_25),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_66),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_56),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_30),
.C(n_33),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_33),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_33),
.C(n_32),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_194),
.B(n_20),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_197),
.C(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_33),
.C(n_32),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_47),
.C(n_29),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_47),
.B1(n_20),
.B2(n_16),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_179),
.B1(n_170),
.B2(n_176),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_202),
.A2(n_162),
.B1(n_177),
.B2(n_183),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_28),
.C(n_22),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_15),
.C(n_1),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_177),
.B1(n_24),
.B2(n_20),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_217),
.B1(n_203),
.B2(n_9),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_28),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_186),
.B(n_192),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_24),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_197),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_0),
.Y(n_214)
);

XOR2x1_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_217),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_15),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_2),
.C(n_3),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_0),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_231),
.Y(n_243)
);

AOI21x1_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_214),
.B(n_206),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_188),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_229),
.B(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_188),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_204),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_198),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_235),
.C(n_204),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_9),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_244),
.C(n_226),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_227),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_211),
.B1(n_219),
.B2(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_3),
.B(n_4),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_15),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_4),
.C(n_15),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_15),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_9),
.B(n_5),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_7),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_10),
.C(n_6),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_256),
.A2(n_241),
.B(n_238),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_264),
.B(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_262),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_249),
.B(n_8),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_15),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_4),
.B(n_7),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_255),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_270),
.C(n_12),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_10),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_7),
.B(n_10),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_272),
.B(n_11),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_266),
.C(n_11),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_12),
.Y(n_277)
);


endmodule