module fake_jpeg_1072_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_0),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_68),
.B1(n_71),
.B2(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_95),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_68),
.B1(n_71),
.B2(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_49),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_65),
.B1(n_69),
.B2(n_58),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_52),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_74),
.B1(n_50),
.B2(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_80),
.B1(n_54),
.B2(n_73),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_80),
.B1(n_60),
.B2(n_78),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_72),
.Y(n_104)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_70),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_78),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_64),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_63),
.Y(n_110)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_123),
.B1(n_124),
.B2(n_133),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_73),
.B1(n_49),
.B2(n_63),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_110),
.B1(n_97),
.B2(n_99),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_66),
.B1(n_55),
.B2(n_53),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_0),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_56),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_56),
.B(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_5),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_139),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_142),
.B(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_115),
.C(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_6),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_6),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_151),
.B(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_23),
.B1(n_44),
.B2(n_43),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_150),
.B1(n_154),
.B2(n_14),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_118),
.B1(n_114),
.B2(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_7),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_130),
.B1(n_22),
.B2(n_24),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_8),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_115),
.B(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_12),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_169),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_141),
.B1(n_150),
.B2(n_140),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_174),
.B1(n_175),
.B2(n_17),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_139),
.B(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_184),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_45),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_18),
.C(n_19),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_16),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_185),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_169),
.B1(n_170),
.B2(n_26),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_30),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_162),
.B(n_164),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_165),
.B(n_159),
.C(n_169),
.D(n_160),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_198),
.B1(n_188),
.B2(n_186),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_189),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_169),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_181),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_193),
.B1(n_199),
.B2(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_208),
.B(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_209),
.C(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_196),
.C(n_21),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_20),
.B(n_27),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_29),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_32),
.Y(n_216)
);


endmodule