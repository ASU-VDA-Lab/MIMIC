module fake_jpeg_1077_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_75),
.Y(n_87)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_72),
.Y(n_90)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_62),
.B1(n_50),
.B2(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_62),
.B1(n_76),
.B2(n_53),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_62),
.B1(n_65),
.B2(n_64),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_67),
.B1(n_66),
.B2(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_57),
.C(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_61),
.C(n_51),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_103),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_105),
.B1(n_107),
.B2(n_61),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_49),
.B(n_77),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_109),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_76),
.B1(n_92),
.B2(n_79),
.Y(n_105)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_1),
.C(n_2),
.Y(n_124)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_0),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_126),
.B1(n_107),
.B2(n_93),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_39),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_11),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_37),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_107),
.B1(n_97),
.B2(n_108),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_9),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_10),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.C(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_11),
.Y(n_145)
);

XOR2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_25),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_12),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_121),
.C(n_28),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_171),
.C(n_155),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_159),
.Y(n_180)
);

NOR4xp25_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_23),
.C(n_35),
.D(n_34),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_160),
.B(n_166),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_12),
.B(n_13),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_13),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_26),
.B(n_32),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_147),
.C(n_146),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_178),
.C(n_167),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_30),
.C(n_31),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_168),
.C(n_36),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

AOI321xp33_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_156),
.A3(n_171),
.B1(n_160),
.B2(n_170),
.C(n_168),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_177),
.B1(n_174),
.B2(n_176),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_16),
.B(n_17),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_182),
.A2(n_172),
.B(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.C(n_184),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_18),
.C(n_19),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_16),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_18),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_19),
.Y(n_198)
);


endmodule