module fake_jpeg_12557_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_51),
.Y(n_87)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_7),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_3),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_64),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_3),
.C(n_4),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_29),
.C(n_35),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_21),
.A2(n_3),
.B(n_4),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_17),
.B1(n_18),
.B2(n_39),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_80),
.B1(n_31),
.B2(n_30),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_97),
.C(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_93),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_18),
.B1(n_17),
.B2(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_96),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_37),
.B1(n_23),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_38),
.B1(n_64),
.B2(n_46),
.Y(n_121)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_23),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_63),
.B1(n_57),
.B2(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_35),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_7),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_37),
.B1(n_24),
.B2(n_22),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_114),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_37),
.B1(n_31),
.B2(n_30),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_117),
.B1(n_123),
.B2(n_74),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_20),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_24),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_33),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_53),
.B1(n_38),
.B2(n_25),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_121),
.B1(n_132),
.B2(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_64),
.B1(n_55),
.B2(n_52),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_76),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_55),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_90),
.C(n_77),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_126),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_52),
.B1(n_46),
.B2(n_9),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_119),
.C(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_86),
.B1(n_101),
.B2(n_67),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_145),
.B1(n_131),
.B2(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_68),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_153),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_124),
.B1(n_122),
.B2(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_91),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_92),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_157),
.Y(n_165)
);

AO22x2_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_84),
.B1(n_94),
.B2(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_160),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_107),
.B1(n_125),
.B2(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_173),
.B1(n_145),
.B2(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_134),
.C(n_152),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_111),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_140),
.B(n_156),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_169),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_157),
.B1(n_129),
.B2(n_12),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_130),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_108),
.B1(n_116),
.B2(n_128),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_116),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_176),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_105),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_151),
.A3(n_158),
.B1(n_146),
.B2(n_157),
.C1(n_15),
.C2(n_16),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_129),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_151),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_179),
.B(n_135),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_177),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_186),
.C(n_195),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_152),
.C(n_136),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_136),
.B1(n_141),
.B2(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_192),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_170),
.Y(n_205)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_158),
.B1(n_146),
.B2(n_140),
.C(n_157),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_175),
.A3(n_167),
.B1(n_176),
.B2(n_174),
.C1(n_170),
.C2(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_166),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_157),
.C(n_11),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_8),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_164),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_165),
.B1(n_161),
.B2(n_173),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_203),
.B(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_167),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_164),
.B(n_178),
.C(n_169),
.D(n_171),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_182),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_160),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_215),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_185),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_229),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_199),
.B(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_225),
.B(n_228),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_209),
.B1(n_199),
.B2(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_196),
.B1(n_195),
.B2(n_194),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_226),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_234),
.B(n_235),
.Y(n_238)
);

HAxp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_187),
.CON(n_235),
.SN(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_223),
.B(n_184),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_183),
.B1(n_192),
.B2(n_230),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_241),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_8),
.C(n_14),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_226),
.B(n_164),
.C(n_159),
.Y(n_240)
);

OAI21x1_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_8),
.B(n_14),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_159),
.B1(n_14),
.B2(n_15),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_15),
.B(n_16),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_238),
.B(n_237),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_242),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_16),
.Y(n_248)
);


endmodule