module fake_netlist_1_8325_n_31 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_31);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g10 ( .A(n_1), .B(n_5), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g11 ( .A(n_3), .B(n_6), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_5), .Y(n_15) );
OR2x2_ASAP7_75t_SL g16 ( .A(n_13), .B(n_2), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_13), .B(n_2), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_14), .B(n_4), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_12), .B1(n_10), .B2(n_15), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_18), .B1(n_20), .B2(n_21), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_16), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_14), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_12), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI322xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_6), .A3(n_7), .B1(n_9), .B2(n_11), .C1(n_22), .C2(n_12), .Y(n_27) );
XNOR2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_11), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_28), .Y(n_30) );
AOI22xp5_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_28), .B1(n_12), .B2(n_29), .Y(n_31) );
endmodule