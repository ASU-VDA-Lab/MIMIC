module fake_netlist_1_8573_n_29 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_4), .B(n_0), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx16_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_2), .B(n_8), .Y(n_14) );
OR2x6_ASAP7_75t_SL g15 ( .A(n_13), .B(n_0), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_9), .B(n_1), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_16), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_14), .Y(n_21) );
OAI211xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B(n_20), .C(n_14), .Y(n_22) );
OAI22xp33_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_15), .B1(n_11), .B2(n_4), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OAI21xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .B(n_11), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_27), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
endmodule