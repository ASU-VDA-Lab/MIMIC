module fake_jpeg_13128_n_537 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_537);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_22),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_67),
.B(n_99),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g162 ( 
.A(n_71),
.Y(n_162)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_74),
.A2(n_44),
.B1(n_56),
.B2(n_53),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_79),
.Y(n_126)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_81),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_82),
.B(n_101),
.Y(n_171)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_0),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_23),
.Y(n_106)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_116),
.Y(n_190)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_119),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_120),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_1),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_19),
.B(n_44),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_19),
.B1(n_27),
.B2(n_36),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_128),
.A2(n_146),
.B1(n_154),
.B2(n_174),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_33),
.B1(n_56),
.B2(n_53),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_131),
.A2(n_161),
.B1(n_199),
.B2(n_200),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_138),
.B(n_139),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_31),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_54),
.B(n_46),
.C(n_57),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_140),
.B(n_148),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_26),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_26),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_152),
.B(n_153),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_20),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_77),
.A2(n_20),
.B1(n_52),
.B2(n_48),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_37),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_78),
.A2(n_37),
.B1(n_41),
.B2(n_52),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_48),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_81),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_45),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_91),
.A2(n_57),
.B(n_54),
.C(n_46),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_188),
.A2(n_51),
.B1(n_12),
.B2(n_13),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_79),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_194),
.B(n_143),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_89),
.A2(n_42),
.B1(n_51),
.B2(n_5),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_94),
.A2(n_51),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_97),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_103),
.B(n_2),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_203),
.Y(n_290)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_204),
.Y(n_301)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_189),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_207),
.A2(n_259),
.B(n_270),
.Y(n_319)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_208),
.Y(n_318)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_209),
.Y(n_283)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_211),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_214),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_173),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_216),
.B(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_217),
.Y(n_303)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_192),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_220),
.B(n_252),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_126),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_221),
.B(n_224),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_140),
.B(n_6),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_223),
.B(n_258),
.Y(n_273)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_125),
.A2(n_118),
.B1(n_104),
.B2(n_69),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_225),
.A2(n_227),
.B1(n_235),
.B2(n_257),
.Y(n_302)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_125),
.A2(n_66),
.B1(n_63),
.B2(n_62),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_142),
.Y(n_229)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_130),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_231),
.B(n_245),
.Y(n_299)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_141),
.A2(n_75),
.B1(n_51),
.B2(n_11),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_234),
.A2(n_254),
.B1(n_225),
.B2(n_227),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_195),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_151),
.Y(n_240)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_243),
.Y(n_281)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_266),
.Y(n_298)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_247),
.B(n_248),
.Y(n_320)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_51),
.B1(n_12),
.B2(n_14),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_250),
.A2(n_256),
.B1(n_160),
.B2(n_134),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_167),
.B(n_8),
.C(n_12),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_235),
.Y(n_305)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_124),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_171),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_255),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_127),
.A2(n_15),
.B1(n_202),
.B2(n_191),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_126),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_188),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_263),
.Y(n_280)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_261),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_186),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_190),
.B(n_123),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_186),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_265),
.Y(n_289)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_269),
.B(n_203),
.Y(n_312)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_182),
.B(n_163),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_311),
.B(n_315),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_180),
.B1(n_191),
.B2(n_183),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_278),
.A2(n_279),
.B1(n_294),
.B2(n_297),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_228),
.A2(n_180),
.B1(n_129),
.B2(n_132),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_207),
.A2(n_128),
.B(n_162),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_293),
.B(n_311),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_215),
.A2(n_129),
.B1(n_132),
.B2(n_196),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_222),
.A2(n_160),
.B1(n_196),
.B2(n_197),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_304),
.A2(n_307),
.B1(n_290),
.B2(n_301),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_219),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_246),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_306),
.A2(n_316),
.B1(n_297),
.B2(n_321),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_251),
.A2(n_163),
.B(n_181),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_321),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_210),
.A2(n_213),
.B(n_238),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_256),
.B(n_234),
.Y(n_321)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_344),
.C(n_352),
.Y(n_375)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_327),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_249),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_328),
.B(n_330),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_279),
.A2(n_250),
.B1(n_267),
.B2(n_226),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_329),
.A2(n_351),
.B1(n_356),
.B2(n_290),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_247),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_298),
.A2(n_236),
.B1(n_257),
.B2(n_264),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_331),
.A2(n_332),
.B1(n_339),
.B2(n_347),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_241),
.B1(n_262),
.B2(n_237),
.Y(n_332)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_294),
.A2(n_261),
.B1(n_230),
.B2(n_239),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_298),
.A2(n_266),
.B1(n_269),
.B2(n_220),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_245),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_354),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_285),
.B(n_282),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_342),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_232),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_302),
.A2(n_209),
.B1(n_268),
.B2(n_273),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_348),
.A2(n_350),
.B1(n_355),
.B2(n_358),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_277),
.A2(n_286),
.B(n_321),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_271),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_305),
.B(n_315),
.C(n_285),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_353),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_306),
.B1(n_293),
.B2(n_273),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_286),
.A2(n_301),
.B1(n_312),
.B2(n_303),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_288),
.A2(n_287),
.B1(n_291),
.B2(n_317),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_313),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_357),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_303),
.A2(n_287),
.B1(n_320),
.B2(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_361),
.Y(n_367)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_274),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_386),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_320),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_373),
.C(n_378),
.Y(n_410)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_271),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_338),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_346),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_344),
.C(n_351),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_291),
.B1(n_308),
.B2(n_296),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_383),
.A2(n_343),
.B1(n_324),
.B2(n_326),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_274),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_353),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_309),
.C(n_281),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_313),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_360),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_395),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_411),
.C(n_375),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_398),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_384),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_403),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_341),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_400),
.B(n_394),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_366),
.A2(n_360),
.B(n_349),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_401),
.A2(n_406),
.B(n_407),
.Y(n_431)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_402),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_377),
.B(n_355),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_413),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_348),
.B(n_350),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_347),
.B(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_409),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_375),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_374),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_414),
.Y(n_438)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_419),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_331),
.B1(n_332),
.B2(n_339),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_369),
.B1(n_365),
.B2(n_376),
.Y(n_425)
);

AOI21x1_ASAP7_75t_L g417 ( 
.A1(n_386),
.A2(n_357),
.B(n_361),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_417),
.A2(n_422),
.B(n_372),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_418),
.A2(n_388),
.B1(n_394),
.B2(n_363),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_383),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_362),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_423),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_393),
.A2(n_343),
.B(n_327),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_427),
.B(n_275),
.C(n_310),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_400),
.A2(n_392),
.B1(n_369),
.B2(n_365),
.Y(n_428)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_364),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_442),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_432),
.A2(n_422),
.B(n_412),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_433),
.B(n_448),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_406),
.A2(n_376),
.B1(n_388),
.B2(n_390),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_443),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_435),
.A2(n_439),
.B1(n_440),
.B2(n_416),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_389),
.C(n_379),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_437),
.C(n_417),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_372),
.C(n_385),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_419),
.A2(n_393),
.B1(n_385),
.B2(n_372),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_418),
.A2(n_391),
.B1(n_381),
.B2(n_382),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_359),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_403),
.A2(n_381),
.B1(n_391),
.B2(n_323),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_308),
.B1(n_345),
.B2(n_337),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_446),
.A2(n_399),
.B1(n_408),
.B2(n_398),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_453),
.C(n_458),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

AO221x1_ASAP7_75t_L g452 ( 
.A1(n_431),
.A2(n_407),
.B1(n_423),
.B2(n_414),
.C(n_415),
.Y(n_452)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_452),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_421),
.C(n_397),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_440),
.Y(n_483)
);

NOR2x1_ASAP7_75t_R g457 ( 
.A(n_426),
.B(n_401),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_466),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_421),
.C(n_397),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_461),
.A2(n_444),
.B(n_447),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_404),
.Y(n_462)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_409),
.C(n_396),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_470),
.C(n_426),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_435),
.A2(n_396),
.B1(n_420),
.B2(n_402),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_441),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_284),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_296),
.B1(n_275),
.B2(n_281),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_431),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_469),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_313),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_478),
.Y(n_491)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_451),
.A2(n_447),
.B1(n_430),
.B2(n_444),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_485),
.B1(n_464),
.B2(n_450),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_441),
.C(n_434),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_479),
.B(n_481),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_455),
.C(n_458),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_448),
.C(n_430),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_482),
.B(n_463),
.Y(n_489)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_460),
.A2(n_438),
.B1(n_443),
.B2(n_424),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_484),
.A2(n_460),
.B1(n_474),
.B2(n_480),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_489),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_473),
.A2(n_468),
.B(n_466),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_493),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_461),
.B(n_453),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_469),
.C(n_456),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_487),
.C(n_471),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g496 ( 
.A(n_475),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_496),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_477),
.Y(n_498)
);

OAI321xp33_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_457),
.A3(n_482),
.B1(n_483),
.B2(n_485),
.C(n_471),
.Y(n_508)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_483),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_497),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_495),
.A2(n_456),
.B1(n_459),
.B2(n_462),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_500),
.A2(n_509),
.B1(n_472),
.B2(n_446),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_508),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_486),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_510),
.Y(n_514)
);

OAI21x1_ASAP7_75t_SL g512 ( 
.A1(n_507),
.A2(n_472),
.B(n_438),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_490),
.A2(n_494),
.B1(n_491),
.B2(n_481),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_486),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_506),
.A2(n_505),
.B1(n_507),
.B2(n_504),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_515),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_424),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_517),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_310),
.Y(n_517)
);

A2O1A1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_503),
.A2(n_292),
.B(n_314),
.C(n_295),
.Y(n_518)
);

INVx11_ASAP7_75t_L g520 ( 
.A(n_518),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_292),
.C(n_276),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_519),
.B(n_501),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_501),
.C(n_510),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_283),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_514),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_514),
.A2(n_276),
.B(n_318),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_517),
.B(n_518),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_528),
.B(n_529),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_525),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_530),
.A2(n_524),
.B(n_520),
.Y(n_532)
);

AOI21x1_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_531),
.B(n_520),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_523),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_523),
.C(n_318),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_322),
.B(n_295),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_322),
.Y(n_537)
);


endmodule