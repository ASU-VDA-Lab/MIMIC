module fake_jpeg_2700_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_48),
.Y(n_60)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_46),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_25),
.B2(n_24),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_67),
.B1(n_64),
.B2(n_55),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_26),
.CI(n_25),
.CON(n_56),
.SN(n_56)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_70),
.A3(n_64),
.B1(n_59),
.B2(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_14),
.B1(n_20),
.B2(n_19),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_66),
.B1(n_73),
.B2(n_8),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_70),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_6),
.C(n_7),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_69),
.C(n_70),
.Y(n_92)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_39),
.CON(n_76),
.SN(n_76)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_46),
.B1(n_45),
.B2(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_61),
.B1(n_56),
.B2(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_62),
.Y(n_105)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_69),
.C(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_74),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_74),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_54),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_68),
.B(n_54),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_102),
.B(n_103),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_89),
.C(n_94),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_62),
.B(n_65),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_84),
.B(n_91),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_65),
.B(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_80),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_118),
.C(n_101),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_104),
.Y(n_125)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_110),
.B1(n_98),
.B2(n_97),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_122),
.C(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_99),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_107),
.C(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_104),
.B1(n_95),
.B2(n_106),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_113),
.B1(n_111),
.B2(n_117),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_120),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_125),
.B(n_126),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_128),
.B(n_131),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.C(n_127),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_127),
.B(n_129),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_124),
.B(n_119),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);


endmodule