module fake_jpeg_9393_n_77 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_2),
.B(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_31),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_12),
.B(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_0),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_52),
.B(n_42),
.C(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_0),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

CKINVDCx11_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_48),
.B(n_46),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_63),
.B1(n_44),
.B2(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_15),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_14),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_68),
.B(n_59),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_60),
.C(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_63),
.B1(n_17),
.B2(n_19),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_16),
.C(n_22),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_23),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_34),
.B(n_25),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_26),
.Y(n_77)
);


endmodule