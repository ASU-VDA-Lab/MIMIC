module fake_jpeg_16082_n_335 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_58),
.Y(n_101)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_67),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_27),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx9p33_ASAP7_75t_R g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_12),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_33),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_86),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_17),
.C(n_35),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_0),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_16),
.B1(n_14),
.B2(n_23),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_78),
.A2(n_92),
.B(n_105),
.Y(n_140)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_18),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_83),
.B(n_99),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_18),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_100),
.Y(n_122)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_39),
.A2(n_44),
.B1(n_40),
.B2(n_50),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_91),
.B1(n_112),
.B2(n_115),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_114),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_37),
.B1(n_26),
.B2(n_33),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_36),
.B1(n_29),
.B2(n_13),
.Y(n_137)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_38),
.A2(n_15),
.B1(n_37),
.B2(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_107),
.B(n_108),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_36),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_36),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_46),
.A2(n_35),
.B1(n_29),
.B2(n_17),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_48),
.A2(n_35),
.B1(n_29),
.B2(n_17),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_13),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_130),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_121),
.B(n_137),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_135),
.Y(n_168)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_36),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_131),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_134),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_13),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_11),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_84),
.A2(n_11),
.B1(n_12),
.B2(n_2),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_136),
.A2(n_145),
.B1(n_162),
.B2(n_70),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_77),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_146),
.Y(n_166)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_161),
.B1(n_151),
.B2(n_130),
.Y(n_173)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_79),
.A2(n_12),
.B1(n_1),
.B2(n_3),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_34),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_34),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_34),
.B(n_1),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_7),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx2_ASAP7_75t_R g153 ( 
.A(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_0),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_1),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_159),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_69),
.B(n_3),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_4),
.Y(n_159)
);

OR2x2_ASAP7_75t_SL g160 ( 
.A(n_72),
.B(n_4),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_102),
.A2(n_4),
.B1(n_7),
.B2(n_94),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_89),
.A2(n_7),
.B1(n_70),
.B2(n_82),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g227 ( 
.A(n_173),
.B(n_90),
.C(n_143),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_75),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_182),
.B(n_168),
.Y(n_234)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_75),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_124),
.B(n_112),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_185),
.B(n_136),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_82),
.B(n_87),
.C(n_89),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_117),
.B(n_73),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_192),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_142),
.B1(n_126),
.B2(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_121),
.C(n_118),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_213),
.C(n_189),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_140),
.B1(n_126),
.B2(n_162),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_206),
.A2(n_211),
.B1(n_223),
.B2(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_171),
.A2(n_151),
.B(n_142),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_214),
.B(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_131),
.C(n_150),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_157),
.B(n_156),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_145),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_216),
.B(n_226),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_180),
.A2(n_72),
.B1(n_141),
.B2(n_144),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_228),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_152),
.B1(n_139),
.B2(n_123),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_187),
.B1(n_186),
.B2(n_175),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_163),
.A2(n_127),
.B1(n_160),
.B2(n_123),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_139),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_234),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

AOI221xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_187),
.B1(n_175),
.B2(n_186),
.C(n_195),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_90),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_163),
.A2(n_196),
.B1(n_173),
.B2(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_197),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_169),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_239),
.C(n_241),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_169),
.B(n_168),
.C(n_176),
.D(n_172),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_249),
.B(n_251),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_169),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_246),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_194),
.C(n_198),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_199),
.C(n_202),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_207),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_260),
.C(n_210),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_256),
.B(n_220),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_170),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_211),
.A2(n_201),
.B1(n_167),
.B2(n_165),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_262),
.B1(n_263),
.B2(n_227),
.Y(n_278)
);

BUFx4f_ASAP7_75t_SL g259 ( 
.A(n_203),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_259),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_199),
.C(n_167),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_206),
.A2(n_165),
.B1(n_183),
.B2(n_200),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_215),
.A2(n_223),
.B1(n_222),
.B2(n_216),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_212),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_270),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_259),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_243),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_274),
.B(n_286),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_275),
.C(n_282),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_224),
.C(n_214),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_233),
.B(n_204),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_253),
.B1(n_251),
.B2(n_247),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_285),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_219),
.A3(n_204),
.B1(n_233),
.B2(n_221),
.C1(n_229),
.C2(n_218),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_261),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_225),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_218),
.C(n_230),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_230),
.C(n_225),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_241),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_250),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_242),
.B(n_253),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_266),
.C(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XOR2x2_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_263),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_262),
.B1(n_258),
.B2(n_260),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_244),
.B1(n_238),
.B2(n_220),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_276),
.A2(n_209),
.B1(n_228),
.B2(n_203),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_271),
.B(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_269),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_293),
.B(n_287),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_282),
.C(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_308),
.Y(n_318)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_275),
.C(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_265),
.B(n_272),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_286),
.C(n_285),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_311),
.B(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_281),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_316),
.B(n_303),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_298),
.B(n_288),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_319),
.B(n_268),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_300),
.B1(n_265),
.B2(n_296),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_312),
.C(n_301),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_292),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_304),
.Y(n_326)
);

NOR2x1_ASAP7_75t_R g329 ( 
.A(n_322),
.B(n_326),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_324),
.B(n_317),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_270),
.B(n_267),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_327),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_306),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_314),
.B(n_283),
.C(n_267),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_283),
.B(n_203),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_332),
.C(n_170),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_326),
.Y(n_335)
);


endmodule