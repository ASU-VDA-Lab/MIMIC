module fake_jpeg_1257_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_7),
.B(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_43),
.B(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_48),
.Y(n_82)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_62),
.Y(n_104)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_66),
.Y(n_83)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_65),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_29),
.B(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_77),
.Y(n_105)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_30),
.B(n_2),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_24),
.B(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_4),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_76),
.Y(n_90)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_3),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_81),
.Y(n_119)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_45),
.A2(n_27),
.B1(n_40),
.B2(n_39),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_32),
.B1(n_40),
.B2(n_39),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_23),
.B1(n_38),
.B2(n_41),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_101),
.B1(n_106),
.B2(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_111),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_21),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_102),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_9),
.B1(n_59),
.B2(n_56),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_97),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_9),
.B1(n_52),
.B2(n_77),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_47),
.B1(n_49),
.B2(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_43),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_45),
.A2(n_34),
.B1(n_42),
.B2(n_50),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_36),
.B1(n_79),
.B2(n_66),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_43),
.B(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_122),
.Y(n_180)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_99),
.Y(n_123)
);

HAxp5_ASAP7_75t_SL g176 ( 
.A(n_123),
.B(n_131),
.CON(n_176),
.SN(n_176)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_115),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_87),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_96),
.B1(n_93),
.B2(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_141),
.B1(n_146),
.B2(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_115),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_147),
.Y(n_157)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_125),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_90),
.B1(n_114),
.B2(n_95),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_152),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_85),
.B1(n_94),
.B2(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_115),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_151),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_107),
.B(n_100),
.C(n_110),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_107),
.B(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_91),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_110),
.B1(n_91),
.B2(n_108),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_167),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_134),
.B1(n_128),
.B2(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_128),
.A2(n_145),
.B1(n_140),
.B2(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_171),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_172),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_179),
.B1(n_173),
.B2(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_191),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_140),
.B(n_150),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_163),
.B(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_126),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_201),
.C(n_210),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_211),
.B1(n_213),
.B2(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_163),
.B(n_150),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_209),
.B(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_162),
.C(n_177),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_173),
.B1(n_161),
.B2(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_170),
.B1(n_159),
.B2(n_139),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_221),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_218),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_192),
.B(n_187),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_212),
.B1(n_184),
.B2(n_202),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_188),
.C(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_188),
.B1(n_186),
.B2(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_203),
.B1(n_212),
.B2(n_214),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_227),
.A2(n_200),
.B1(n_219),
.B2(n_223),
.Y(n_235)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_206),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_206),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_226),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_235),
.A2(n_226),
.B1(n_231),
.B2(n_230),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_217),
.C(n_210),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_199),
.C(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_200),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_236),
.B(n_233),
.Y(n_243)
);

OAI221xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_225),
.B1(n_234),
.B2(n_182),
.C(n_183),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_247),
.B(n_245),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_242),
.Y(n_249)
);


endmodule