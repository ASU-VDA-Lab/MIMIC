module fake_jpeg_21210_n_31 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_31);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

AND2x2_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx2_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_5),
.B(n_10),
.C(n_13),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

AO21x2_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_17),
.B(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_27),
.B(n_28),
.Y(n_30)
);

AOI211xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_24),
.B(n_25),
.C(n_23),
.Y(n_31)
);


endmodule