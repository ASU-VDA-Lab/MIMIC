module fake_jpeg_5835_n_244 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_19),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_25),
.B1(n_19),
.B2(n_28),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_52),
.B1(n_57),
.B2(n_59),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_25),
.B1(n_36),
.B2(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_27),
.B1(n_34),
.B2(n_21),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_24),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_33),
.B1(n_28),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_31),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_71),
.B(n_78),
.Y(n_99)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_59),
.B1(n_65),
.B2(n_23),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_24),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_18),
.B1(n_29),
.B2(n_17),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_84),
.B1(n_86),
.B2(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_81),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_48),
.B(n_29),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_29),
.B1(n_17),
.B2(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_48),
.B1(n_62),
.B2(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_20),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_41),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_102),
.B(n_80),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_85),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_110),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_54),
.B1(n_63),
.B2(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_113),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_54),
.C(n_15),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_77),
.B1(n_73),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_124),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_123),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_111),
.B1(n_90),
.B2(n_110),
.Y(n_142)
);

BUFx6f_ASAP7_75t_SL g127 ( 
.A(n_92),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_69),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_102),
.B(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_141),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_101),
.C(n_102),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_156),
.B1(n_136),
.B2(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_111),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_111),
.B(n_95),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_80),
.B1(n_112),
.B2(n_74),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_134),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_15),
.B1(n_98),
.B2(n_6),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_3),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_138),
.B1(n_151),
.B2(n_153),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_120),
.A3(n_116),
.B1(n_118),
.B2(n_130),
.C1(n_124),
.C2(n_122),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_116),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_120),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_74),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_120),
.C(n_6),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_183),
.B1(n_154),
.B2(n_145),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_147),
.C(n_157),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_138),
.B1(n_142),
.B2(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_139),
.C(n_140),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_158),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_188),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_186),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_137),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_166),
.C(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_195),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_206),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_165),
.C(n_194),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_199),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_191),
.B(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_167),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_209),
.C(n_204),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_204),
.B(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_171),
.B(n_172),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_171),
.B(n_172),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_150),
.B1(n_178),
.B2(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_127),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_182),
.C(n_188),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_185),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_195),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_216),
.A2(n_207),
.B(n_6),
.C(n_8),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_196),
.C(n_186),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_92),
.C(n_98),
.Y(n_218)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_226),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_216),
.B1(n_9),
.B2(n_10),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_5),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_8),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_8),
.B(n_9),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_222),
.B1(n_11),
.B2(n_12),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_10),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_10),
.B(n_11),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_238),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_235),
.A3(n_229),
.B1(n_232),
.B2(n_12),
.C1(n_13),
.C2(n_11),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_12),
.C(n_13),
.Y(n_244)
);


endmodule