module fake_jpeg_24112_n_264 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_152;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx8_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_32),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_18),
.Y(n_62)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_48),
.B(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_63),
.Y(n_91)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_53),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_30),
.B(n_27),
.C(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_55),
.B(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_20),
.B1(n_27),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_65),
.B(n_80),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_30),
.B(n_34),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_29),
.B1(n_34),
.B2(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_72),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_21),
.B1(n_35),
.B2(n_31),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_73),
.B(n_77),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_21),
.B1(n_35),
.B2(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_18),
.B1(n_36),
.B2(n_31),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_18),
.B1(n_36),
.B2(n_33),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_38),
.A2(n_35),
.B1(n_26),
.B2(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_25),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_97),
.B1(n_100),
.B2(n_52),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_105),
.B1(n_112),
.B2(n_64),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_36),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_96),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_24),
.C(n_23),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_6),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_24),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_23),
.B1(n_19),
.B2(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_115),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_19),
.B1(n_28),
.B2(n_32),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_51),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_78),
.C(n_79),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_51),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_73),
.B1(n_69),
.B2(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_5),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_69),
.B1(n_72),
.B2(n_49),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_118),
.A2(n_134),
.B1(n_137),
.B2(n_140),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_125),
.B(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_126),
.A2(n_128),
.B1(n_139),
.B2(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_52),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_85),
.B1(n_64),
.B2(n_86),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_60),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_107),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_141),
.B1(n_104),
.B2(n_101),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_60),
.B1(n_8),
.B2(n_9),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_6),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_145),
.C(n_95),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_88),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_16),
.B1(n_11),
.B2(n_12),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_10),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_111),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_154),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_96),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_110),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_159),
.Y(n_179)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_172),
.B(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_96),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_145),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_141),
.B(n_109),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_91),
.C(n_92),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_129),
.C(n_109),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_109),
.Y(n_176)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_178),
.B(n_185),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_175),
.B(n_160),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_122),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_190),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_163),
.B(n_172),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_186),
.B(n_187),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_137),
.B(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_91),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_129),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_197),
.C(n_176),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_134),
.B(n_122),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_112),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_200),
.C(n_205),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_165),
.C(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_179),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_167),
.B1(n_160),
.B2(n_155),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_206),
.B1(n_212),
.B2(n_213),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_175),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_209),
.C(n_197),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_165),
.C(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_105),
.B1(n_150),
.B2(n_171),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_171),
.B1(n_157),
.B2(n_156),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_188),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_222),
.Y(n_229)
);

NOR2x1_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_194),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_224),
.B(n_181),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_226),
.C(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_184),
.C(n_197),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_195),
.B1(n_193),
.B2(n_177),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_181),
.B1(n_182),
.B2(n_190),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_221),
.C(n_228),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_211),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_239),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_212),
.B1(n_206),
.B2(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_201),
.B1(n_189),
.B2(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_237),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_220),
.B(n_217),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_205),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_187),
.B(n_178),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_200),
.C(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.C(n_247),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_218),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_224),
.A3(n_234),
.B1(n_187),
.B2(n_237),
.C1(n_239),
.C2(n_184),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_191),
.C(n_219),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_238),
.B(n_232),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_252),
.B(n_182),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_152),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_248),
.C(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_257),
.C(n_186),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_158),
.B1(n_251),
.B2(n_101),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_260),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_92),
.B(n_89),
.Y(n_261)
);

OAI311xp33_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_89),
.A3(n_104),
.B1(n_133),
.C1(n_262),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_104),
.Y(n_264)
);


endmodule