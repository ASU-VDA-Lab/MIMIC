module real_jpeg_5832_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_1),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_124),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_1),
.A2(n_124),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_3),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_4),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_77),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_5),
.A2(n_43),
.B1(n_244),
.B2(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_5),
.A2(n_43),
.B1(n_92),
.B2(n_282),
.Y(n_281)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_7),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_142),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_8),
.A2(n_65),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_8),
.B(n_246),
.C(n_250),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_8),
.B(n_23),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_8),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_8),
.B(n_133),
.Y(n_284)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_11),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_11),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_11),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_12),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_12),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_13),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_14),
.A2(n_50),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_14),
.A2(n_50),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_14),
.A2(n_50),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_228),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_226),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_157),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_18),
.B(n_157),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_98),
.C(n_134),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_19),
.A2(n_20),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_21),
.B(n_64),
.C(n_72),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_36),
.B(n_44),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_22),
.A2(n_36),
.B1(n_54),
.B2(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_22),
.B(n_46),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_55),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_25),
.Y(n_140)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_29),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_29),
.Y(n_244)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_32),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_32),
.Y(n_223)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_32),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_37),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_39),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_39),
.Y(n_217)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_53),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_47),
.B(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_49),
.Y(n_164)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_53),
.A2(n_305),
.B(n_307),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_58),
.Y(n_142)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_175),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_65),
.A2(n_166),
.B(n_174),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_65),
.A2(n_178),
.B(n_260),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_SL g305 ( 
.A1(n_65),
.A2(n_216),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_66),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_66),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_79),
.B1(n_88),
.B2(n_95),
.Y(n_72)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_79),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_86),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_89),
.Y(n_259)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_96),
.A2(n_152),
.B(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_98),
.B(n_134),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_119),
.B(n_125),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_99),
.A2(n_125),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_99),
.A2(n_119),
.B1(n_219),
.B2(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_100),
.B(n_126),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_104),
.Y(n_222)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_106),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_110),
.A2(n_224),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_116),
.B2(n_118),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_116),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_146),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_135),
.B(n_146),
.Y(n_308)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.A3(n_139),
.B1(n_141),
.B2(n_143),
.Y(n_135)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_144),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_141),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_151),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_153),
.B(n_181),
.Y(n_260)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_194),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_176),
.B2(n_177),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.A3(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_183),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_178),
.A2(n_255),
.B(n_260),
.Y(n_254)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_211),
.B2(n_225),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_204),
.B(n_205),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B(n_224),
.Y(n_218)
);

INVx5_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AO21x1_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_310),
.B(n_315),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_297),
.B(n_309),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_270),
.B(n_296),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_253),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_232),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_241),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_233),
.A2(n_241),
.B1(n_242),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_262),
.C(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_268),
.B2(n_269),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_286),
.B(n_295),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_279),
.B(n_285),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_284),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_293),
.Y(n_295)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_299),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_308),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.C(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);


endmodule