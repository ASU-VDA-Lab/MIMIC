module fake_jpeg_27663_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_9),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_7),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_11),
.B2(n_14),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_10),
.C(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_31),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_10),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_27),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_42),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_44),
.B(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_33),
.B(n_34),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_41),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_14),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_43),
.C(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_58),
.B1(n_57),
.B2(n_51),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_0),
.C(n_1),
.Y(n_54)
);

BUFx24_ASAP7_75t_SL g60 ( 
.A(n_55),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_12),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.C(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_50),
.B1(n_10),
.B2(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_5),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.A3(n_8),
.B1(n_2),
.B2(n_3),
.C1(n_1),
.C2(n_32),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_32),
.B1(n_40),
.B2(n_3),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_1),
.C(n_3),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_67),
.B(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);


endmodule