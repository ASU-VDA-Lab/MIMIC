module fake_jpeg_26260_n_287 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_20),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_20),
.C(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_41),
.B1(n_32),
.B2(n_33),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_15),
.B1(n_31),
.B2(n_30),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_33),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_38),
.B(n_46),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_40),
.B1(n_44),
.B2(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_36),
.C(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_62),
.Y(n_72)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_20),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_41),
.B1(n_38),
.B2(n_47),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_39),
.B1(n_55),
.B2(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_79),
.B1(n_86),
.B2(n_78),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_40),
.B1(n_41),
.B2(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_47),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_29),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_39),
.B1(n_26),
.B2(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_92),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_104),
.B(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_99),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_60),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_61),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_62),
.B1(n_59),
.B2(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_76),
.B1(n_81),
.B2(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_0),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_109),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_82),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_99),
.B(n_100),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_125),
.B1(n_104),
.B2(n_71),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_122),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_84),
.C(n_29),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_67),
.Y(n_154)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_79),
.B1(n_68),
.B2(n_74),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_127),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_93),
.B(n_98),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_139),
.B(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_151),
.B(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_138),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_95),
.B1(n_106),
.B2(n_74),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_125),
.B1(n_123),
.B2(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_126),
.B1(n_120),
.B2(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_58),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_106),
.B1(n_74),
.B2(n_71),
.Y(n_146)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_45),
.B(n_27),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_30),
.B(n_67),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_145),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_114),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_161),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_176),
.B(n_144),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_108),
.C(n_29),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_165),
.C(n_172),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_108),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_179),
.B(n_174),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_30),
.B(n_71),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_174),
.B(n_0),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_175),
.B1(n_177),
.B2(n_146),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_58),
.B1(n_45),
.B2(n_54),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_171),
.B1(n_150),
.B2(n_130),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_45),
.B1(n_54),
.B2(n_51),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_28),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_12),
.B(n_18),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_66),
.B1(n_51),
.B2(n_52),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_52),
.B1(n_37),
.B2(n_29),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_28),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_149),
.C(n_130),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_197),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_137),
.C(n_136),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_192),
.C(n_158),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_143),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_193),
.B(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_191),
.B(n_195),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_132),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_137),
.C(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_141),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_63),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_0),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_200),
.A2(n_164),
.B1(n_166),
.B2(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_63),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_215),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_168),
.B1(n_167),
.B2(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_207),
.B1(n_213),
.B2(n_214),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_178),
.C(n_161),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_219),
.C(n_28),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_167),
.B1(n_193),
.B2(n_182),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_17),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_172),
.B1(n_37),
.B2(n_63),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_63),
.B1(n_29),
.B2(n_37),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_180),
.B1(n_181),
.B2(n_185),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_1),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_24),
.C(n_34),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_228),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_197),
.B(n_196),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_231),
.B(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_24),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_28),
.B(n_18),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_232),
.C(n_233),
.Y(n_241)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_206),
.B(n_3),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_34),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_34),
.C(n_17),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_216),
.C(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

OAI322xp33_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_220),
.A3(n_212),
.B1(n_209),
.B2(n_219),
.C1(n_217),
.C2(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_240),
.B(n_226),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_244),
.A2(n_247),
.B1(n_5),
.B2(n_7),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_204),
.C(n_34),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_241),
.C(n_244),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_230),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_246),
.B(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_227),
.B1(n_229),
.B2(n_224),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_232),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_256),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_233),
.B1(n_235),
.B2(n_8),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_257),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_12),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_242),
.B(n_239),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_260),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_266),
.B1(n_10),
.B2(n_11),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_241),
.B(n_247),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_7),
.C(n_8),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_5),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_7),
.B(n_8),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_253),
.C(n_258),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_272),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_274),
.B(n_264),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_9),
.B(n_10),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_267),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_264),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_271),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_34),
.B(n_10),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_10),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_11),
.C(n_34),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_11),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_34),
.Y(n_287)
);


endmodule