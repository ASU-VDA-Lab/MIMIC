module fake_jpeg_13625_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_11),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_43),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_21),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_26),
.B1(n_49),
.B2(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_50),
.B1(n_69),
.B2(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_0),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_96),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_20),
.B1(n_47),
.B2(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_92),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_67),
.B1(n_62),
.B2(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_58),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_67),
.B1(n_50),
.B2(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_72),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_71),
.B1(n_57),
.B2(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_59),
.B1(n_63),
.B2(n_51),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_113),
.B1(n_35),
.B2(n_42),
.Y(n_137)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_73),
.C(n_56),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_5),
.C(n_6),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_33),
.B(n_44),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_118),
.Y(n_128)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_114),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_8),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_1),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_6),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_10),
.Y(n_131)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_126),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_132),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_30),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_129),
.C(n_13),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_138),
.B(n_17),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_12),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_10),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_11),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_108),
.B1(n_107),
.B2(n_15),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_29),
.B(n_41),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

NOR4xp25_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_149),
.C(n_150),
.D(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_146),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_12),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_148),
.C(n_151),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

OR2x4_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_39),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_136),
.C(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_157),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_SL g158 ( 
.A1(n_156),
.A2(n_144),
.A3(n_145),
.B1(n_150),
.B2(n_142),
.C1(n_147),
.C2(n_128),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_148),
.B(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_156),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_154),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_161),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_158),
.Y(n_167)
);


endmodule