module real_jpeg_15263_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_0),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_0),
.A2(n_87),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22x1_ASAP7_75t_SL g314 ( 
.A1(n_0),
.A2(n_87),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_0),
.A2(n_87),
.B1(n_229),
.B2(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_52),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_3),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_4),
.B(n_84),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_4),
.A2(n_22),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_22),
.B1(n_157),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_4),
.B(n_332),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_4),
.A2(n_358),
.A3(n_360),
.B1(n_362),
.B2(n_364),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_4),
.B(n_306),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_4),
.B(n_246),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_5),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_5),
.Y(n_306)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_6),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_6),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_6),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_6),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_7),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_8),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_127),
.B1(n_193),
.B2(n_196),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_8),
.A2(n_127),
.B1(n_215),
.B2(n_219),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_10),
.Y(n_231)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_261),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_259),
.Y(n_13)
);

INVxp33_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_222),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_16),
.B(n_222),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_149),
.C(n_199),
.Y(n_16)
);

INVxp67_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_18),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_19),
.B(n_80),
.C(n_121),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_46),
.Y(n_19)
);

XOR2x2_ASAP7_75t_SL g268 ( 
.A(n_20),
.B(n_46),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_36),
.B2(n_39),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_22),
.B(n_106),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_22),
.A2(n_36),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_22),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_22),
.B(n_363),
.Y(n_362)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_23),
.A2(n_120),
.A3(n_290),
.B1(n_292),
.B2(n_297),
.Y(n_289)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_32),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_35),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_38),
.Y(n_142)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_45),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_59),
.B(n_63),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_47),
.A2(n_69),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_51),
.Y(n_388)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_62),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_63),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_64),
.A2(n_227),
.B(n_232),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_65),
.A2(n_203),
.B(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_69),
.B(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_69),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_69),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_71),
.Y(n_205)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_121),
.B2(n_122),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_117),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_81),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_92),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_82),
.B(n_93),
.Y(n_190)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_107),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_92),
.Y(n_254)
);

NOR2x1p5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_105),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_93),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_93),
.B(n_192),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_93),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_100),
.B2(n_102),
.Y(n_93)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_101),
.Y(n_291)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_104),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_114),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_112),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_137),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_124),
.B(n_138),
.Y(n_257)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_130),
.B(n_143),
.Y(n_185)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_130),
.Y(n_274)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_138),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_150),
.B(n_199),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_184),
.C(n_189),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_151),
.A2(n_152),
.B1(n_189),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_165),
.B(n_177),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_153),
.B(n_314),
.Y(n_353)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_160),
.B2(n_163),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_167),
.B1(n_171),
.B2(n_175),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_161),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_164),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_177),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_214),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_165),
.B(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_176),
.Y(n_318)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_177),
.Y(n_312)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_184),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_185),
.B(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_190),
.B(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_211),
.Y(n_199)
);

NAND2x1p5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_211),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_202),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_202),
.B(n_336),
.Y(n_392)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_207),
.Y(n_335)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_212),
.B(n_353),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_213),
.B(n_313),
.Y(n_330)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_250),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g302 ( 
.A1(n_227),
.A2(n_303),
.B(n_307),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_227),
.A2(n_335),
.B(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_231),
.Y(n_361)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp67_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_247),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_249),
.B(n_352),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

XOR2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

AOI21x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B(n_255),
.Y(n_252)
);

NOR2x1p5_ASAP7_75t_SL g349 ( 
.A(n_254),
.B(n_255),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_280),
.B(n_405),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_278),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_264),
.B(n_278),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_265),
.B(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.C(n_275),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_275),
.B1(n_276),
.B2(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_277),
.B(n_378),
.Y(n_390)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_325),
.B(n_404),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_322),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_284),
.B(n_322),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.C(n_308),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_285),
.B(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_288),
.A2(n_308),
.B1(n_309),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_302),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_289),
.A2(n_302),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_398),
.B(n_403),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_354),
.B(n_397),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_341),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_341),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.C(n_333),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_347),
.C(n_350),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_374),
.B(n_396),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_371),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_356),
.B(n_371),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_370),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_370),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_382),
.B(n_395),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_381),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_381),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_391),
.B(n_394),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_390),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_393),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_402),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);


endmodule