module fake_netlist_1_1546_n_792 (n_117, n_44, n_133, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_98, n_74, n_7, n_29, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_139, n_16, n_13, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_145, n_61, n_21, n_99, n_109, n_93, n_132, n_51, n_140, n_96, n_39, n_792, n_769);
input n_117;
input n_44;
input n_133;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_139;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_145;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_51;
input n_140;
input n_96;
input n_39;
output n_792;
output n_769;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_43), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_146), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_41), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_48), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_74), .Y(n_152) );
INVxp67_ASAP7_75t_L g153 ( .A(n_123), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_105), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_73), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_134), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_14), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
INVxp33_ASAP7_75t_SL g161 ( .A(n_126), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_77), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_30), .Y(n_163) );
INVxp33_ASAP7_75t_SL g164 ( .A(n_10), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_80), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_39), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_122), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_14), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_15), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_108), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_70), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_22), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_84), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_121), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_88), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_136), .B(n_102), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_8), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_35), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_81), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_23), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_30), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_92), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_18), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_49), .Y(n_185) );
BUFx5_ASAP7_75t_L g186 ( .A(n_37), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_93), .Y(n_188) );
INVxp33_ASAP7_75t_SL g189 ( .A(n_133), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_15), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_119), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_9), .Y(n_193) );
INVx1_ASAP7_75t_SL g194 ( .A(n_42), .Y(n_194) );
INVxp33_ASAP7_75t_SL g195 ( .A(n_76), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_89), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_71), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_116), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_34), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_67), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_112), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_86), .Y(n_204) );
INVxp67_ASAP7_75t_SL g205 ( .A(n_55), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_120), .Y(n_206) );
INVxp33_ASAP7_75t_SL g207 ( .A(n_47), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_94), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_26), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_87), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_78), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_83), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_75), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_27), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_56), .Y(n_215) );
INVxp33_ASAP7_75t_SL g216 ( .A(n_60), .Y(n_216) );
INVxp33_ASAP7_75t_SL g217 ( .A(n_79), .Y(n_217) );
INVxp67_ASAP7_75t_SL g218 ( .A(n_33), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_54), .Y(n_219) );
INVxp67_ASAP7_75t_SL g220 ( .A(n_46), .Y(n_220) );
INVxp33_ASAP7_75t_L g221 ( .A(n_58), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_11), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_140), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_132), .Y(n_224) );
INVxp33_ASAP7_75t_SL g225 ( .A(n_82), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_143), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_72), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_91), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_106), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_113), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_45), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_12), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_5), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_101), .Y(n_235) );
BUFx2_ASAP7_75t_SL g236 ( .A(n_11), .Y(n_236) );
INVxp33_ASAP7_75t_SL g237 ( .A(n_16), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_118), .Y(n_238) );
INVxp33_ASAP7_75t_SL g239 ( .A(n_139), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_124), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_85), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_33), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_110), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_13), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_37), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_117), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_69), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_135), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_227), .B(n_0), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_186), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_159), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_186), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_240), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_240), .Y(n_256) );
AND2x6_ASAP7_75t_L g257 ( .A(n_192), .B(n_62), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_167), .B(n_0), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_221), .B(n_1), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_150), .Y(n_261) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_154), .A2(n_1), .B(n_2), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_149), .B(n_2), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_148), .A2(n_64), .B(n_63), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_169), .B(n_3), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_149), .B(n_3), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_219), .B(n_4), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_240), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_186), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_192), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_186), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_186), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_240), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_186), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_154), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_248), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_248), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_156), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_156), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_248), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_248), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_248), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_238), .B(n_5), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_249), .B(n_153), .Y(n_285) );
INVx4_ASAP7_75t_L g286 ( .A(n_257), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_251), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_260), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_251), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_257), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_252), .B(n_148), .Y(n_293) );
INVx5_ASAP7_75t_L g294 ( .A(n_257), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_253), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_252), .B(n_188), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_263), .A2(n_147), .B1(n_209), .B2(n_181), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_252), .B(n_197), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_255), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_253), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_254), .Y(n_301) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_250), .A2(n_236), .B1(n_170), .B2(n_171), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_276), .A2(n_166), .B1(n_177), .B2(n_168), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_260), .A2(n_164), .B1(n_216), .B2(n_207), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_265), .B(n_159), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_261), .B(n_150), .Y(n_307) );
BUFx10_ASAP7_75t_L g308 ( .A(n_257), .Y(n_308) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_262), .B(n_165), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_276), .B(n_151), .Y(n_311) );
INVx6_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_261), .B(n_161), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_259), .A2(n_182), .B1(n_242), .B2(n_222), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_257), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_276), .B(n_279), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_279), .A2(n_168), .B1(n_177), .B2(n_166), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_258), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_258), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_257), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_258), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_269), .Y(n_322) );
INVx4_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
AND2x6_ASAP7_75t_L g324 ( .A(n_263), .B(n_165), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_263), .B(n_233), .Y(n_325) );
AND3x2_ASAP7_75t_SL g326 ( .A(n_302), .B(n_184), .C(n_172), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_298), .B(n_279), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_289), .B(n_280), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_296), .A2(n_265), .B1(n_267), .B2(n_250), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_289), .B(n_280), .Y(n_330) );
INVx4_ASAP7_75t_L g331 ( .A(n_324), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_306), .B(n_280), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_312), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_306), .B(n_265), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_285), .B(n_267), .Y(n_336) );
INVx5_ASAP7_75t_L g337 ( .A(n_324), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_297), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_324), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_316), .A2(n_266), .B(n_264), .C(n_269), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_286), .B(n_266), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_312), .Y(n_345) );
INVx5_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_296), .B(n_284), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_313), .B(n_284), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_293), .B(n_266), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_325), .B(n_266), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_308), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_314), .A2(n_297), .B(n_311), .C(n_304), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_325), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_314), .B(n_182), .Y(n_357) );
AND2x6_ASAP7_75t_L g358 ( .A(n_320), .B(n_266), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_325), .B(n_271), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_304), .B(n_264), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_317), .B(n_264), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_317), .B(n_264), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_302), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_286), .Y(n_367) );
BUFx6f_ASAP7_75t_SL g368 ( .A(n_286), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_302), .Y(n_370) );
NAND3xp33_ASAP7_75t_L g371 ( .A(n_305), .B(n_242), .C(n_222), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_302), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_294), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_294), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_292), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_292), .B(n_178), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_315), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_315), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_288), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_323), .B(n_178), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_294), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_323), .B(n_185), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_294), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_291), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_323), .A2(n_237), .B1(n_207), .B2(n_244), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_295), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_295), .B(n_271), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_337), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_354), .A2(n_350), .B(n_364), .C(n_360), .Y(n_390) );
NOR2xp33_ASAP7_75t_R g391 ( .A(n_331), .B(n_202), .Y(n_391) );
BUFx10_ASAP7_75t_L g392 ( .A(n_335), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_331), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_352), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_342), .A2(n_301), .B(n_300), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_352), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_340), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_331), .A2(n_235), .B1(n_189), .B2(n_195), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_338), .A2(n_236), .B1(n_262), .B2(n_214), .Y(n_399) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_371), .B(n_233), .Y(n_400) );
INVx5_ASAP7_75t_L g401 ( .A(n_337), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_356), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_355), .A2(n_262), .B1(n_257), .B2(n_272), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_341), .A2(n_303), .B(n_301), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_334), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_334), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_335), .B(n_205), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_356), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_364), .A2(n_273), .B(n_275), .C(n_272), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_332), .Y(n_410) );
AO21x2_ASAP7_75t_L g411 ( .A1(n_341), .A2(n_171), .B(n_170), .Y(n_411) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_343), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_346), .Y(n_413) );
AO21x1_ASAP7_75t_L g414 ( .A1(n_363), .A2(n_175), .B(n_174), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_347), .B(n_218), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_346), .B(n_294), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_338), .A2(n_231), .B1(n_232), .B2(n_191), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_328), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_357), .B(n_220), .Y(n_419) );
CKINVDCx8_ASAP7_75t_R g420 ( .A(n_358), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_333), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_329), .B(n_163), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_336), .B(n_189), .Y(n_423) );
INVx5_ASAP7_75t_L g424 ( .A(n_358), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_349), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_358), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_359), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_330), .B(n_193), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_386), .B(n_195), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_358), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_327), .B(n_194), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_333), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_351), .B(n_215), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_345), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_361), .A2(n_225), .B1(n_239), .B2(n_217), .Y(n_438) );
BUFx8_ASAP7_75t_L g439 ( .A(n_368), .Y(n_439) );
INVx5_ASAP7_75t_SL g440 ( .A(n_376), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
INVx4_ASAP7_75t_L g442 ( .A(n_358), .Y(n_442) );
OAI22xp33_ASAP7_75t_L g443 ( .A1(n_370), .A2(n_231), .B1(n_232), .B2(n_191), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_362), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_372), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_369), .B(n_365), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_344), .Y(n_447) );
NAND2x2_ASAP7_75t_L g448 ( .A(n_326), .B(n_226), .Y(n_448) );
BUFx8_ASAP7_75t_L g449 ( .A(n_368), .Y(n_449) );
O2A1O1Ixp5_ASAP7_75t_SL g450 ( .A1(n_366), .A2(n_155), .B(n_158), .C(n_157), .Y(n_450) );
NOR2x1_ASAP7_75t_R g451 ( .A(n_381), .B(n_152), .Y(n_451) );
NOR2xp33_ASAP7_75t_R g452 ( .A(n_368), .B(n_152), .Y(n_452) );
O2A1O1Ixp5_ASAP7_75t_L g453 ( .A1(n_388), .A2(n_173), .B(n_208), .C(n_151), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_385), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_387), .Y(n_455) );
BUFx4_ASAP7_75t_SL g456 ( .A(n_326), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_381), .B(n_245), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_383), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_375), .A2(n_318), .B(n_310), .Y(n_459) );
NOR2x1_ASAP7_75t_SL g460 ( .A(n_362), .B(n_174), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_379), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_362), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_374), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_375), .A2(n_257), .B1(n_239), .B2(n_200), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_377), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_390), .A2(n_378), .B(n_377), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_410), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_433), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_457), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_412), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
AOI21x1_ASAP7_75t_L g474 ( .A1(n_414), .A2(n_180), .B(n_179), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_434), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_432), .B(n_319), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_394), .B(n_367), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_446), .A2(n_203), .B1(n_212), .B2(n_204), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_458), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_396), .B(n_367), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_415), .B(n_321), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_391), .A2(n_445), .B1(n_448), .B2(n_398), .Y(n_483) );
AOI322xp5_ASAP7_75t_L g484 ( .A1(n_417), .A2(n_419), .A3(n_422), .B1(n_407), .B2(n_429), .C1(n_430), .C2(n_423), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_390), .A2(n_162), .B(n_196), .C(n_160), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_446), .A2(n_246), .B1(n_322), .B2(n_183), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_420), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_436), .B(n_6), .Y(n_489) );
BUFx8_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_455), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_442), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_409), .A2(n_199), .B(n_201), .C(n_198), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_422), .A2(n_230), .B1(n_187), .B2(n_190), .C1(n_234), .C2(n_241), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_440), .A2(n_229), .B1(n_230), .B2(n_228), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_454), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_443), .A2(n_208), .B(n_223), .C(n_173), .Y(n_497) );
AO31x2_ASAP7_75t_L g498 ( .A1(n_409), .A2(n_256), .A3(n_278), .B(n_270), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_449), .A2(n_210), .B1(n_211), .B2(n_206), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_443), .A2(n_224), .B1(n_243), .B2(n_247), .C(n_213), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_438), .B(n_6), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_442), .B(n_382), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_405), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_392), .B(n_7), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_453), .A2(n_223), .B(n_176), .C(n_256), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_447), .Y(n_507) );
CKINVDCx12_ASAP7_75t_R g508 ( .A(n_451), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_453), .A2(n_270), .B(n_256), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_406), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_424), .B(n_339), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_452), .Y(n_512) );
CKINVDCx8_ASAP7_75t_R g513 ( .A(n_463), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_424), .B(n_348), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_428), .A2(n_278), .B1(n_281), .B2(n_270), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_456), .A2(n_281), .B1(n_278), .B2(n_10), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_424), .B(n_353), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_401), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_399), .A2(n_281), .B1(n_353), .B2(n_268), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_411), .A2(n_353), .B1(n_268), .B2(n_274), .Y(n_520) );
INVx4_ASAP7_75t_L g521 ( .A(n_401), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_400), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_393), .Y(n_523) );
OAI21xp33_ASAP7_75t_L g524 ( .A1(n_464), .A2(n_384), .B(n_373), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_425), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_411), .A2(n_431), .B1(n_402), .B2(n_408), .Y(n_526) );
AND2x6_ASAP7_75t_L g527 ( .A(n_397), .B(n_373), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_427), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_404), .A2(n_268), .B1(n_274), .B2(n_255), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_465), .A2(n_268), .B1(n_274), .B2(n_255), .Y(n_530) );
CKINVDCx8_ASAP7_75t_R g531 ( .A(n_401), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_401), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_459), .A2(n_395), .B(n_403), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_472), .A2(n_435), .B1(n_437), .B2(n_421), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_467), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_483), .A2(n_435), .B1(n_441), .B2(n_437), .Y(n_537) );
OR2x6_ASAP7_75t_L g538 ( .A(n_485), .B(n_397), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_527), .Y(n_539) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_506), .A2(n_486), .B(n_533), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
OAI211xp5_ASAP7_75t_L g542 ( .A1(n_499), .A2(n_389), .B(n_268), .C(n_274), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g543 ( .A1(n_497), .A2(n_462), .B(n_444), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_484), .B(n_450), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_508), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_531), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_469), .B(n_462), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_489), .A2(n_274), .B1(n_277), .B2(n_255), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_533), .A2(n_416), .B(n_299), .Y(n_549) );
OR2x6_ASAP7_75t_L g550 ( .A(n_512), .B(n_17), .Y(n_550) );
AO21x1_ASAP7_75t_L g551 ( .A1(n_516), .A2(n_299), .B(n_287), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_476), .B(n_18), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_491), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_501), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_502), .A2(n_277), .B1(n_282), .B2(n_283), .Y(n_555) );
OR2x6_ASAP7_75t_L g556 ( .A(n_488), .B(n_24), .Y(n_556) );
AO31x2_ASAP7_75t_L g557 ( .A1(n_466), .A2(n_25), .A3(n_28), .B(n_29), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_466), .A2(n_28), .B(n_31), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_494), .B(n_32), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_490), .A2(n_487), .B1(n_505), .B2(n_523), .Y(n_561) );
INVx5_ASAP7_75t_SL g562 ( .A(n_470), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_468), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_521), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_521), .B(n_36), .Y(n_565) );
CKINVDCx6p67_ASAP7_75t_R g566 ( .A(n_513), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_500), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_567) );
OAI21xp33_ASAP7_75t_SL g568 ( .A1(n_496), .A2(n_40), .B(n_41), .Y(n_568) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_509), .A2(n_66), .B(n_65), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_479), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_482), .B(n_44), .Y(n_571) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_474), .A2(n_98), .B(n_145), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_495), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_524), .A2(n_99), .B(n_144), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_471), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_478), .A2(n_51), .B1(n_52), .B2(n_53), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_507), .Y(n_577) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_534), .A2(n_57), .B(n_58), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_480), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_478), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_475), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_477), .Y(n_582) );
BUFx3_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
OR2x6_ASAP7_75t_L g584 ( .A(n_532), .B(n_68), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_559), .A2(n_522), .B1(n_481), .B2(n_519), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_556), .A2(n_492), .B1(n_532), .B2(n_528), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_554), .A2(n_493), .B1(n_526), .B2(n_519), .C(n_515), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_561), .A2(n_525), .B1(n_520), .B2(n_510), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_563), .B(n_504), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_560), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_560), .B(n_498), .Y(n_591) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_549), .A2(n_529), .B(n_530), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_575), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_536), .B(n_498), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_581), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_582), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_570), .B(n_503), .Y(n_597) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_542), .A2(n_517), .B(n_514), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_553), .Y(n_600) );
AO21x2_ASAP7_75t_L g601 ( .A1(n_558), .A2(n_511), .B(n_527), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_539), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_539), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_584), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_557), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_577), .B(n_95), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_552), .B(n_96), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g609 ( .A1(n_537), .A2(n_97), .B1(n_100), .B2(n_103), .C(n_104), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_557), .Y(n_610) );
AO21x2_ASAP7_75t_L g611 ( .A1(n_540), .A2(n_107), .B(n_109), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_541), .B(n_114), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_557), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_540), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_547), .Y(n_615) );
OA21x2_ASAP7_75t_L g616 ( .A1(n_549), .A2(n_127), .B(n_128), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_579), .Y(n_617) );
NAND2xp33_ASAP7_75t_R g618 ( .A(n_550), .B(n_130), .Y(n_618) );
CKINVDCx8_ASAP7_75t_R g619 ( .A(n_545), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_539), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_568), .B(n_578), .C(n_548), .Y(n_621) );
INVx6_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_571), .B(n_544), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_565), .B(n_564), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_576), .A2(n_580), .B(n_573), .C(n_567), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_572), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_564), .B(n_583), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_569), .Y(n_628) );
AO21x2_ASAP7_75t_L g629 ( .A1(n_574), .A2(n_543), .B(n_551), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_562), .B(n_535), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_538), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_605), .Y(n_632) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_604), .Y(n_633) );
AOI31xp33_ASAP7_75t_L g634 ( .A1(n_618), .A2(n_548), .A3(n_555), .B(n_566), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_594), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_589), .B(n_562), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_600), .B(n_569), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_605), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_604), .B(n_594), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_590), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_606), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_617), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_617), .B(n_593), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_606), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_610), .Y(n_645) );
NOR2xp33_ASAP7_75t_SL g646 ( .A(n_619), .B(n_597), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_588), .A2(n_586), .B1(n_623), .B2(n_585), .C(n_597), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_610), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_593), .B(n_595), .Y(n_649) );
OR2x6_ASAP7_75t_L g650 ( .A(n_598), .B(n_630), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_591), .B(n_615), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_625), .A2(n_587), .B1(n_624), .B2(n_621), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_591), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_595), .B(n_596), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_613), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_596), .B(n_615), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_624), .B(n_631), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_614), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_630), .B(n_603), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_614), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_627), .B(n_607), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_607), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_599), .B(n_603), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_608), .B(n_620), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_626), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_601), .B(n_629), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_626), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_601), .B(n_629), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_629), .B(n_602), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_628), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_599), .B(n_603), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_602), .B(n_611), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_628), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_612), .B(n_611), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_611), .B(n_592), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_622), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_592), .B(n_609), .Y(n_677) );
BUFx3_ASAP7_75t_L g678 ( .A(n_622), .Y(n_678) );
BUFx3_ASAP7_75t_L g679 ( .A(n_616), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_594), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_635), .B(n_680), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_640), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_653), .B(n_651), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_635), .B(n_680), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_632), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_639), .B(n_656), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_638), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_651), .B(n_640), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_639), .B(n_656), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_643), .B(n_649), .Y(n_690) );
AO21x1_ASAP7_75t_L g691 ( .A1(n_634), .A2(n_652), .B(n_633), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_641), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_642), .B(n_647), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_645), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_649), .B(n_654), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_645), .Y(n_696) );
INVxp33_ASAP7_75t_L g697 ( .A(n_646), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_654), .B(n_637), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_662), .B(n_657), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_657), .B(n_661), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_648), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_637), .B(n_659), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_664), .B(n_636), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_659), .B(n_669), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_641), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_644), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_644), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_655), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_663), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_671), .B(n_650), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_672), .B(n_668), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_655), .Y(n_712) );
BUFx2_ASAP7_75t_L g713 ( .A(n_663), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_660), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_660), .B(n_658), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_663), .B(n_676), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_658), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_678), .B(n_677), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_665), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_665), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_670), .B(n_673), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_672), .A2(n_675), .B1(n_674), .B2(n_666), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_673), .Y(n_723) );
AOI31xp33_ASAP7_75t_L g724 ( .A1(n_691), .A2(n_667), .A3(n_679), .B(n_697), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_683), .B(n_688), .Y(n_725) );
INVx2_ASAP7_75t_SL g726 ( .A(n_713), .Y(n_726) );
INVx2_ASAP7_75t_SL g727 ( .A(n_713), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_721), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_711), .B(n_698), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_695), .B(n_690), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_699), .B(n_695), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_693), .B(n_700), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_702), .B(n_704), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_703), .B(n_682), .Y(n_734) );
AOI211x1_ASAP7_75t_L g735 ( .A1(n_718), .A2(n_710), .B(n_716), .C(n_704), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_721), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_702), .B(n_686), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_689), .B(n_722), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_681), .B(n_684), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_715), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_709), .Y(n_741) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_709), .B(n_714), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_685), .A2(n_687), .B1(n_714), .B2(n_720), .C(n_719), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_694), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_692), .B(n_712), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_692), .B(n_712), .Y(n_746) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_717), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_717), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_742), .Y(n_749) );
INVx3_ASAP7_75t_L g750 ( .A(n_745), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_744), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_744), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_735), .B(n_696), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_741), .B(n_705), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_729), .B(n_723), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_740), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_748), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_735), .B(n_701), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_725), .B(n_706), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_743), .B(n_707), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_730), .B(n_708), .Y(n_761) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_724), .B(n_708), .Y(n_762) );
XNOR2xp5_ASAP7_75t_L g763 ( .A(n_738), .B(n_731), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_742), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_732), .B(n_734), .Y(n_765) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_726), .B(n_727), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_739), .B(n_728), .Y(n_767) );
XNOR2x1_ASAP7_75t_L g768 ( .A(n_737), .B(n_733), .Y(n_768) );
UNKNOWN g769 ( );
INVx1_ASAP7_75t_L g770 ( .A(n_736), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_746), .B(n_741), .Y(n_771) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_766), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_765), .Y(n_773) );
XNOR2xp5_ASAP7_75t_L g774 ( .A(n_768), .B(n_763), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_SL g775 ( .A1(n_769), .A2(n_758), .B(n_753), .C(n_760), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_757), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_756), .B(n_760), .Y(n_777) );
OA22x2_ASAP7_75t_L g778 ( .A1(n_774), .A2(n_762), .B1(n_764), .B2(n_749), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_775), .B(n_755), .Y(n_779) );
AO22x2_ASAP7_75t_L g780 ( .A1(n_776), .A2(n_764), .B1(n_749), .B2(n_757), .Y(n_780) );
XNOR2x1_ASAP7_75t_L g781 ( .A(n_773), .B(n_767), .Y(n_781) );
OAI211xp5_ASAP7_75t_SL g782 ( .A1(n_777), .A2(n_771), .B(n_750), .C(n_749), .Y(n_782) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_781), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_778), .B(n_772), .Y(n_784) );
NAND3xp33_ASAP7_75t_SL g785 ( .A(n_779), .B(n_772), .C(n_759), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_783), .A2(n_780), .B1(n_782), .B2(n_772), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_786), .A2(n_784), .B1(n_785), .B2(n_770), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_786), .B(n_761), .Y(n_788) );
BUFx2_ASAP7_75t_L g789 ( .A(n_788), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_789), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_790), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_791), .A2(n_787), .B1(n_751), .B2(n_752), .C(n_754), .Y(n_792) );
endmodule