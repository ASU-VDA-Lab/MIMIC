module real_jpeg_24765_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_244;
wire n_167;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_1),
.A2(n_40),
.B1(n_46),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_71),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_40),
.B1(n_46),
.B2(n_71),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_7),
.A2(n_40),
.B1(n_46),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_8),
.A2(n_40),
.B1(n_46),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_8),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_11),
.A2(n_29),
.B1(n_63),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_11),
.A2(n_40),
.B1(n_46),
.B2(n_63),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_12),
.A2(n_35),
.B1(n_66),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_12),
.A2(n_40),
.B1(n_46),
.B2(n_66),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_13),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_13),
.B(n_75),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_56),
.C(n_58),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_111),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_67),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_111),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_13),
.B(n_40),
.C(n_95),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_13),
.A2(n_39),
.B(n_202),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_15),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_99),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_15),
.A2(n_40),
.B1(n_46),
.B2(n_99),
.Y(n_157)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_16),
.B(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_21),
.B(n_114),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_83),
.C(n_101),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_22),
.B(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_23),
.B(n_52),
.C(n_68),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_24),
.B(n_37),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.A3(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_26),
.B(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_29),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_82)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_38),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_39),
.A2(n_86),
.B1(n_88),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_39),
.A2(n_45),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_39),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_39),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_40),
.A2(n_46),
.B1(n_95),
.B2(n_96),
.Y(n_97)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_46),
.B(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_48),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_68),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_64),
.Y(n_52)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_53),
.A2(n_64),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_54),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_54),
.A2(n_138),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_56),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_56),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_67),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_65),
.B(n_108),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B(n_76),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_75),
.B1(n_81),
.B2(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_83),
.B(n_101),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_91),
.Y(n_139)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_90),
.B(n_111),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_92),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_92),
.A2(n_190),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_93),
.A2(n_125),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_98),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_97),
.A2(n_104),
.B(n_175),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_97),
.B(n_111),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_109),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_107),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_245),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_162),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_160),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_145),
.B(n_160),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_146),
.A2(n_147),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_150),
.B(n_151),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_239),
.B(n_244),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_191),
.B(n_238),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_180),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_165),
.B(n_180),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.C(n_177),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_173),
.A2(n_177),
.B1(n_178),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_187),
.C(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_232),
.B(n_237),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_210),
.B(n_231),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_204),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_204),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_199),
.C(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_201),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_220),
.B(n_230),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_218),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_216),
.B(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_225),
.B(n_229),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_243),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);


endmodule