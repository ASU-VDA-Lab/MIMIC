module fake_jpeg_6821_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_36),
.Y(n_62)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_20),
.CON(n_52),
.SN(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_73)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_30),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_58),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_32),
.C(n_16),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_64),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_16),
.B1(n_29),
.B2(n_15),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_59),
.B1(n_60),
.B2(n_19),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_31),
.B1(n_18),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_17),
.B1(n_19),
.B2(n_26),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_17),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_42),
.B1(n_41),
.B2(n_33),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_83),
.B1(n_30),
.B2(n_26),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_84),
.Y(n_90)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_55),
.B1(n_58),
.B2(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_23),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_57),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_19),
.B1(n_18),
.B2(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_102),
.Y(n_118)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_93),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_92),
.B1(n_104),
.B2(n_82),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_98),
.B(n_103),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_56),
.B(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_49),
.B1(n_55),
.B2(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_55),
.B1(n_30),
.B2(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_106),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_128),
.B1(n_104),
.B2(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_119),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_68),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_71),
.C(n_62),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_96),
.C(n_85),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_66),
.C(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_39),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_83),
.B1(n_79),
.B2(n_61),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_88),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_89),
.B1(n_92),
.B2(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_141),
.B1(n_149),
.B2(n_118),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_88),
.C(n_106),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_151),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_109),
.B(n_117),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_100),
.B1(n_85),
.B2(n_91),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_150),
.C(n_116),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_89),
.B1(n_100),
.B2(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_106),
.B1(n_100),
.B2(n_89),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_93),
.B(n_96),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_109),
.B(n_120),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_100),
.B1(n_106),
.B2(n_101),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_88),
.C(n_48),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_103),
.B1(n_79),
.B2(n_61),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_131),
.C(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_151),
.B1(n_143),
.B2(n_144),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_161),
.B(n_162),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_132),
.A2(n_110),
.B(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_146),
.B(n_138),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_107),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_190),
.B1(n_156),
.B2(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_139),
.B1(n_142),
.B2(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_180),
.C(n_185),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_153),
.C(n_131),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_136),
.B1(n_148),
.B2(n_107),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_48),
.C(n_39),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_61),
.B1(n_65),
.B2(n_40),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_152),
.B1(n_162),
.B2(n_163),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_37),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_65),
.B1(n_80),
.B2(n_48),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_37),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

AO221x1_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_80),
.B1(n_48),
.B2(n_154),
.C(n_152),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_24),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_15),
.B1(n_24),
.B2(n_27),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_166),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_176),
.B1(n_183),
.B2(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_199),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_182),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_203),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_172),
.B1(n_48),
.B2(n_18),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_202),
.A2(n_180),
.B1(n_188),
.B2(n_22),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_0),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_31),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_48),
.B1(n_22),
.B2(n_31),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_210),
.B1(n_212),
.B2(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_191),
.C(n_187),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.C(n_214),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_187),
.C(n_181),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_22),
.B1(n_24),
.B2(n_15),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_39),
.C(n_37),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_195),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_224),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_223),
.B(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_226),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_200),
.B(n_198),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_37),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_37),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_0),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_0),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_218),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_234),
.Y(n_243)
);

AOI31xp33_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_210),
.A3(n_211),
.B(n_10),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_10),
.B(n_14),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_211),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_1),
.C(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_227),
.C(n_3),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_239),
.B(n_242),
.Y(n_245)
);

OAI311xp33_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_10),
.A3(n_14),
.B1(n_13),
.C1(n_12),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_241),
.A3(n_11),
.B1(n_12),
.B2(n_6),
.C1(n_4),
.C2(n_5),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_242)
);

OAI221xp5_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_233),
.B1(n_230),
.B2(n_236),
.C(n_237),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_247),
.B(n_4),
.C(n_6),
.Y(n_249)
);

AOI321xp33_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_27),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_245),
.B(n_6),
.Y(n_250)
);

AOI221xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_27),
.B1(n_248),
.B2(n_225),
.C(n_245),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_251),
.Y(n_252)
);


endmodule