module fake_jpeg_18919_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_19),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_0),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_19),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_18),
.B1(n_32),
.B2(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_52),
.B1(n_66),
.B2(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_21),
.B1(n_20),
.B2(n_26),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_63),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_34),
.B1(n_18),
.B2(n_32),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_24),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_21),
.B1(n_26),
.B2(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_30),
.B(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_34),
.B1(n_18),
.B2(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_80),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_85),
.B1(n_92),
.B2(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_43),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_36),
.B1(n_43),
.B2(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_61),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_96),
.B1(n_90),
.B2(n_82),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_103),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_105),
.Y(n_142)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_111),
.Y(n_132)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_43),
.C(n_67),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_43),
.C(n_83),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_91),
.B1(n_46),
.B2(n_50),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_57),
.B(n_55),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_53),
.B1(n_64),
.B2(n_54),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_80),
.B(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_71),
.B(n_33),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_79),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_130),
.Y(n_154)
);

AO21x2_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_80),
.B(n_36),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_131),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_71),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_147),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_151),
.B1(n_114),
.B2(n_105),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_95),
.C(n_87),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_148),
.C(n_124),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_50),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_94),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_36),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_29),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_110),
.B(n_108),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_61),
.B(n_27),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_99),
.B1(n_114),
.B2(n_121),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_89),
.B1(n_17),
.B2(n_23),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_160),
.B1(n_178),
.B2(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_170),
.B1(n_175),
.B2(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_171),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_109),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_177),
.B(n_127),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_110),
.B1(n_108),
.B2(n_106),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_174),
.B1(n_176),
.B2(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_131),
.B(n_33),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_106),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_120),
.B1(n_111),
.B2(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_102),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_148),
.B1(n_125),
.B2(n_149),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_104),
.B(n_97),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_102),
.B1(n_17),
.B2(n_23),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_192),
.B1(n_193),
.B2(n_160),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_138),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_201),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_155),
.B1(n_174),
.B2(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_197),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_196),
.B(n_203),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_126),
.C(n_127),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_150),
.B1(n_133),
.B2(n_142),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_156),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_179),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_150),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_33),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_177),
.C(n_176),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_141),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_204),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_134),
.B(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_97),
.C(n_134),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_93),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_93),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_209),
.B1(n_181),
.B2(n_192),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_186),
.B1(n_184),
.B2(n_29),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_152),
.B1(n_161),
.B2(n_167),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_171),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_214),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_180),
.Y(n_214)
);

NAND2x1_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_172),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_203),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_183),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_221),
.B(n_227),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_156),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_229),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_17),
.B1(n_28),
.B2(n_22),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_28),
.B1(n_22),
.B2(n_97),
.Y(n_223)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_183),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_184),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_198),
.B1(n_205),
.B2(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_224),
.B(n_227),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_189),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_244),
.B(n_254),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_234),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_182),
.C(n_201),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_238),
.C(n_242),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_236),
.A2(n_237),
.B1(n_247),
.B2(n_0),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_198),
.B(n_186),
.C(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_204),
.C(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_230),
.B1(n_220),
.B2(n_3),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_33),
.C(n_29),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_33),
.C(n_29),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_226),
.C(n_225),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_10),
.B(n_16),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_28),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_263),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_229),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_262),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_219),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_208),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_265),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_252),
.C(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_243),
.C(n_233),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_225),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_29),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_270),
.A2(n_272),
.B1(n_247),
.B2(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_230),
.B1(n_220),
.B2(n_12),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_245),
.B1(n_237),
.B2(n_234),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_259),
.C(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_236),
.C(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_281),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_248),
.C(n_237),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_244),
.B(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_248),
.B1(n_12),
.B2(n_13),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_261),
.B1(n_14),
.B2(n_15),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_262),
.B(n_8),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_263),
.C(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_2),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_290),
.A2(n_287),
.B1(n_9),
.B2(n_14),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_260),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_292),
.B(n_298),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_264),
.B(n_4),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_284),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_299),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_8),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_27),
.C(n_15),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_9),
.C(n_14),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_277),
.B1(n_278),
.B2(n_275),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_274),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_285),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_307),
.A2(n_297),
.B(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_296),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_285),
.C(n_9),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_319),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_4),
.B(n_5),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_317),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_302),
.C(n_5),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_4),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_320),
.B(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_321),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_325),
.B(n_6),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_5),
.B(n_6),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_7),
.B(n_317),
.Y(n_331)
);


endmodule