module real_aes_3810_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1106;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_1123;
wire n_549;
wire n_571;
wire n_491;
wire n_694;
wire n_894;
wire n_1034;
wire n_923;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1053;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_726;
wire n_369;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_725;
wire n_455;
wire n_504;
wire n_973;
wire n_1081;
wire n_671;
wire n_1084;
wire n_960;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_1031;
wire n_1103;
wire n_880;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1014;
wire n_1028;
wire n_366;
wire n_346;
wire n_1083;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_1043;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_1102;
wire n_601;
wire n_463;
wire n_661;
wire n_396;
wire n_804;
wire n_1076;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_1104;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_0), .A2(n_176), .B1(n_480), .B2(n_482), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_1), .A2(n_130), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_2), .A2(n_219), .B1(n_391), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_3), .A2(n_143), .B1(n_527), .B2(n_664), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_4), .A2(n_266), .B1(n_587), .B2(n_588), .Y(n_1116) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_5), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_6), .A2(n_227), .B1(n_818), .B2(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g598 ( .A(n_7), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_8), .A2(n_280), .B1(n_558), .B2(n_664), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_9), .A2(n_253), .B1(n_419), .B2(n_573), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_10), .A2(n_21), .B1(n_376), .B2(n_456), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_11), .B(n_339), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_12), .A2(n_283), .B1(n_480), .B2(n_527), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_13), .A2(n_209), .B1(n_505), .B2(n_506), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_14), .A2(n_150), .B1(n_391), .B2(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_15), .B(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_16), .A2(n_181), .B1(n_508), .B2(n_509), .Y(n_739) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_17), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_18), .A2(n_57), .B1(n_471), .B2(n_545), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_19), .A2(n_128), .B1(n_451), .B2(n_523), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_20), .A2(n_32), .B1(n_332), .B2(n_358), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_22), .A2(n_129), .B1(n_372), .B2(n_484), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_23), .A2(n_191), .B1(n_408), .B2(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g611 ( .A(n_24), .Y(n_611) );
INVx1_ASAP7_75t_L g463 ( .A(n_25), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_26), .A2(n_533), .B(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g536 ( .A(n_27), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_28), .A2(n_81), .B1(n_509), .B2(n_736), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_29), .A2(n_180), .B1(n_371), .B2(n_376), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_30), .A2(n_308), .B1(n_508), .B2(n_509), .Y(n_507) );
XOR2x2_ASAP7_75t_L g728 ( .A(n_31), .B(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_31), .A2(n_142), .B1(n_870), .B2(n_878), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_33), .A2(n_38), .B1(n_371), .B2(n_376), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_34), .A2(n_126), .B1(n_560), .B2(n_664), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_35), .A2(n_89), .B1(n_419), .B2(n_757), .Y(n_784) );
INVx1_ASAP7_75t_L g567 ( .A(n_36), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_37), .A2(n_110), .B1(n_419), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_39), .A2(n_119), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_40), .A2(n_145), .B1(n_333), .B2(n_372), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_41), .A2(n_157), .B1(n_529), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_42), .A2(n_86), .B1(n_505), .B2(n_506), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_43), .A2(n_167), .B1(n_391), .B2(n_394), .Y(n_452) );
OA22x2_ASAP7_75t_L g345 ( .A1(n_44), .A2(n_141), .B1(n_339), .B2(n_343), .Y(n_345) );
INVx1_ASAP7_75t_L g366 ( .A(n_44), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_45), .A2(n_259), .B1(n_359), .B2(n_523), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_46), .A2(n_52), .B1(n_428), .B2(n_438), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_47), .A2(n_50), .B1(n_505), .B2(n_506), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_48), .A2(n_248), .B1(n_480), .B2(n_482), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_49), .A2(n_296), .B1(n_682), .B2(n_818), .Y(n_817) );
XNOR2x2_ASAP7_75t_L g640 ( .A(n_51), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g856 ( .A(n_51), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_53), .A2(n_215), .B1(n_499), .B2(n_501), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_54), .A2(n_133), .B1(n_844), .B2(n_847), .Y(n_843) );
INVx1_ASAP7_75t_L g675 ( .A(n_55), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_56), .A2(n_85), .B1(n_482), .B2(n_557), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_58), .A2(n_163), .B1(n_603), .B2(n_631), .C(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g858 ( .A(n_59), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_60), .B(n_158), .Y(n_322) );
INVx1_ASAP7_75t_L g342 ( .A(n_60), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_60), .A2(n_141), .B(n_368), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_61), .A2(n_473), .B(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_62), .A2(n_131), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_63), .A2(n_250), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_64), .A2(n_230), .B1(n_391), .B2(n_394), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_65), .A2(n_122), .B1(n_451), .B2(n_621), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_66), .A2(n_97), .B1(n_868), .B2(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_67), .A2(n_161), .B1(n_621), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_68), .A2(n_185), .B1(n_451), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_69), .A2(n_132), .B1(n_633), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_70), .A2(n_277), .B1(n_469), .B2(n_471), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_71), .A2(n_104), .B1(n_371), .B2(n_376), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_72), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_73), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g839 ( .A(n_74), .Y(n_839) );
AND2x4_ASAP7_75t_L g842 ( .A(n_74), .B(n_228), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_75), .A2(n_203), .B1(n_451), .B2(n_527), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_76), .A2(n_265), .B1(n_841), .B2(n_868), .Y(n_895) );
INVx1_ASAP7_75t_L g1076 ( .A(n_76), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_76), .A2(n_1104), .B1(n_1106), .B2(n_1124), .Y(n_1103) );
INVx1_ASAP7_75t_L g822 ( .A(n_77), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_78), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_79), .A2(n_80), .B1(n_454), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_82), .A2(n_173), .B1(n_498), .B2(n_499), .Y(n_497) );
AO22x2_ASAP7_75t_L g867 ( .A1(n_83), .A2(n_247), .B1(n_841), .B2(n_868), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_84), .A2(n_88), .B1(n_414), .B2(n_490), .C(n_820), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_87), .A2(n_565), .B(n_566), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g670 ( .A(n_90), .B(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_90), .A2(n_115), .B1(n_847), .B2(n_888), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_91), .A2(n_490), .B(n_493), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_92), .A2(n_267), .B1(n_565), .B2(n_587), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_93), .B(n_755), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_94), .A2(n_116), .B1(n_870), .B2(n_878), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_95), .A2(n_460), .B(n_462), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_96), .A2(n_134), .B1(n_667), .B2(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g821 ( .A(n_98), .Y(n_821) );
AND2x4_ASAP7_75t_L g840 ( .A(n_99), .B(n_318), .Y(n_840) );
INVx1_ASAP7_75t_L g846 ( .A(n_99), .Y(n_846) );
INVx1_ASAP7_75t_SL g871 ( .A(n_99), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_100), .A2(n_220), .B1(n_419), .B2(n_498), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_101), .A2(n_243), .B1(n_522), .B2(n_524), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_102), .A2(n_169), .B1(n_654), .B2(n_655), .Y(n_653) );
XNOR2x2_ASAP7_75t_SL g578 ( .A(n_103), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g1119 ( .A(n_105), .Y(n_1119) );
INVx1_ASAP7_75t_L g789 ( .A(n_106), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_107), .A2(n_223), .B1(n_560), .B2(n_667), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_108), .A2(n_125), .B1(n_841), .B2(n_868), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_109), .A2(n_286), .B1(n_380), .B2(n_529), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_111), .A2(n_302), .B1(n_602), .B2(n_603), .C(n_605), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_112), .A2(n_310), .B1(n_844), .B2(n_868), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_113), .A2(n_127), .B1(n_482), .B2(n_664), .Y(n_663) );
XNOR2x1_ASAP7_75t_L g476 ( .A(n_114), .B(n_477), .Y(n_476) );
OAI22x1_ASAP7_75t_L g701 ( .A1(n_116), .A2(n_702), .B1(n_725), .B2(n_726), .Y(n_701) );
NAND3xp33_ASAP7_75t_SL g725 ( .A(n_116), .B(n_714), .C(n_722), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g1106 ( .A(n_117), .B(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g486 ( .A(n_118), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_120), .A2(n_156), .B1(n_735), .B2(n_736), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_121), .A2(n_301), .B1(n_505), .B2(n_506), .Y(n_1113) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_123), .A2(n_473), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g592 ( .A(n_124), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_135), .B(n_460), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_136), .A2(n_263), .B1(n_529), .B2(n_562), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_137), .A2(n_252), .B1(n_662), .B2(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g474 ( .A(n_138), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_139), .A2(n_289), .B1(n_508), .B2(n_509), .Y(n_1114) );
INVx1_ASAP7_75t_L g357 ( .A(n_140), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_140), .B(n_188), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_140), .B(n_364), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_141), .B(n_237), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_144), .A2(n_257), .B1(n_359), .B2(n_583), .Y(n_1089) );
INVx1_ASAP7_75t_L g627 ( .A(n_146), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_147), .A2(n_231), .B1(n_572), .B2(n_573), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_148), .A2(n_159), .B1(n_414), .B2(n_690), .C(n_691), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_149), .A2(n_258), .B1(n_562), .B2(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_151), .A2(n_155), .B1(n_573), .B2(n_783), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_152), .A2(n_205), .B1(n_562), .B2(n_662), .Y(n_813) );
INVx1_ASAP7_75t_L g760 ( .A(n_153), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_154), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_158), .B(n_350), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_160), .A2(n_184), .B1(n_372), .B2(n_560), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_162), .A2(n_309), .B1(n_562), .B2(n_662), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_164), .A2(n_311), .B1(n_454), .B2(n_662), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_165), .A2(n_197), .B1(n_333), .B2(n_451), .Y(n_665) );
INVx1_ASAP7_75t_L g495 ( .A(n_166), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_168), .A2(n_211), .B1(n_545), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_170), .A2(n_251), .B1(n_667), .B2(n_668), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_171), .B(n_595), .Y(n_594) );
AOI21xp33_ASAP7_75t_SL g1082 ( .A1(n_172), .A2(n_757), .B(n_1083), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_174), .A2(n_291), .B1(n_573), .B2(n_753), .Y(n_752) );
INVxp33_ASAP7_75t_SL g863 ( .A(n_175), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_177), .A2(n_771), .B1(n_772), .B2(n_790), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_177), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_178), .A2(n_295), .B1(n_835), .B2(n_841), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g1085 ( .A(n_179), .B(n_1086), .Y(n_1085) );
XNOR2x1_ASAP7_75t_L g552 ( .A(n_182), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_183), .A2(n_293), .B1(n_419), .B2(n_659), .Y(n_1087) );
INVx1_ASAP7_75t_L g692 ( .A(n_186), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_187), .A2(n_288), .B1(n_372), .B2(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g340 ( .A(n_188), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_189), .A2(n_213), .B1(n_456), .B2(n_457), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_190), .B(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_192), .A2(n_304), .B1(n_380), .B2(n_386), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_193), .A2(n_212), .B1(n_386), .B2(n_454), .Y(n_453) );
XNOR2x1_ASAP7_75t_L g791 ( .A(n_194), .B(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_195), .A2(n_285), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g1084 ( .A(n_196), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_198), .A2(n_234), .B1(n_540), .B2(n_542), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g1111 ( .A1(n_199), .A2(n_204), .B1(n_542), .B2(n_659), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_200), .B(n_461), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_201), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_202), .A2(n_271), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_206), .A2(n_221), .B1(n_735), .B2(n_736), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_207), .A2(n_260), .B1(n_584), .B2(n_621), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_208), .A2(n_244), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_210), .A2(n_290), .B1(n_844), .B2(n_872), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_214), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_216), .A2(n_240), .B1(n_499), .B2(n_501), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_217), .A2(n_241), .B1(n_372), .B2(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_218), .A2(n_294), .B1(n_583), .B2(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_222), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_224), .A2(n_254), .B1(n_588), .B2(n_735), .Y(n_801) );
INVx1_ASAP7_75t_L g600 ( .A(n_225), .Y(n_600) );
AO22x1_ASAP7_75t_L g869 ( .A1(n_226), .A2(n_233), .B1(n_870), .B2(n_872), .Y(n_869) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_228), .Y(n_323) );
AND2x4_ASAP7_75t_L g838 ( .A(n_228), .B(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_229), .B(n_690), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_232), .A2(n_305), .B1(n_418), .B2(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g677 ( .A(n_235), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_236), .A2(n_273), .B1(n_502), .B2(n_565), .Y(n_740) );
INVx1_ASAP7_75t_L g355 ( .A(n_237), .Y(n_355) );
INVxp67_ASAP7_75t_L g437 ( .A(n_237), .Y(n_437) );
INVx1_ASAP7_75t_L g732 ( .A(n_238), .Y(n_732) );
INVx1_ASAP7_75t_L g1123 ( .A(n_239), .Y(n_1123) );
AOI22xp5_ASAP7_75t_SL g722 ( .A1(n_242), .A2(n_281), .B1(n_533), .B2(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g318 ( .A(n_245), .Y(n_318) );
INVxp33_ASAP7_75t_SL g966 ( .A(n_246), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_249), .A2(n_644), .B(n_647), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_255), .A2(n_256), .B1(n_502), .B2(n_508), .Y(n_795) );
AO221x2_ASAP7_75t_L g962 ( .A1(n_261), .A2(n_262), .B1(n_835), .B2(n_963), .C(n_964), .Y(n_962) );
INVx1_ASAP7_75t_L g606 ( .A(n_264), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g797 ( .A1(n_268), .A2(n_604), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_269), .Y(n_799) );
INVx1_ASAP7_75t_L g679 ( .A(n_270), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_272), .A2(n_300), .B1(n_380), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_274), .A2(n_287), .B1(n_419), .B2(n_488), .Y(n_568) );
INVx1_ASAP7_75t_L g749 ( .A(n_275), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_276), .A2(n_519), .B(n_546), .Y(n_518) );
INVx1_ASAP7_75t_L g548 ( .A(n_276), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_278), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_279), .B(n_651), .Y(n_650) );
XNOR2x2_ASAP7_75t_L g329 ( .A(n_282), .B(n_330), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_284), .A2(n_298), .B1(n_391), .B2(n_394), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_292), .A2(n_306), .B1(n_333), .B2(n_451), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_297), .A2(n_492), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g648 ( .A(n_299), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_303), .Y(n_399) );
AOI21xp33_ASAP7_75t_SL g787 ( .A1(n_307), .A2(n_658), .B(n_788), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_324), .B(n_827), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_316), .B(n_1101), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_316), .B(n_1102), .Y(n_1105) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OA21x2_ASAP7_75t_L g1125 ( .A1(n_317), .A2(n_871), .B(n_1126), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g845 ( .A(n_318), .B(n_846), .Y(n_845) );
AND3x4_ASAP7_75t_L g870 ( .A(n_318), .B(n_838), .C(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g1101 ( .A(n_319), .B(n_1102), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_320), .A2(n_442), .B(n_443), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g1102 ( .A(n_323), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_696), .B2(n_697), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
XNOR2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_511), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OA22x2_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_445), .B1(n_446), .B2(n_510), .Y(n_328) );
INVx3_ASAP7_75t_L g510 ( .A(n_329), .Y(n_510) );
NAND3xp33_ASAP7_75t_SL g330 ( .A(n_331), .B(n_369), .C(n_397), .Y(n_330) );
BUFx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_334), .Y(n_523) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_334), .Y(n_583) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_334), .Y(n_621) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_346), .Y(n_334) );
AND2x4_ASAP7_75t_L g373 ( .A(n_335), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g383 ( .A(n_335), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g387 ( .A(n_335), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g505 ( .A(n_335), .B(n_384), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_335), .B(n_388), .Y(n_506) );
AND2x4_ASAP7_75t_L g508 ( .A(n_335), .B(n_396), .Y(n_508) );
AND2x4_ASAP7_75t_L g735 ( .A(n_335), .B(n_374), .Y(n_735) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_344), .Y(n_335) );
AND2x2_ASAP7_75t_L g404 ( .A(n_336), .B(n_345), .Y(n_404) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g393 ( .A(n_337), .B(n_345), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
NAND2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g343 ( .A(n_339), .Y(n_343) );
INVx3_ASAP7_75t_L g350 ( .A(n_339), .Y(n_350) );
NAND2xp33_ASAP7_75t_L g356 ( .A(n_339), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_339), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_340), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_342), .A2(n_368), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g435 ( .A(n_345), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g361 ( .A(n_346), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g509 ( .A(n_346), .B(n_362), .Y(n_509) );
AND2x4_ASAP7_75t_L g588 ( .A(n_346), .B(n_393), .Y(n_588) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g396 ( .A(n_347), .Y(n_396) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_352), .Y(n_347) );
AND2x4_ASAP7_75t_L g374 ( .A(n_348), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g384 ( .A(n_348), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g389 ( .A(n_348), .Y(n_389) );
AND2x2_ASAP7_75t_L g431 ( .A(n_348), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_350), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g364 ( .A(n_350), .Y(n_364) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_351), .B(n_363), .C(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx5_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g524 ( .A(n_360), .Y(n_524) );
INVx3_ASAP7_75t_L g584 ( .A(n_360), .Y(n_584) );
INVx2_ASAP7_75t_L g763 ( .A(n_360), .Y(n_763) );
INVx6_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx12f_ASAP7_75t_L g451 ( .A(n_361), .Y(n_451) );
AND2x4_ASAP7_75t_L g378 ( .A(n_362), .B(n_374), .Y(n_378) );
AND2x4_ASAP7_75t_L g420 ( .A(n_362), .B(n_388), .Y(n_420) );
AND2x4_ASAP7_75t_L g502 ( .A(n_362), .B(n_388), .Y(n_502) );
AND2x4_ASAP7_75t_L g736 ( .A(n_362), .B(n_374), .Y(n_736) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_367), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND3x1_ASAP7_75t_L g369 ( .A(n_370), .B(n_379), .C(n_390), .Y(n_369) );
BUFx12f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx12f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_373), .Y(n_456) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_373), .Y(n_667) );
AND2x2_ASAP7_75t_L g392 ( .A(n_374), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g481 ( .A(n_374), .B(n_393), .Y(n_481) );
AND2x4_ASAP7_75t_L g587 ( .A(n_374), .B(n_393), .Y(n_587) );
INVx4_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g457 ( .A(n_377), .Y(n_457) );
INVx1_ASAP7_75t_L g484 ( .A(n_377), .Y(n_484) );
INVx2_ASAP7_75t_L g560 ( .A(n_377), .Y(n_560) );
INVx4_ASAP7_75t_L g668 ( .A(n_377), .Y(n_668) );
INVx2_ASAP7_75t_L g780 ( .A(n_377), .Y(n_780) );
INVx8_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx4f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g775 ( .A(n_382), .Y(n_775) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_383), .Y(n_454) );
BUFx12f_ASAP7_75t_L g562 ( .A(n_383), .Y(n_562) );
AND2x4_ASAP7_75t_L g403 ( .A(n_384), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g410 ( .A(n_384), .B(n_393), .Y(n_410) );
AND2x4_ASAP7_75t_L g501 ( .A(n_384), .B(n_393), .Y(n_501) );
AND2x4_ASAP7_75t_L g565 ( .A(n_384), .B(n_404), .Y(n_565) );
AND2x4_ASAP7_75t_L g388 ( .A(n_385), .B(n_389), .Y(n_388) );
BUFx5_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g529 ( .A(n_387), .Y(n_529) );
INVx1_ASAP7_75t_L g617 ( .A(n_387), .Y(n_617) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_387), .Y(n_662) );
AND2x4_ASAP7_75t_L g415 ( .A(n_388), .B(n_404), .Y(n_415) );
AND2x2_ASAP7_75t_L g426 ( .A(n_388), .B(n_393), .Y(n_426) );
AND2x2_ASAP7_75t_L g492 ( .A(n_388), .B(n_393), .Y(n_492) );
AND2x2_ASAP7_75t_L g604 ( .A(n_388), .B(n_404), .Y(n_604) );
BUFx8_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_392), .Y(n_664) );
AND2x4_ASAP7_75t_L g395 ( .A(n_393), .B(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_395), .Y(n_482) );
BUFx12f_ASAP7_75t_L g527 ( .A(n_395), .Y(n_527) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_395), .Y(n_558) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_395), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_411), .C(n_421), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_405), .B2(n_406), .Y(n_398) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g658 ( .A(n_402), .Y(n_658) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_403), .Y(n_473) );
BUFx3_ASAP7_75t_L g498 ( .A(n_403), .Y(n_498) );
BUFx3_ASAP7_75t_L g818 ( .A(n_403), .Y(n_818) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_409), .Y(n_541) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g573 ( .A(n_410), .Y(n_573) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_410), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_416), .B2(n_417), .Y(n_411) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
BUFx8_ASAP7_75t_SL g654 ( .A(n_415), .Y(n_654) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_415), .Y(n_757) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g676 ( .A(n_419), .Y(n_676) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_420), .Y(n_471) );
INVx3_ASAP7_75t_L g656 ( .A(n_420), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx3_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g570 ( .A(n_425), .Y(n_570) );
INVx2_ASAP7_75t_L g631 ( .A(n_425), .Y(n_631) );
INVx2_ASAP7_75t_L g755 ( .A(n_425), .Y(n_755) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g461 ( .A(n_426), .Y(n_461) );
INVx2_ASAP7_75t_L g646 ( .A(n_426), .Y(n_646) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_429), .A2(n_463), .B(n_464), .Y(n_462) );
INVx3_ASAP7_75t_L g542 ( .A(n_429), .Y(n_542) );
INVx2_ASAP7_75t_L g633 ( .A(n_429), .Y(n_633) );
INVx2_ASAP7_75t_L g753 ( .A(n_429), .Y(n_753) );
INVx4_ASAP7_75t_L g783 ( .A(n_429), .Y(n_783) );
INVx5_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g572 ( .A(n_430), .Y(n_572) );
BUFx4f_ASAP7_75t_L g682 ( .A(n_430), .Y(n_682) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_430), .Y(n_1081) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_435), .Y(n_430) );
AND2x2_ASAP7_75t_L g499 ( .A(n_431), .B(n_435), .Y(n_499) );
AND2x4_ASAP7_75t_L g595 ( .A(n_431), .B(n_435), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g442 ( .A(n_433), .Y(n_442) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_439), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_439), .B(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_439), .B(n_1123), .Y(n_1122) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx4_ASAP7_75t_L g652 ( .A(n_440), .Y(n_652) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_441), .Y(n_467) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_475), .Y(n_446) );
XNOR2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_474), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_458), .Y(n_448) );
NAND4xp25_ASAP7_75t_SL g449 ( .A(n_450), .B(n_452), .C(n_453), .D(n_455), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_468), .C(n_472), .Y(n_458) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_466), .B(n_760), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g1083 ( .A(n_466), .B(n_1084), .Y(n_1083) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
INVx2_ASAP7_75t_L g538 ( .A(n_467), .Y(n_538) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g545 ( .A(n_470), .Y(n_545) );
INVx4_ASAP7_75t_L g711 ( .A(n_471), .Y(n_711) );
INVx4_ASAP7_75t_L g680 ( .A(n_473), .Y(n_680) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND4xp75_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .C(n_496), .D(n_503), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx4f_ASAP7_75t_L g557 ( .A(n_481), .Y(n_557) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_489), .Y(n_485) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_492), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_494), .B(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_494), .B(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_494), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .Y(n_496) );
INVx2_ASAP7_75t_L g534 ( .A(n_498), .Y(n_534) );
INVx1_ASAP7_75t_L g597 ( .A(n_501), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_502), .Y(n_599) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_575), .B2(n_695), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OA22x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_550), .B2(n_574), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
INVxp67_ASAP7_75t_L g549 ( .A(n_520), .Y(n_549) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .C(n_528), .D(n_530), .Y(n_520) );
BUFx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_531), .B(n_548), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .C(n_543), .D(n_544), .Y(n_531) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g634 ( .A(n_541), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g574 ( .A(n_552), .Y(n_574) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_563), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_559), .D(n_561), .Y(n_554) );
NAND4xp25_ASAP7_75t_SL g563 ( .A(n_564), .B(n_568), .C(n_569), .D(n_571), .Y(n_563) );
INVx2_ASAP7_75t_L g593 ( .A(n_565), .Y(n_593) );
INVx2_ASAP7_75t_L g724 ( .A(n_573), .Y(n_724) );
INVx1_ASAP7_75t_L g695 ( .A(n_575), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_637), .B2(n_638), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AO22x2_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_607), .B1(n_635), .B2(n_636), .Y(n_577) );
INVx2_ASAP7_75t_L g635 ( .A(n_578), .Y(n_635) );
NAND4xp75_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .C(n_590), .D(n_601), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_596), .Y(n_590) );
OAI21xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_594), .Y(n_591) );
INVx4_ASAP7_75t_L g649 ( .A(n_595), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_596) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g636 ( .A(n_609), .Y(n_636) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
XNOR2x1_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_613), .B(n_622), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .C(n_619), .D(n_620), .Y(n_613) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g720 ( .A(n_616), .Y(n_720) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_629), .C(n_632), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .Y(n_624) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OA22x2_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_669), .B2(n_694), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_660), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_653), .C(n_657), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
INVx1_ASAP7_75t_L g1086 ( .A(n_645), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g708 ( .A(n_646), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_650), .Y(n_647) );
INVx2_ASAP7_75t_L g693 ( .A(n_651), .Y(n_693) );
INVx4_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g713 ( .A(n_652), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_652), .B(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_652), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1120 ( .A(n_654), .Y(n_1120) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g674 ( .A(n_659), .Y(n_674) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .C(n_665), .D(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g694 ( .A(n_669), .Y(n_694) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND4xp75_ASAP7_75t_L g671 ( .A(n_672), .B(n_683), .C(n_686), .D(n_689), .Y(n_671) );
NOR2xp67_ASAP7_75t_L g672 ( .A(n_673), .B(n_678), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B(n_681), .Y(n_678) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_744), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AO22x2_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_727), .B2(n_743), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_714), .C(n_722), .Y(n_703) );
INVx1_ASAP7_75t_L g726 ( .A(n_704), .Y(n_726) );
AND3x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_709), .C(n_712), .Y(n_704) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND4x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .C(n_718), .D(n_721), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_728), .Y(n_743) );
NAND3x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .C(n_738), .Y(n_729) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
AND4x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .C(n_741), .D(n_742), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_767), .B1(n_825), .B2(n_826), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_746), .Y(n_826) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NOR2xp67_ASAP7_75t_L g750 ( .A(n_751), .B(n_761), .Y(n_750) );
NAND4xp25_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .C(n_756), .D(n_758), .Y(n_751) );
NAND4xp25_ASAP7_75t_SL g761 ( .A(n_762), .B(n_764), .C(n_765), .D(n_766), .Y(n_761) );
INVx1_ASAP7_75t_L g825 ( .A(n_767), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B1(n_805), .B2(n_823), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
XOR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_791), .Y(n_769) );
INVx1_ASAP7_75t_L g790 ( .A(n_772), .Y(n_790) );
NAND4xp75_ASAP7_75t_L g772 ( .A(n_773), .B(n_777), .C(n_781), .D(n_785), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
OR2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_800), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .C(n_796), .D(n_797), .Y(n_793) );
NAND4xp25_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .C(n_803), .D(n_804), .Y(n_800) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx3_ASAP7_75t_L g824 ( .A(n_807), .Y(n_824) );
XNOR2x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_822), .Y(n_807) );
NAND4xp75_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .C(n_815), .D(n_819), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_1068), .B1(n_1070), .B2(n_1099), .C(n_1103), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_974), .B(n_1022), .Y(n_828) );
OAI211xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_848), .B(n_907), .C(n_941), .Y(n_829) );
CKINVDCx14_ASAP7_75t_R g985 ( .A(n_830), .Y(n_985) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_830), .A2(n_938), .B1(n_1009), .B2(n_1011), .C(n_1018), .Y(n_1008) );
O2A1O1Ixp33_ASAP7_75t_L g1023 ( .A1(n_830), .A2(n_1024), .B(n_1027), .C(n_1031), .Y(n_1023) );
OAI222xp33_ASAP7_75t_L g1040 ( .A1(n_830), .A2(n_958), .B1(n_993), .B2(n_1041), .C1(n_1043), .C2(n_1046), .Y(n_1040) );
INVx5_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_831), .B(n_920), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_831), .B(n_957), .Y(n_956) );
INVx3_ASAP7_75t_L g1050 ( .A(n_831), .Y(n_1050) );
INVx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
AND2x2_ASAP7_75t_L g908 ( .A(n_832), .B(n_909), .Y(n_908) );
AND2x2_ASAP7_75t_L g996 ( .A(n_832), .B(n_873), .Y(n_996) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_832), .B(n_924), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_832), .B(n_865), .Y(n_1065) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_832), .B(n_866), .Y(n_1067) );
INVx3_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g934 ( .A(n_833), .B(n_924), .Y(n_934) );
OR2x2_ASAP7_75t_L g939 ( .A(n_833), .B(n_940), .Y(n_939) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_833), .B(n_973), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_843), .Y(n_833) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
AND2x4_ASAP7_75t_L g837 ( .A(n_838), .B(n_840), .Y(n_837) );
AND2x4_ASAP7_75t_L g844 ( .A(n_838), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_838), .B(n_840), .Y(n_862) );
AND2x4_ASAP7_75t_L g868 ( .A(n_838), .B(n_840), .Y(n_868) );
AND2x4_ASAP7_75t_L g841 ( .A(n_840), .B(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g876 ( .A(n_840), .B(n_842), .Y(n_876) );
AND2x2_ASAP7_75t_L g888 ( .A(n_840), .B(n_842), .Y(n_888) );
INVx2_ASAP7_75t_L g857 ( .A(n_841), .Y(n_857) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_841), .Y(n_1069) );
AND2x4_ASAP7_75t_L g847 ( .A(n_842), .B(n_845), .Y(n_847) );
AND2x2_ASAP7_75t_L g872 ( .A(n_842), .B(n_845), .Y(n_872) );
AND2x2_ASAP7_75t_L g878 ( .A(n_842), .B(n_845), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g1126 ( .A(n_842), .Y(n_1126) );
INVx3_ASAP7_75t_L g860 ( .A(n_844), .Y(n_860) );
INVx3_ASAP7_75t_L g855 ( .A(n_847), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_865), .B1(n_879), .B2(n_890), .C(n_897), .Y(n_848) );
INVxp67_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_864), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_851), .B(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_851), .B(n_916), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_851), .B(n_921), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_851), .B(n_929), .Y(n_1025) );
INVx1_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
AND2x2_ASAP7_75t_L g915 ( .A(n_852), .B(n_916), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_852), .B(n_874), .Y(n_928) );
AND2x2_ASAP7_75t_L g971 ( .A(n_852), .B(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_852), .B(n_886), .Y(n_1060) );
INVx3_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g903 ( .A(n_853), .Y(n_903) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_853), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_853), .B(n_896), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_853), .B(n_874), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_853), .B(n_957), .Y(n_1007) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_853), .B(n_866), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_853), .B(n_900), .Y(n_1052) );
OR2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_859), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_855), .A2(n_857), .B1(n_965), .B2(n_966), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_859) );
INVx1_ASAP7_75t_L g963 ( .A(n_860), .Y(n_963) );
INVx1_ASAP7_75t_L g1016 ( .A(n_864), .Y(n_1016) );
AND2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_873), .Y(n_864) );
OAI211xp5_ASAP7_75t_SL g913 ( .A1(n_865), .A2(n_914), .B(n_917), .C(n_931), .Y(n_913) );
INVx1_ASAP7_75t_L g1002 ( .A(n_865), .Y(n_1002) );
CKINVDCx6p67_ASAP7_75t_R g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g920 ( .A(n_866), .B(n_874), .Y(n_920) );
INVx1_ASAP7_75t_L g925 ( .A(n_866), .Y(n_925) );
AND2x2_ASAP7_75t_L g957 ( .A(n_866), .B(n_900), .Y(n_957) );
OR2x2_ASAP7_75t_L g973 ( .A(n_866), .B(n_874), .Y(n_973) );
OAI322xp33_ASAP7_75t_L g976 ( .A1(n_866), .A2(n_950), .A3(n_960), .B1(n_977), .B2(n_978), .C1(n_979), .C2(n_981), .Y(n_976) );
OR2x6_ASAP7_75t_L g866 ( .A(n_867), .B(n_869), .Y(n_866) );
BUFx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_874), .Y(n_900) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_874), .Y(n_1028) );
AND2x4_ASAP7_75t_L g874 ( .A(n_875), .B(n_877), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_879), .B(n_948), .Y(n_947) );
CKINVDCx16_ASAP7_75t_R g978 ( .A(n_879), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_879), .B(n_1006), .Y(n_1005) );
AND2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_884), .Y(n_879) );
AND2x2_ASAP7_75t_L g916 ( .A(n_880), .B(n_893), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_880), .B(n_896), .Y(n_922) );
OR2x2_ASAP7_75t_L g930 ( .A(n_880), .B(n_896), .Y(n_930) );
OR2x2_ASAP7_75t_L g951 ( .A(n_880), .B(n_893), .Y(n_951) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_880), .B(n_884), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
OR2x2_ASAP7_75t_L g906 ( .A(n_881), .B(n_893), .Y(n_906) );
AND2x2_ASAP7_75t_L g933 ( .A(n_881), .B(n_893), .Y(n_933) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_884), .B(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g932 ( .A(n_884), .B(n_933), .Y(n_932) );
AND2x2_ASAP7_75t_L g937 ( .A(n_884), .B(n_916), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_884), .B(n_954), .Y(n_988) );
O2A1O1Ixp33_ASAP7_75t_SL g1031 ( .A1(n_884), .A2(n_1032), .B(n_1035), .C(n_1037), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_884), .B(n_1003), .Y(n_1036) );
AND3x1_ASAP7_75t_L g1042 ( .A(n_884), .B(n_909), .C(n_915), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_884), .B(n_893), .Y(n_1045) );
INVx3_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx3_ASAP7_75t_L g896 ( .A(n_886), .Y(n_896) );
OR2x2_ASAP7_75t_L g983 ( .A(n_886), .B(n_893), .Y(n_983) );
AND2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AOI31xp33_ASAP7_75t_L g1024 ( .A1(n_891), .A2(n_1016), .A3(n_1025), .B(n_1026), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1017 ( .A(n_892), .Y(n_1017) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
OR2x2_ASAP7_75t_L g905 ( .A(n_896), .B(n_906), .Y(n_905) );
AND2x2_ASAP7_75t_L g911 ( .A(n_896), .B(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_896), .B(n_950), .Y(n_949) );
AND2x2_ASAP7_75t_L g959 ( .A(n_896), .B(n_933), .Y(n_959) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_896), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_896), .B(n_951), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_901), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_898), .B(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g909 ( .A(n_899), .Y(n_909) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
AND2x2_ASAP7_75t_L g910 ( .A(n_902), .B(n_911), .Y(n_910) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_902), .B(n_932), .C(n_934), .Y(n_931) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_903), .B(n_951), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_903), .B(n_983), .Y(n_982) );
O2A1O1Ixp33_ASAP7_75t_L g1018 ( .A1(n_903), .A2(n_978), .B(n_1019), .C(n_1021), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_903), .B(n_933), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_903), .B(n_959), .Y(n_1063) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g912 ( .A(n_906), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_906), .B(n_1034), .Y(n_1033) );
AOI211xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_910), .B(n_913), .C(n_935), .Y(n_907) );
INVx1_ASAP7_75t_L g1021 ( .A(n_908), .Y(n_1021) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_909), .A2(n_1000), .B1(n_1001), .B2(n_1003), .C(n_1004), .Y(n_999) );
INVx1_ASAP7_75t_L g994 ( .A(n_911), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_914), .Y(n_984) );
AND2x2_ASAP7_75t_L g969 ( .A(n_916), .B(n_970), .Y(n_969) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_916), .B(n_1030), .Y(n_1029) );
AOI21xp33_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_921), .B(n_923), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx2_ASAP7_75t_L g940 ( .A(n_920), .Y(n_940) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_922), .B(n_928), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_926), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_924), .B(n_980), .Y(n_993) );
AOI211xp5_ASAP7_75t_L g1038 ( .A1(n_924), .A2(n_1039), .B(n_1040), .C(n_1047), .Y(n_1038) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AOI21xp33_ASAP7_75t_SL g1066 ( .A1(n_926), .A2(n_997), .B(n_1067), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_929), .Y(n_926) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_927), .B(n_937), .Y(n_1039) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g1055 ( .A(n_932), .Y(n_1055) );
INVx1_ASAP7_75t_L g1034 ( .A(n_933), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_934), .B(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g1046 ( .A(n_934), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g935 ( .A(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_937), .B(n_972), .Y(n_991) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
AOI211xp5_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_946), .B(n_952), .C(n_967), .Y(n_941) );
INVxp67_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVxp67_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g968 ( .A1(n_950), .A2(n_969), .B(n_971), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_950), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .B1(n_958), .B2(n_960), .C(n_961), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g960 ( .A(n_957), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_958), .B(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NOR3xp33_ASAP7_75t_L g989 ( .A(n_961), .B(n_990), .C(n_992), .Y(n_989) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g1026 ( .A(n_969), .Y(n_1026) );
INVx2_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
NAND5xp2_ASAP7_75t_SL g974 ( .A(n_975), .B(n_986), .C(n_989), .D(n_999), .E(n_1008), .Y(n_974) );
OAI21xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_984), .B(n_985), .Y(n_975) );
INVx1_ASAP7_75t_L g1030 ( .A(n_977), .Y(n_1030) );
INVxp67_ASAP7_75t_SL g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVxp67_ASAP7_75t_SL g986 ( .A(n_987), .Y(n_986) );
INVxp67_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_994), .B1(n_995), .B2(n_997), .Y(n_992) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
CKINVDCx14_ASAP7_75t_R g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
AOI21xp5_ASAP7_75t_L g1047 ( .A1(n_1007), .A2(n_1048), .B(n_1053), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1014), .B1(n_1016), .B2(n_1017), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1019 ( .A(n_1020), .Y(n_1019) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1038), .C(n_1056), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1026), .B(n_1055), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1044 ( .A(n_1028), .B(n_1045), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_1028), .B(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1043 ( .A(n_1044), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1051), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1061), .B1(n_1062), .B2(n_1064), .C(n_1066), .Y(n_1056) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
OAI21x1_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1077), .B(n_1093), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1075), .B(n_1087), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g1075 ( .A(n_1076), .Y(n_1075) );
NOR2xp67_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1088), .Y(n_1077) );
NAND3xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1085), .C(n_1087), .Y(n_1078) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1079), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1082), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1095 ( .A(n_1085), .Y(n_1095) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1088), .Y(n_1098) );
NAND4xp25_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1090), .C(n_1091), .D(n_1092), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1098), .Y(n_1093) );
NOR3xp33_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1096), .C(n_1097), .Y(n_1094) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
NOR4xp75_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1112), .C(n_1115), .D(n_1118), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
NAND2xp5_ASAP7_75t_SL g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
OAI21x1_ASAP7_75t_SL g1118 ( .A1(n_1119), .A2(n_1120), .B(n_1121), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
endmodule