module fake_jpeg_11138_n_135 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_50),
.B1(n_21),
.B2(n_28),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_32),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_19),
.B(n_16),
.C(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_27),
.B(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_27),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_21),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_25),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_5),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_73),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_20),
.B1(n_19),
.B2(n_31),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_26),
.B1(n_22),
.B2(n_14),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_20),
.B1(n_14),
.B2(n_26),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_72),
.Y(n_89)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_11),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_37),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_35),
.B1(n_37),
.B2(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_88),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_44),
.C(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_92),
.Y(n_98)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_103),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_67),
.B1(n_75),
.B2(n_83),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_67),
.B1(n_75),
.B2(n_83),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_83),
.B1(n_86),
.B2(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_96),
.B(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_96),
.B(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_100),
.B1(n_99),
.B2(n_86),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_126),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_64),
.B(n_131),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_64),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_64),
.Y(n_135)
);


endmodule