module fake_jpeg_17368_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_0),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_17),
.B(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_20),
.B(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_12),
.C(n_8),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_7),
.B1(n_16),
.B2(n_17),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_27),
.B(n_1),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_19),
.B1(n_13),
.B2(n_20),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_22),
.C(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_34),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_32),
.B(n_28),
.Y(n_37)
);

AOI222xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_35),
.B1(n_30),
.B2(n_6),
.C1(n_5),
.C2(n_22),
.Y(n_38)
);


endmodule