module fake_jpeg_15391_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_46),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_58),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_27),
.B1(n_22),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_73)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_16),
.Y(n_106)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_22),
.B1(n_27),
.B2(n_32),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_19),
.B(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_23),
.B(n_29),
.C(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_19),
.B1(n_20),
.B2(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_36),
.B1(n_38),
.B2(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_36),
.B1(n_38),
.B2(n_25),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_23),
.B1(n_29),
.B2(n_24),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_56),
.B1(n_47),
.B2(n_19),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_28),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_58),
.A3(n_43),
.B1(n_24),
.B2(n_31),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_86),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_47),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_87),
.A2(n_107),
.B(n_30),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_76),
.B1(n_72),
.B2(n_79),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_63),
.B1(n_16),
.B2(n_7),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_108),
.B(n_44),
.Y(n_136)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_109),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_0),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_21),
.B1(n_16),
.B2(n_30),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_48),
.B1(n_51),
.B2(n_44),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_81),
.B1(n_63),
.B2(n_61),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_60),
.B1(n_72),
.B2(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_119),
.B1(n_99),
.B2(n_98),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_83),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_121),
.B(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_118),
.B1(n_122),
.B2(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_61),
.B1(n_78),
.B2(n_81),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_87),
.B(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_63),
.B1(n_48),
.B2(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_51),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_87),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_136),
.B(n_68),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_30),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_93),
.C(n_85),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_89),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_110),
.B1(n_97),
.B2(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_165),
.B1(n_166),
.B2(n_1),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_110),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_146),
.B(n_154),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_111),
.Y(n_144)
);

NAND2xp67_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_107),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_157),
.B(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_153),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_103),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_118),
.A2(n_48),
.B1(n_44),
.B2(n_68),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_156),
.A2(n_117),
.B1(n_147),
.B2(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_1),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_112),
.B1(n_120),
.B2(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_9),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_174),
.C(n_175),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_184),
.B(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_122),
.B1(n_113),
.B2(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_123),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_119),
.B1(n_133),
.B2(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_124),
.B1(n_135),
.B2(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

OAI22x1_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_180),
.B(n_186),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_148),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_150),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_145),
.B(n_10),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_206),
.B1(n_210),
.B2(n_169),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_200),
.B(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NOR4xp25_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_146),
.C(n_161),
.D(n_151),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_157),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_175),
.C(n_174),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_140),
.B(n_154),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_165),
.B(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_149),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_207),
.Y(n_217)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_166),
.B1(n_3),
.B2(n_6),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_173),
.B1(n_177),
.B2(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_223),
.C(n_225),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_191),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_172),
.B1(n_182),
.B2(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_226),
.B1(n_193),
.B2(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_201),
.C(n_205),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_179),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_176),
.B1(n_183),
.B2(n_178),
.Y(n_226)
);

OAI21x1_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_210),
.B(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_210),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_233),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_203),
.B(n_193),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_205),
.C(n_202),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_220),
.C(n_216),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_221),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_228),
.B(n_221),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_225),
.C(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_232),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_254),
.A3(n_244),
.B1(n_252),
.B2(n_253),
.C1(n_246),
.C2(n_239),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_231),
.B1(n_215),
.B2(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_199),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_255),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_235),
.C(n_213),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_198),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_245),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_209),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_260),
.B1(n_8),
.B2(n_5),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_239),
.A3(n_198),
.B1(n_214),
.B2(n_209),
.C1(n_196),
.C2(n_189),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_261),
.B(n_7),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_6),
.C(n_7),
.Y(n_265)
);

OAI311xp33_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_266),
.A3(n_260),
.B1(n_11),
.C1(n_12),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_11),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_12),
.C(n_13),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_14),
.Y(n_272)
);


endmodule