module fake_jpeg_30396_n_405 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_405);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_21),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_46),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_66),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_21),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_49),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_67),
.Y(n_86)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_28),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_76),
.Y(n_109)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

CKINVDCx9p33_ASAP7_75t_R g127 ( 
.A(n_79),
.Y(n_127)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_41),
.Y(n_123)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_42),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_97),
.Y(n_155)
);

INVx2_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_113),
.Y(n_132)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_61),
.A2(n_31),
.B1(n_28),
.B2(n_42),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_125),
.B1(n_69),
.B2(n_52),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_111),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_41),
.Y(n_113)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_48),
.B1(n_25),
.B2(n_34),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_25),
.B1(n_34),
.B2(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_49),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_51),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_82),
.B1(n_81),
.B2(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_50),
.B(n_32),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_131),
.A2(n_105),
.B1(n_36),
.B2(n_39),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_22),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_40),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_149),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_39),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_97),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_127),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_93),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_75),
.C(n_65),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_22),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_22),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_104),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_94),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_172),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_119),
.B1(n_57),
.B2(n_102),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_181),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_128),
.B1(n_122),
.B2(n_115),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_180),
.B1(n_185),
.B2(n_145),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_99),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_128),
.B1(n_64),
.B2(n_62),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

INVx5_ASAP7_75t_SL g189 ( 
.A(n_182),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_143),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_194),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_193),
.B(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_134),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_172),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_186),
.B1(n_170),
.B2(n_173),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_112),
.B1(n_115),
.B2(n_122),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_139),
.B1(n_148),
.B2(n_165),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_175),
.A2(n_144),
.B1(n_166),
.B2(n_130),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_185),
.B1(n_155),
.B2(n_174),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_168),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_226),
.B1(n_200),
.B2(n_166),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_179),
.C(n_150),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_164),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_221),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_166),
.B1(n_189),
.B2(n_190),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_186),
.B(n_156),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_174),
.B(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_186),
.B1(n_166),
.B2(n_180),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_195),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_227),
.A2(n_229),
.B(n_169),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_243),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_195),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_230),
.A2(n_151),
.B1(n_158),
.B2(n_147),
.Y(n_270)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_247),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_208),
.B(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_226),
.B1(n_201),
.B2(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_235),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_204),
.B1(n_144),
.B2(n_141),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_99),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_132),
.Y(n_243)
);

CKINVDCx10_ASAP7_75t_R g244 ( 
.A(n_219),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_203),
.B1(n_205),
.B2(n_189),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_171),
.B1(n_204),
.B2(n_184),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_191),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_211),
.B1(n_223),
.B2(n_217),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_260),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_211),
.C(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_250),
.C(n_247),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_242),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_217),
.B(n_206),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_187),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_116),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_269),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_231),
.A2(n_165),
.B1(n_144),
.B2(n_138),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_149),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_31),
.B1(n_44),
.B2(n_30),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_160),
.B1(n_159),
.B2(n_177),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_238),
.B(n_37),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_37),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_248),
.B1(n_227),
.B2(n_229),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_236),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_276),
.B(n_281),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_279),
.C(n_301),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_249),
.C(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_288),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_239),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_273),
.B(n_263),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_244),
.C(n_232),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_285),
.A2(n_162),
.B(n_152),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_292),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_163),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_SL g289 ( 
.A(n_259),
.B(n_245),
.C(n_202),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_290),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_129),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_271),
.B1(n_254),
.B2(n_178),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_202),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_163),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_263),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_44),
.Y(n_297)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_256),
.A2(n_31),
.B1(n_47),
.B2(n_27),
.Y(n_298)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_177),
.C(n_146),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_270),
.B1(n_274),
.B2(n_267),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_305),
.A2(n_314),
.B1(n_318),
.B2(n_320),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_307),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_251),
.C(n_273),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_102),
.C(n_98),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_311),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_289),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_294),
.A2(n_254),
.B1(n_271),
.B2(n_264),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_299),
.B1(n_277),
.B2(n_286),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_278),
.A2(n_138),
.B1(n_154),
.B2(n_178),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_284),
.A2(n_39),
.B(n_36),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_319),
.A2(n_1),
.B(n_2),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_283),
.A2(n_154),
.B1(n_159),
.B2(n_140),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_92),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_339),
.B1(n_47),
.B2(n_84),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_292),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_332),
.Y(n_355)
);

NAND5xp2_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_276),
.C(n_287),
.D(n_295),
.E(n_161),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_90),
.B(n_114),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_333),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_36),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_96),
.C(n_88),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_338),
.C(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_103),
.C(n_118),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_313),
.A2(n_321),
.B1(n_312),
.B2(n_316),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_2),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_317),
.A2(n_104),
.B(n_161),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_322),
.B1(n_318),
.B2(n_314),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_345),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_315),
.B1(n_304),
.B2(n_322),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_344),
.A2(n_347),
.B1(n_4),
.B2(n_6),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_335),
.A2(n_340),
.B(n_329),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_346),
.B(n_334),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_337),
.A2(n_305),
.B1(n_303),
.B2(n_320),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_349),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_327),
.B(n_1),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_339),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_3),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_161),
.C(n_47),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_342),
.C(n_330),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_356),
.A2(n_337),
.B1(n_326),
.B2(n_338),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_358),
.A2(n_355),
.B(n_354),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_364),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_363),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_86),
.B1(n_8),
.B2(n_9),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_365),
.A2(n_35),
.B1(n_29),
.B2(n_34),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_47),
.C(n_48),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_368),
.C(n_86),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_353),
.A2(n_114),
.B(n_108),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_367),
.A2(n_4),
.B(n_6),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_84),
.C(n_90),
.Y(n_368)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_369),
.Y(n_386)
);

AOI221xp5_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_347),
.B1(n_356),
.B2(n_352),
.C(n_8),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_370),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_372),
.B(n_373),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_108),
.B(n_58),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_374),
.B(n_375),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_357),
.A2(n_56),
.B(n_34),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_377),
.B(n_378),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_34),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_366),
.C(n_35),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_7),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_7),
.Y(n_385)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_385),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_9),
.C(n_10),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_388),
.A2(n_389),
.B(n_376),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_10),
.C(n_12),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_391),
.B(n_392),
.Y(n_396)
);

O2A1O1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_387),
.A2(n_376),
.B(n_370),
.C(n_15),
.Y(n_393)
);

AOI322xp5_ASAP7_75t_L g398 ( 
.A1(n_393),
.A2(n_383),
.A3(n_384),
.B1(n_382),
.B2(n_17),
.C1(n_18),
.C2(n_14),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_12),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_14),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_397),
.A2(n_398),
.B(n_399),
.Y(n_400)
);

AOI322xp5_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_19),
.C1(n_29),
.C2(n_35),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_396),
.A2(n_390),
.B(n_16),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_402),
.A2(n_400),
.B(n_16),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_15),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_19),
.Y(n_405)
);


endmodule