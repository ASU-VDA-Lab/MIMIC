module fake_jpeg_13955_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_16),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

CKINVDCx6p67_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_62),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_72),
.Y(n_89)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_75),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_52),
.C(n_58),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_71),
.B(n_70),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_78),
.B1(n_50),
.B2(n_51),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_51),
.B1(n_50),
.B2(n_63),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_114),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_61),
.Y(n_140)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_123),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_124),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_87),
.B(n_66),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_25),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_129),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_0),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_67),
.C(n_66),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_145),
.C(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_1),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_61),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_2),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_2),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_3),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_5),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_6),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_6),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_67),
.B1(n_27),
.B2(n_30),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_133),
.C(n_129),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_163),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_126),
.B1(n_130),
.B2(n_147),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_12),
.C(n_13),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_15),
.C(n_17),
.Y(n_164)
);

NOR4xp25_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_19),
.C(n_21),
.D(n_22),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_170),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_26),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_175),
.B1(n_172),
.B2(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_154),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_176),
.C(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_160),
.B1(n_152),
.B2(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_168),
.B(n_160),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_155),
.A3(n_156),
.B1(n_169),
.B2(n_40),
.C1(n_41),
.C2(n_42),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_181),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_32),
.B(n_33),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_39),
.Y(n_184)
);


endmodule