module fake_jpeg_1424_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_7),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_19),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_39),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_0),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_3),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_27),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_25),
.B1(n_14),
.B2(n_16),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_28),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_60),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_30),
.A2(n_13),
.A3(n_15),
.B1(n_20),
.B2(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_61),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_0),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_31),
.B(n_35),
.C(n_36),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_39),
.B(n_33),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_44),
.B(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_35),
.B1(n_6),
.B2(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_44),
.B1(n_63),
.B2(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_6),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_46),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_88),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_75),
.B1(n_68),
.B2(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_69),
.Y(n_101)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_46),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_74),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_74),
.B1(n_68),
.B2(n_64),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_92),
.B1(n_66),
.B2(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_46),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_84),
.B(n_88),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_86),
.B(n_89),
.Y(n_104)
);

INVxp33_ASAP7_75t_SL g112 ( 
.A(n_104),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_108),
.C(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_93),
.B(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_100),
.B1(n_96),
.B2(n_95),
.Y(n_116)
);

AO221x1_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_98),
.B1(n_85),
.B2(n_90),
.C(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_110),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_104),
.C(n_93),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_91),
.C(n_80),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_112),
.B(n_113),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_124),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_91),
.B1(n_56),
.B2(n_45),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_125),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_76),
.Y(n_129)
);


endmodule