module fake_netlist_6_2783_n_918 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_918);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_918;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_859;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_386;
wire n_201;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_816;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_9),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_31),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_52),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_86),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_44),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_73),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_17),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_46),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_133),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_28),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_79),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_18),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_67),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_87),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_135),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_101),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_70),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_56),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_127),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_128),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_42),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_81),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_98),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_111),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_106),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_24),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_182),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_59),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_80),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_69),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_76),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_97),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_4),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_164),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_75),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_144),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_162),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_110),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_66),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_161),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

BUFx8_ASAP7_75t_SL g262 ( 
.A(n_137),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_45),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_104),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_130),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_117),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_134),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_183),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_141),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_77),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_27),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_35),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_15),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_4),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_116),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_48),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_1),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_109),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_38),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_9),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_185),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_216),
.B(n_0),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_0),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_191),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_248),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_1),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_195),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_199),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_201),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_204),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_214),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_197),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_206),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_207),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_208),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_233),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_197),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_203),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_211),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_213),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_203),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_233),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_220),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_215),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_232),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_189),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_278),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_190),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_222),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_223),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_227),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_228),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_193),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_268),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_194),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_196),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_268),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_221),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_198),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_283),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_283),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_205),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_231),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_234),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_231),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_210),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_219),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_236),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_287),
.B(n_296),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_300),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_345),
.B(n_192),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_286),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_305),
.B(n_273),
.Y(n_364)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_340),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_273),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_312),
.B(n_273),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_292),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_345),
.A2(n_264),
.B1(n_209),
.B2(n_217),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_304),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_289),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_290),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_284),
.B(n_221),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_230),
.B(n_192),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_303),
.Y(n_383)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_230),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_298),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_299),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_301),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_322),
.B(n_263),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_320),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_272),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_293),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_285),
.A2(n_272),
.B(n_229),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_329),
.A2(n_235),
.B(n_225),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_307),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_313),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_314),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_348),
.B(n_221),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_241),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_319),
.B(n_238),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_397),
.A2(n_267),
.B1(n_350),
.B2(n_246),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_267),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_370),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_394),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_394),
.B(n_302),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_367),
.B(n_327),
.Y(n_417)
);

NOR2x1p5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_336),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_267),
.B1(n_243),
.B2(n_247),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_330),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_375),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_332),
.C(n_331),
.Y(n_424)
);

BUFx10_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_R g431 ( 
.A(n_362),
.B(n_346),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_387),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_396),
.B(n_336),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_316),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_338),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_224),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_394),
.Y(n_442)
);

OAI22xp33_ASAP7_75t_L g443 ( 
.A1(n_371),
.A2(n_394),
.B1(n_407),
.B2(n_395),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_408),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_338),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_385),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_386),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_404),
.B(n_368),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_365),
.B(n_342),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_342),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_389),
.B(n_250),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_368),
.B(n_267),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_365),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_390),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_259),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_377),
.B(n_367),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_367),
.B(n_261),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_361),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_380),
.B(n_239),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_359),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_380),
.A2(n_265),
.B1(n_240),
.B2(n_266),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

INVx4_ASAP7_75t_SL g473 ( 
.A(n_380),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_392),
.B(n_343),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_357),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_360),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_392),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_364),
.Y(n_481)
);

OAI221xp5_ASAP7_75t_L g482 ( 
.A1(n_410),
.A2(n_384),
.B1(n_378),
.B2(n_360),
.C(n_379),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_477),
.Y(n_484)
);

AO22x2_ASAP7_75t_L g485 ( 
.A1(n_414),
.A2(n_364),
.B1(n_369),
.B2(n_291),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

AOI22x1_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_369),
.B1(n_409),
.B2(n_378),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_415),
.B(n_379),
.Y(n_491)
);

OAI221xp5_ASAP7_75t_L g492 ( 
.A1(n_420),
.A2(n_384),
.B1(n_374),
.B2(n_366),
.C(n_372),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_423),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_427),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_466),
.A2(n_380),
.B1(n_382),
.B2(n_398),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_452),
.B(n_353),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_439),
.B(n_409),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_417),
.B(n_421),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_437),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

BUFx8_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_455),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_478),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

OAI221xp5_ASAP7_75t_L g508 ( 
.A1(n_470),
.A2(n_366),
.B1(n_372),
.B2(n_374),
.C(n_405),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_463),
.A2(n_343),
.B1(n_291),
.B2(n_310),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_448),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_450),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_439),
.A2(n_451),
.B1(n_415),
.B2(n_443),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_432),
.Y(n_513)
);

AO22x2_ASAP7_75t_L g514 ( 
.A1(n_426),
.A2(n_294),
.B1(n_310),
.B2(n_334),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_445),
.B(n_400),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_431),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_451),
.A2(n_380),
.B1(n_400),
.B2(n_242),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_455),
.B(n_294),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_430),
.B(n_366),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_436),
.A2(n_334),
.B1(n_3),
.B2(n_5),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_459),
.B(n_372),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_471),
.B(n_382),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_449),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_425),
.B(n_374),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_469),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_451),
.B(n_472),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_438),
.B(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_464),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_380),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_458),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_425),
.B(n_365),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_456),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_458),
.B(n_380),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_458),
.B(n_359),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_434),
.A2(n_424),
.B1(n_458),
.B2(n_416),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_441),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_441),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_517),
.B(n_418),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_479),
.B(n_467),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_SL g549 ( 
.A(n_481),
.B(n_433),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_479),
.B(n_473),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_499),
.B(n_473),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_SL g552 ( 
.A(n_504),
.B(n_460),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_544),
.B(n_468),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_457),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_497),
.B(n_441),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_534),
.B(n_454),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_498),
.B(n_454),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_530),
.B(n_454),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_529),
.B(n_244),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_491),
.B(n_461),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_491),
.B(n_461),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_522),
.B(n_461),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_521),
.B(n_245),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_522),
.B(n_249),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_532),
.B(n_251),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_SL g566 ( 
.A(n_509),
.B(n_252),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_512),
.B(n_254),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_486),
.B(n_255),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_503),
.B(n_487),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_490),
.B(n_256),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_493),
.B(n_257),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_494),
.B(n_269),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_496),
.B(n_270),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_500),
.B(n_271),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_501),
.B(n_276),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_489),
.B(n_515),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_515),
.B(n_277),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_480),
.B(n_413),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_488),
.B(n_279),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_480),
.B(n_413),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_505),
.B(n_280),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_510),
.B(n_355),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_511),
.B(n_355),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_516),
.B(n_356),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_533),
.B(n_537),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_538),
.B(n_356),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_518),
.B(n_351),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_524),
.B(n_351),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_485),
.B(n_457),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_413),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_483),
.B(n_352),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_484),
.B(n_352),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_484),
.B(n_357),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_519),
.B(n_357),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_485),
.B(n_462),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_525),
.B(n_358),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_525),
.B(n_413),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_528),
.B(n_358),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_528),
.B(n_358),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_462),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_506),
.B(n_354),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_545),
.B(n_354),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_495),
.B(n_354),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_536),
.B(n_29),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_535),
.B(n_32),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_548),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_566),
.A2(n_482),
.B(n_508),
.C(n_540),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_553),
.A2(n_546),
.B(n_545),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_558),
.B(n_546),
.Y(n_609)
);

OAI21x1_ASAP7_75t_SL g610 ( 
.A1(n_600),
.A2(n_541),
.B(n_542),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_554),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_576),
.A2(n_507),
.B(n_527),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_591),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_603),
.A2(n_543),
.B(n_531),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_569),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_555),
.B(n_526),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_560),
.B(n_526),
.Y(n_617)
);

AO31x2_ASAP7_75t_L g618 ( 
.A1(n_578),
.A2(n_492),
.A3(n_539),
.B(n_526),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_567),
.B(n_539),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_550),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_556),
.B(n_577),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_594),
.A2(n_523),
.B(n_95),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_547),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_561),
.A2(n_523),
.B(n_94),
.Y(n_624)
);

OAI22x1_ASAP7_75t_L g625 ( 
.A1(n_589),
.A2(n_514),
.B1(n_502),
.B2(n_7),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_602),
.A2(n_93),
.B(n_188),
.Y(n_626)
);

AO31x2_ASAP7_75t_L g627 ( 
.A1(n_580),
.A2(n_514),
.A3(n_6),
.B(n_7),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_604),
.A2(n_502),
.B(n_8),
.C(n_10),
.Y(n_628)
);

AOI221x1_ASAP7_75t_L g629 ( 
.A1(n_585),
.A2(n_595),
.B1(n_565),
.B2(n_574),
.C(n_572),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_562),
.B(n_2),
.Y(n_630)
);

AOI221xp5_ASAP7_75t_SL g631 ( 
.A1(n_605),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_557),
.B(n_593),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_570),
.B(n_12),
.Y(n_633)
);

O2A1O1Ixp5_ASAP7_75t_L g634 ( 
.A1(n_586),
.A2(n_100),
.B(n_181),
.C(n_180),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_592),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_549),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_552),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_R g638 ( 
.A(n_563),
.B(n_34),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_604),
.A2(n_99),
.B(n_177),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_590),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_551),
.A2(n_96),
.B(n_176),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_597),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_605),
.A2(n_92),
.B(n_173),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_564),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_596),
.A2(n_91),
.B(n_172),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_571),
.A2(n_90),
.B(n_171),
.Y(n_646)
);

AO32x2_ASAP7_75t_L g647 ( 
.A1(n_568),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_601),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_573),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_598),
.A2(n_102),
.B(n_170),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_599),
.A2(n_89),
.B(n_168),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_575),
.B(n_13),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_612),
.A2(n_588),
.B(n_587),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_620),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_L g655 ( 
.A1(n_644),
.A2(n_628),
.B1(n_622),
.B2(n_624),
.C(n_649),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_611),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_621),
.A2(n_581),
.B1(n_579),
.B2(n_582),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_606),
.Y(n_658)
);

AO31x2_ASAP7_75t_L g659 ( 
.A1(n_607),
.A2(n_584),
.A3(n_583),
.B(n_559),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_609),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_615),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_620),
.B(n_36),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_636),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_609),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_633),
.B(n_16),
.C(n_17),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_614),
.A2(n_105),
.B(n_167),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_636),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_608),
.A2(n_103),
.B(n_166),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_37),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_619),
.B(n_19),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_613),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_652),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_625),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_620),
.Y(n_674)
);

AO22x2_ASAP7_75t_L g675 ( 
.A1(n_629),
.A2(n_647),
.B1(n_610),
.B2(n_631),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_642),
.A2(n_108),
.B(n_158),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_642),
.A2(n_85),
.B(n_157),
.Y(n_677)
);

OA21x2_ASAP7_75t_L g678 ( 
.A1(n_631),
.A2(n_23),
.B(n_25),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_623),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_SL g680 ( 
.A1(n_616),
.A2(n_25),
.B(n_26),
.C(n_39),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_617),
.A2(n_113),
.B(n_40),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_618),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_645),
.A2(n_114),
.B(n_41),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_626),
.A2(n_115),
.B(n_43),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_640),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_635),
.Y(n_686)
);

AO21x2_ASAP7_75t_L g687 ( 
.A1(n_650),
.A2(n_118),
.B(n_49),
.Y(n_687)
);

OAI21x1_ASAP7_75t_SL g688 ( 
.A1(n_650),
.A2(n_119),
.B(n_50),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_630),
.A2(n_120),
.B(n_51),
.Y(n_689)
);

AO21x2_ASAP7_75t_L g690 ( 
.A1(n_651),
.A2(n_121),
.B(n_53),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_638),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_639),
.A2(n_123),
.B(n_54),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_634),
.A2(n_632),
.B(n_643),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_648),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_660),
.B(n_618),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_686),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_682),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_656),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_618),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_661),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_656),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_686),
.Y(n_702)
);

BUFx5_ASAP7_75t_L g703 ( 
.A(n_664),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_655),
.A2(n_641),
.B(n_646),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_675),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_671),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_654),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_694),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_675),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_679),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_666),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_653),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_659),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_662),
.B(n_659),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_675),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_667),
.A2(n_651),
.B1(n_648),
.B2(n_647),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_678),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_678),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_678),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_670),
.B(n_627),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_659),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_683),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_676),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_663),
.B(n_627),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_677),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_684),
.A2(n_627),
.B(n_647),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_684),
.A2(n_124),
.B(n_55),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_687),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_687),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_659),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_693),
.A2(n_131),
.B(n_57),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_690),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_658),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_690),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_662),
.B(n_139),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_679),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_658),
.Y(n_738)
);

CKINVDCx11_ASAP7_75t_R g739 ( 
.A(n_669),
.Y(n_739)
);

NAND2x1_ASAP7_75t_L g740 ( 
.A(n_688),
.B(n_184),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_700),
.B(n_685),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_R g743 ( 
.A(n_735),
.B(n_691),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_SL g744 ( 
.A(n_736),
.B(n_691),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_710),
.B(n_685),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_710),
.B(n_669),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_710),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_706),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_737),
.B(n_738),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_698),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_R g751 ( 
.A(n_735),
.B(n_669),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_736),
.B(n_654),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_698),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_R g754 ( 
.A(n_739),
.B(n_674),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_R g755 ( 
.A(n_720),
.B(n_674),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_698),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_706),
.B(n_673),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_701),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_733),
.B(n_673),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_R g760 ( 
.A(n_720),
.B(n_714),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_R g761 ( 
.A(n_714),
.B(n_689),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_696),
.B(n_665),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_701),
.Y(n_763)
);

XNOR2xp5_ASAP7_75t_L g764 ( 
.A(n_701),
.B(n_657),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_707),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_696),
.B(n_672),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_736),
.B(n_654),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_697),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_736),
.B(n_654),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_702),
.B(n_680),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_707),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_702),
.B(n_681),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_695),
.B(n_668),
.Y(n_773)
);

XNOR2xp5_ASAP7_75t_L g774 ( 
.A(n_714),
.B(n_692),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_R g775 ( 
.A(n_703),
.B(n_112),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_708),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_703),
.B(n_156),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_708),
.B(n_83),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_750),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_768),
.B(n_715),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_769),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_748),
.B(n_705),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_773),
.B(n_705),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_769),
.B(n_714),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_764),
.A2(n_704),
.B1(n_716),
.B2(n_740),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_776),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_742),
.B(n_695),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_755),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_770),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_751),
.A2(n_741),
.B1(n_703),
.B2(n_740),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_772),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_749),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_774),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_762),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_766),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_753),
.B(n_709),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_756),
.B(n_26),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_758),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_763),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_745),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_746),
.A2(n_724),
.B1(n_741),
.B2(n_703),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_778),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_759),
.B(n_703),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_746),
.A2(n_703),
.B1(n_709),
.B2(n_715),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_745),
.B(n_713),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_765),
.B(n_703),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_747),
.B(n_703),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_779),
.Y(n_809)
);

AND2x2_ASAP7_75t_SL g810 ( 
.A(n_788),
.B(n_760),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_780),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_780),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_796),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_786),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_795),
.B(n_703),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_782),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_795),
.B(n_697),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_786),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_782),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_795),
.B(n_728),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_798),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_793),
.B(n_754),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_783),
.B(n_721),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_784),
.B(n_712),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_810),
.B(n_790),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_816),
.B(n_793),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_813),
.B(n_783),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_813),
.B(n_803),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_816),
.B(n_784),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_821),
.B(n_787),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_819),
.B(n_814),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_811),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_810),
.B(n_784),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_824),
.B(n_784),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_SL g835 ( 
.A(n_833),
.B(n_743),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_834),
.B(n_822),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_826),
.B(n_818),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_825),
.A2(n_785),
.B1(n_790),
.B2(n_801),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_830),
.B(n_804),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_825),
.B(n_775),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_839),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_SL g842 ( 
.A1(n_838),
.A2(n_797),
.B(n_792),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_837),
.B(n_828),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_836),
.B(n_829),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_840),
.B(n_809),
.Y(n_845)
);

AOI311xp33_ASAP7_75t_L g846 ( 
.A1(n_841),
.A2(n_804),
.A3(n_794),
.B(n_789),
.C(n_812),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_843),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_845),
.A2(n_835),
.B1(n_827),
.B2(n_809),
.Y(n_848)
);

OAI221xp5_ASAP7_75t_L g849 ( 
.A1(n_842),
.A2(n_794),
.B1(n_832),
.B2(n_800),
.C(n_744),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_847),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_849),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_848),
.B(n_844),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_850),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_851),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_852),
.B(n_845),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_850),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_853),
.B(n_831),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_856),
.B(n_846),
.C(n_771),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_855),
.B(n_854),
.C(n_809),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_SL g860 ( 
.A(n_855),
.B(n_777),
.C(n_808),
.Y(n_860)
);

NOR4xp25_ASAP7_75t_SL g861 ( 
.A(n_853),
.B(n_761),
.C(n_799),
.D(n_789),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_L g862 ( 
.A(n_853),
.B(n_791),
.C(n_798),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_853),
.B(n_799),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_858),
.A2(n_791),
.B(n_807),
.Y(n_864)
);

AOI222xp33_ASAP7_75t_L g865 ( 
.A1(n_860),
.A2(n_734),
.B1(n_728),
.B2(n_729),
.C1(n_732),
.C2(n_798),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_859),
.A2(n_781),
.B1(n_779),
.B2(n_802),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_863),
.B(n_857),
.Y(n_867)
);

OAI221xp5_ASAP7_75t_SL g868 ( 
.A1(n_862),
.A2(n_861),
.B1(n_779),
.B2(n_805),
.C(n_820),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_857),
.Y(n_869)
);

AOI221xp5_ASAP7_75t_L g870 ( 
.A1(n_858),
.A2(n_734),
.B1(n_729),
.B2(n_732),
.C(n_817),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_859),
.A2(n_824),
.B1(n_781),
.B2(n_796),
.Y(n_871)
);

AND2x2_ASAP7_75t_SL g872 ( 
.A(n_859),
.B(n_781),
.Y(n_872)
);

NOR2x1_ASAP7_75t_L g873 ( 
.A(n_869),
.B(n_752),
.Y(n_873)
);

OAI211xp5_ASAP7_75t_SL g874 ( 
.A1(n_870),
.A2(n_802),
.B(n_815),
.C(n_725),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_867),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_871),
.B(n_58),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_872),
.Y(n_877)
);

NOR2x1_ASAP7_75t_L g878 ( 
.A(n_864),
.B(n_767),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_L g879 ( 
.A(n_868),
.B(n_731),
.C(n_727),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_865),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_SL g881 ( 
.A(n_875),
.B(n_866),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_SL g882 ( 
.A(n_877),
.B(n_802),
.C(n_725),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_880),
.B(n_873),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_R g884 ( 
.A(n_876),
.B(n_60),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_879),
.B(n_820),
.C(n_781),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_878),
.B(n_781),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_R g887 ( 
.A(n_874),
.B(n_62),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_875),
.B(n_824),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_875),
.B(n_63),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_R g890 ( 
.A(n_875),
.B(n_64),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_883),
.A2(n_731),
.B(n_727),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_881),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_886),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_888),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_889),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_890),
.B(n_884),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_885),
.Y(n_897)
);

XOR2xp5_ASAP7_75t_L g898 ( 
.A(n_882),
.B(n_65),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_887),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_888),
.B(n_823),
.Y(n_900)
);

XOR2x1_ASAP7_75t_L g901 ( 
.A(n_899),
.B(n_68),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_892),
.A2(n_820),
.B1(n_767),
.B2(n_752),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_893),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_894),
.A2(n_723),
.B1(n_699),
.B2(n_719),
.Y(n_904)
);

NAND4xp25_ASAP7_75t_L g905 ( 
.A(n_896),
.B(n_723),
.C(n_823),
.D(n_806),
.Y(n_905)
);

AOI21xp33_ASAP7_75t_L g906 ( 
.A1(n_897),
.A2(n_72),
.B(n_74),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_903),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_901),
.B(n_895),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_905),
.A2(n_898),
.B1(n_900),
.B2(n_891),
.Y(n_909)
);

AOI31xp33_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_908),
.A3(n_906),
.B(n_909),
.Y(n_910)
);

AOI31xp33_ASAP7_75t_L g911 ( 
.A1(n_907),
.A2(n_898),
.A3(n_902),
.B(n_904),
.Y(n_911)
);

OAI322xp33_ASAP7_75t_L g912 ( 
.A1(n_910),
.A2(n_718),
.A3(n_717),
.B1(n_719),
.B2(n_711),
.C1(n_143),
.C2(n_147),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_911),
.A2(n_806),
.B1(n_722),
.B2(n_717),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_912),
.A2(n_722),
.B1(n_713),
.B2(n_730),
.Y(n_914)
);

AOI222xp33_ASAP7_75t_L g915 ( 
.A1(n_913),
.A2(n_718),
.B1(n_726),
.B2(n_722),
.C1(n_142),
.C2(n_148),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_915),
.Y(n_916)
);

AOI221xp5_ASAP7_75t_L g917 ( 
.A1(n_916),
.A2(n_914),
.B1(n_82),
.B2(n_140),
.C(n_151),
.Y(n_917)
);

AOI211xp5_ASAP7_75t_L g918 ( 
.A1(n_917),
.A2(n_78),
.B(n_153),
.C(n_154),
.Y(n_918)
);


endmodule