module fake_netlist_6_895_n_28 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_28);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_28;

wire n_16;
wire n_21;
wire n_10;
wire n_24;
wire n_18;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_19;
wire n_25;

INVx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

AND2x4_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

OAI21x1_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_12),
.B(n_11),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_7),
.B(n_9),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

OAI221xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_13),
.B1(n_11),
.B2(n_19),
.C(n_10),
.Y(n_23)
);

NAND3x1_ASAP7_75t_SL g24 ( 
.A(n_23),
.B(n_15),
.C(n_1),
.Y(n_24)
);

AOI211xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_19),
.B(n_12),
.C(n_15),
.Y(n_25)
);

OR3x2_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_0),
.C(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_25),
.Y(n_27)
);

AOI222xp33_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_0),
.B1(n_13),
.B2(n_15),
.C1(n_18),
.C2(n_26),
.Y(n_28)
);


endmodule