module fake_jpeg_15446_n_166 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_166);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_64),
.B1(n_48),
.B2(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_102),
.Y(n_120)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_59),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_51),
.B1(n_64),
.B2(n_60),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_113),
.B1(n_114),
.B2(n_0),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_63),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_58),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_59),
.B1(n_65),
.B2(n_50),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_54),
.B(n_62),
.C(n_53),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_114),
.B(n_108),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_104),
.B1(n_125),
.B2(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_57),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_123),
.B1(n_99),
.B2(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_126),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_3),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_96),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_128),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_131),
.B(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_21),
.B1(n_45),
.B2(n_44),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_124),
.B1(n_115),
.B2(n_103),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_120),
.C(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_133),
.B(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_139),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_139),
.B(n_22),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_151),
.C(n_146),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_148),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_152),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_46),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_20),
.Y(n_158)
);

NAND4xp25_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_19),
.C(n_40),
.D(n_37),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_18),
.C(n_35),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_15),
.B(n_33),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_10),
.C(n_32),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_42),
.B(n_31),
.C(n_30),
.D(n_24),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_4),
.B(n_7),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_4),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_7),
.B(n_8),
.Y(n_166)
);


endmodule