module fake_ariane_1269_n_170 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_170);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_170;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

NOR2xp67_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_36),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_0),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_1),
.Y(n_73)
);

BUFx6f_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_2),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_7),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_11),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NAND2x1p5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_13),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_17),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_39),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_52),
.B(n_22),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_55),
.B(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_57),
.B(n_46),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_58),
.B(n_56),
.C(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_56),
.B(n_49),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_24),
.B(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_28),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_30),
.B(n_32),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_37),
.C(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_79),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_71),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_85),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_87),
.B(n_73),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_91),
.C(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_77),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_90),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_90),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_116),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_115),
.C(n_118),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_75),
.B1(n_122),
.B2(n_99),
.C(n_101),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_108),
.B(n_90),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_108),
.C(n_74),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_108),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_90),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_129),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_126),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_129),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_144),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_154),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_141),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_152),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_143),
.C(n_158),
.Y(n_162)
);

NOR3x1_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_140),
.C(n_149),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_157),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_162),
.Y(n_166)
);

AOI211xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_163),
.B(n_157),
.C(n_155),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_148),
.B1(n_153),
.B2(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_150),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_126),
.B1(n_142),
.B2(n_147),
.C(n_75),
.Y(n_170)
);


endmodule