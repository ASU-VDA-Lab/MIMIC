module fake_jpeg_31453_n_434 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_434);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_434;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_50),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g153 ( 
.A(n_51),
.Y(n_153)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_14),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_70),
.B(n_82),
.Y(n_144)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_14),
.B(n_10),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_90),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_89),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_24),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_38),
.Y(n_155)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_38),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_95),
.Y(n_117)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_43),
.A2(n_10),
.B(n_3),
.Y(n_94)
);

NAND2x1p5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_38),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_103),
.A2(n_111),
.B1(n_34),
.B2(n_23),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_41),
.B1(n_24),
.B2(n_44),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_105),
.A2(n_106),
.B1(n_116),
.B2(n_131),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_24),
.B1(n_44),
.B2(n_23),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_13),
.B(n_3),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_108),
.A2(n_11),
.B(n_3),
.C(n_6),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_22),
.B1(n_37),
.B2(n_36),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_113),
.B(n_138),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_20),
.B1(n_35),
.B2(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_135),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_17),
.B1(n_35),
.B2(n_20),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_22),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_32),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_34),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_47),
.A2(n_15),
.B1(n_33),
.B2(n_30),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_73),
.B1(n_69),
.B2(n_80),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_50),
.B(n_32),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_78),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_61),
.B(n_30),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_17),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_171),
.Y(n_209)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_170),
.A2(n_177),
.B(n_193),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_176),
.B1(n_179),
.B2(n_105),
.Y(n_207)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_128),
.A2(n_89),
.B1(n_86),
.B2(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_180),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_126),
.A2(n_76),
.B1(n_68),
.B2(n_9),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_186),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_183),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_101),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_113),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_192),
.B1(n_11),
.B2(n_12),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_6),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_178),
.B1(n_183),
.B2(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_195),
.Y(n_227)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_115),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_196),
.Y(n_215)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_177),
.B1(n_193),
.B2(n_172),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_207),
.A2(n_165),
.B1(n_139),
.B2(n_199),
.Y(n_260)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_187),
.A3(n_161),
.B1(n_167),
.B2(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_160),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_134),
.C(n_129),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_220),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_219),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_216),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_116),
.C(n_131),
.Y(n_220)
);

AO22x2_ASAP7_75t_L g224 ( 
.A1(n_159),
.A2(n_100),
.B1(n_106),
.B2(n_133),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_173),
.Y(n_238)
);

AOI22x1_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_185),
.B1(n_100),
.B2(n_194),
.Y(n_235)
);

AOI22x1_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_145),
.B1(n_132),
.B2(n_164),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_260),
.B1(n_228),
.B2(n_214),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_240),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_241),
.B(n_242),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_222),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_243),
.B(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_166),
.B1(n_170),
.B2(n_187),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_252),
.B1(n_211),
.B2(n_221),
.Y(n_265)
);

NAND2x1p5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_162),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_263),
.B(n_224),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_227),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_253),
.B(n_254),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_212),
.B1(n_204),
.B2(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_166),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_181),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_195),
.B(n_139),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_267),
.B1(n_273),
.B2(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_211),
.B1(n_224),
.B2(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_287),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_210),
.C(n_215),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_288),
.C(n_248),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_224),
.B1(n_235),
.B2(n_233),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_284),
.B(n_273),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_283),
.B1(n_252),
.B2(n_253),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_202),
.B1(n_223),
.B2(n_228),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_202),
.B(n_229),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_205),
.B(n_218),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_237),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_229),
.C(n_236),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_254),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_291),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_293),
.A2(n_294),
.B1(n_301),
.B2(n_282),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_246),
.B1(n_252),
.B2(n_260),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_251),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_300),
.C(n_269),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_256),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_303),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_302),
.B(n_268),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_240),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_308),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_246),
.B1(n_239),
.B2(n_234),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_255),
.B(n_262),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_307),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_274),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_268),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_201),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_267),
.A2(n_239),
.B1(n_217),
.B2(n_242),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_280),
.B1(n_285),
.B2(n_276),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_236),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_297),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_328),
.Y(n_353)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_322),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_301),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_290),
.B(n_286),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_332),
.C(n_336),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_326),
.A2(n_294),
.B1(n_304),
.B2(n_309),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_334),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_289),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_278),
.C(n_285),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_280),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_270),
.C(n_265),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_298),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_345),
.C(n_352),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_296),
.Y(n_341)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_343),
.A2(n_351),
.B1(n_333),
.B2(n_327),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_304),
.B1(n_292),
.B2(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_292),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_329),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_356),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_337),
.B(n_334),
.C(n_315),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_331),
.A2(n_290),
.B1(n_311),
.B2(n_286),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_243),
.C(n_217),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_200),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_335),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_218),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_358),
.C(n_330),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_231),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_335),
.C(n_315),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_359),
.A2(n_361),
.B1(n_349),
.B2(n_346),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_323),
.B(n_337),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_363),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_357),
.B1(n_348),
.B2(n_351),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_340),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_365),
.A2(n_346),
.B(n_349),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_368),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_326),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_345),
.B(n_319),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_366),
.Y(n_383)
);

XOR2x2_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_319),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_373),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_372),
.C(n_355),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_330),
.C(n_231),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_347),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_370),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_382),
.C(n_387),
.Y(n_390)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_380),
.A2(n_368),
.B1(n_359),
.B2(n_361),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_384),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_350),
.C(n_352),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_389),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_353),
.B1(n_249),
.B2(n_206),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_353),
.B1(n_249),
.B2(n_206),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_385),
.B(n_374),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_205),
.C(n_157),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_188),
.C(n_168),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_169),
.C(n_189),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_230),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_391),
.A2(n_400),
.B1(n_387),
.B2(n_376),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_360),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_395),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_397),
.B1(n_402),
.B2(n_383),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_360),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_369),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_104),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_365),
.B(n_230),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_399),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_191),
.B1(n_175),
.B2(n_184),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_388),
.A2(n_112),
.B(n_102),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_401),
.B(n_98),
.Y(n_409)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_405),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_376),
.C(n_133),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_143),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_104),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_410),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_121),
.C(n_152),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_412),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_391),
.C(n_392),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_406),
.A2(n_400),
.B(n_399),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_414),
.A2(n_12),
.B(n_13),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_417),
.A2(n_411),
.B1(n_152),
.B2(n_119),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_412),
.B(n_12),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_418),
.B(n_419),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_405),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_420),
.C(n_416),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_421),
.A2(n_423),
.B(n_425),
.Y(n_427)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_422),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_408),
.C(n_120),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_415),
.C(n_417),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_119),
.C(n_120),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_SL g431 ( 
.A(n_429),
.B(n_430),
.C(n_427),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_SL g430 ( 
.A1(n_426),
.A2(n_13),
.B(n_0),
.C(n_154),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_154),
.B(n_123),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_154),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_0),
.Y(n_434)
);


endmodule