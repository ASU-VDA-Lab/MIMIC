module fake_aes_1664_n_44 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_44);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
BUFx6f_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_4), .B(n_5), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_15), .B(n_0), .C(n_1), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_17), .B(n_0), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_14), .B(n_1), .Y(n_22) );
BUFx12f_ASAP7_75t_L g23 ( .A(n_11), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_16), .B1(n_11), .B2(n_13), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_13), .B1(n_11), .B2(n_4), .Y(n_25) );
BUFx12f_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_22), .A2(n_2), .B1(n_3), .B2(n_7), .Y(n_27) );
NOR4xp25_ASAP7_75t_SL g28 ( .A(n_27), .B(n_19), .C(n_20), .D(n_21), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_24), .B(n_20), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_25), .B(n_21), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_30), .B(n_26), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_18), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_31), .Y(n_35) );
NAND4xp75_ASAP7_75t_L g36 ( .A(n_33), .B(n_28), .C(n_3), .D(n_23), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NAND2xp5_ASAP7_75t_SL g38 ( .A(n_34), .B(n_18), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_37), .B(n_18), .Y(n_39) );
NAND2xp5_ASAP7_75t_L g40 ( .A(n_36), .B(n_38), .Y(n_40) );
NAND2xp5_ASAP7_75t_L g41 ( .A(n_36), .B(n_23), .Y(n_41) );
OR2x6_ASAP7_75t_L g42 ( .A(n_41), .B(n_40), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_39), .Y(n_43) );
XOR2xp5_ASAP7_75t_L g44 ( .A(n_43), .B(n_42), .Y(n_44) );
endmodule