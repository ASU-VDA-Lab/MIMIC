module real_jpeg_9228_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_341, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_341;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_1),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_49),
.B1(n_51),
.B2(n_94),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_94),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_69),
.B1(n_70),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_3),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_49),
.B1(n_51),
.B2(n_99),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_99),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_99),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_4),
.A2(n_35),
.B1(n_69),
.B2(n_70),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_4),
.A2(n_35),
.B1(n_49),
.B2(n_51),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_23),
.B1(n_25),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_10),
.A2(n_61),
.B1(n_69),
.B2(n_70),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_49),
.B1(n_51),
.B2(n_61),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_49),
.B1(n_51),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_11),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_106),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_106),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_51),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_12),
.B(n_51),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_12),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_12),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_26),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_12),
.A2(n_28),
.B(n_30),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_115),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_24),
.B1(n_49),
.B2(n_51),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_14),
.A2(n_24),
.B1(n_69),
.B2(n_70),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_15),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_15),
.A2(n_49),
.B1(n_51),
.B2(n_63),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_339),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_81),
.B(n_337),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_21),
.A2(n_37),
.B(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_22),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_22),
.A2(n_26),
.B(n_36),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_27),
.B(n_32),
.C(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_32),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_23),
.A2(n_32),
.B(n_115),
.C(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_34),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_26),
.A2(n_36),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_27),
.A2(n_37),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_27),
.A2(n_37),
.B1(n_212),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_27),
.A2(n_37),
.B1(n_221),
.B2(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_27),
.A2(n_33),
.B(n_60),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_30),
.A2(n_46),
.B(n_47),
.C(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_47),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g145 ( 
.A(n_30),
.B(n_115),
.CON(n_145),
.SN(n_145)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_36),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_37),
.A2(n_78),
.B(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_40),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_75),
.C(n_79),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_41),
.A2(n_42),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_58),
.C(n_64),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_43),
.A2(n_44),
.B1(n_64),
.B2(n_312),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_53),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_45),
.A2(n_164),
.B(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_52),
.B(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_46),
.A2(n_54),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_46),
.A2(n_54),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_47),
.B(n_51),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_49),
.A2(n_55),
.B1(n_145),
.B2(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_66),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_52),
.A2(n_54),
.B(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_53),
.A2(n_131),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_54),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_57),
.B(n_131),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_58),
.A2(n_59),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_64),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_64),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_68),
.B(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_68),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_65),
.A2(n_68),
.B1(n_105),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_65),
.A2(n_68),
.B1(n_133),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_65),
.A2(n_143),
.B(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_65),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_65),
.A2(n_68),
.B1(n_227),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_65),
.A2(n_247),
.B(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_68),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_68),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_68),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_69),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_74),
.B(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_74),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_75),
.A2(n_79),
.B1(n_80),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_75),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_330),
.B(n_336),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_302),
.A3(n_323),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_82)
);

AOI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_255),
.A3(n_277),
.B1(n_295),
.B2(n_301),
.C(n_342),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_214),
.C(n_251),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_185),
.B(n_213),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_158),
.B(n_184),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_138),
.B(n_157),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_126),
.B(n_137),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_112),
.B(n_125),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_100),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_95),
.B(n_155),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_118),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_107),
.B2(n_111),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_120),
.B(n_124),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_118),
.A2(n_119),
.B1(n_170),
.B2(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_118),
.A2(n_154),
.B(n_195),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_118),
.A2(n_119),
.B(n_153),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_128),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_139),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.CI(n_134),
.CON(n_129),
.SN(n_129)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_131),
.A2(n_164),
.B1(n_166),
.B2(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_135),
.B(n_171),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_136),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_149),
.B2(n_156),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_144),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_148),
.C(n_156),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_160),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_176),
.B2(n_177),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_179),
.C(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_175),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_164),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_173),
.C(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_180),
.B(n_228),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_187),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_199),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_198),
.C(n_199),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_209),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_206),
.B2(n_207),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_206),
.C(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_204),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_233),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_215),
.B(n_233),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_224),
.C(n_231),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_219),
.C(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_225),
.B1(n_231),
.B2(n_232),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_230),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_244),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_244),
.C(n_248),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_238),
.C(n_242),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_243),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_256),
.A2(n_296),
.B(n_300),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_257),
.B(n_258),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_269),
.B2(n_270),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_270),
.C(n_276),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_264),
.C(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_267),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_275),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_272),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_271),
.A2(n_284),
.B(n_287),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_278),
.B(n_279),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_279),
.Y(n_324)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.CI(n_294),
.CON(n_279),
.SN(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_292),
.B(n_293),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_292),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_293),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_293),
.A2(n_304),
.B1(n_314),
.B2(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B(n_299),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_316),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_314),
.C(n_315),
.Y(n_303)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_306),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_312),
.C(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_318),
.C(n_322),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_309),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule