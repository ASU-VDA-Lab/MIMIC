module fake_jpeg_28219_n_106 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_15),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_40),
.B1(n_20),
.B2(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_58),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_44),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_9),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_20),
.B1(n_32),
.B2(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_42),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_41),
.B(n_1),
.Y(n_63)
);

AOI21x1_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_0),
.B(n_3),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_32),
.B1(n_24),
.B2(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_24),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_68),
.B(n_74),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_29),
.B(n_32),
.C(n_31),
.D(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_73),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_24),
.C(n_9),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.C(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_11),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_29),
.C(n_14),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_29),
.C(n_14),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_63),
.C(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_59),
.B(n_65),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_85),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_72),
.B1(n_76),
.B2(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_82),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_16),
.B1(n_18),
.B2(n_7),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_86),
.B1(n_85),
.B2(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_3),
.C(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_96),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_92),
.C(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_82),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_7),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_87),
.B1(n_101),
.B2(n_100),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_103),
.Y(n_106)
);


endmodule