module fake_jpeg_19125_n_201 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_43),
.Y(n_59)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_51),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_23),
.B1(n_27),
.B2(n_34),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_31),
.C(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_57),
.B(n_9),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_22),
.B1(n_18),
.B2(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_22),
.B1(n_34),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_36),
.B1(n_24),
.B2(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_24),
.B1(n_32),
.B2(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_72),
.B1(n_29),
.B2(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_7),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_29),
.B1(n_28),
.B2(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_86),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_51),
.A3(n_49),
.B1(n_42),
.B2(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_68),
.Y(n_107)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_54),
.B1(n_26),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_31),
.B1(n_4),
.B2(n_6),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_31),
.B1(n_6),
.B2(n_7),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_12),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_12),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_106),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_65),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_81),
.B1(n_83),
.B2(n_76),
.Y(n_127)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_76),
.B1(n_71),
.B2(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_65),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_79),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_104),
.B1(n_81),
.B2(n_115),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_134),
.B1(n_115),
.B2(n_112),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_106),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_114),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_118),
.B1(n_108),
.B2(n_116),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_74),
.B(n_61),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_145),
.B1(n_135),
.B2(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_146),
.B1(n_129),
.B2(n_128),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_114),
.B(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_108),
.B1(n_100),
.B2(n_109),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_88),
.B1(n_91),
.B2(n_90),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_149),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_117),
.B1(n_89),
.B2(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_148),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_156),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_158),
.B1(n_140),
.B2(n_146),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_147),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_149),
.B(n_145),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_134),
.B1(n_136),
.B2(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_148),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_139),
.B1(n_148),
.B2(n_131),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_154),
.B1(n_160),
.B2(n_89),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_82),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_148),
.C(n_133),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_162),
.C(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_117),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_155),
.B(n_154),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_10),
.B(n_14),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_177),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_167),
.B1(n_170),
.B2(n_173),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_160),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_86),
.B(n_82),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_79),
.B(n_77),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_92),
.C(n_74),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.C(n_75),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_183),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_164),
.B1(n_163),
.B2(n_92),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_185),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_174),
.B(n_178),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_180),
.Y(n_194)
);

OAI321xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_179),
.A3(n_187),
.B1(n_175),
.B2(n_177),
.C(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_186),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_190),
.B(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_181),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_197),
.C(n_15),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_15),
.Y(n_201)
);


endmodule