module real_aes_18464_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_501;
wire n_488;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_948;
wire n_700;
wire n_399;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1699;
wire n_419;
wire n_730;
wire n_1023;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1802;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g556 ( .A(n_0), .Y(n_556) );
AO22x1_ASAP7_75t_L g608 ( .A1(n_0), .A2(n_234), .B1(n_609), .B2(n_611), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_1), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g396 ( .A(n_1), .Y(n_396) );
AND2x2_ASAP7_75t_L g540 ( .A(n_1), .B(n_497), .Y(n_540) );
AND2x2_ASAP7_75t_L g617 ( .A(n_1), .B(n_253), .Y(n_617) );
INVx1_ASAP7_75t_L g568 ( .A(n_2), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_2), .A2(n_128), .B1(n_513), .B2(n_606), .Y(n_605) );
XOR2x2_ASAP7_75t_L g347 ( .A(n_3), .B(n_348), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g1494 ( .A1(n_3), .A2(n_59), .B1(n_1477), .B2(n_1495), .Y(n_1494) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_4), .Y(n_1419) );
INVx1_ASAP7_75t_L g1282 ( .A(n_5), .Y(n_1282) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_6), .A2(n_225), .B1(n_922), .B2(n_923), .Y(n_921) );
INVxp67_ASAP7_75t_SL g959 ( .A(n_6), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_7), .A2(n_298), .B1(n_696), .B2(n_706), .C(n_1294), .Y(n_1293) );
AOI22xp33_ASAP7_75t_SL g1310 ( .A1(n_7), .A2(n_318), .B1(n_782), .B2(n_791), .Y(n_1310) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_8), .Y(n_847) );
AND4x1_ASAP7_75t_L g895 ( .A(n_8), .B(n_849), .C(n_852), .D(n_877), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_9), .A2(n_282), .B1(n_1016), .B2(n_1125), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_9), .A2(n_82), .B1(n_606), .B2(n_862), .C(n_998), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_10), .A2(n_321), .B1(n_636), .B2(n_1097), .Y(n_1209) );
INVx1_ASAP7_75t_L g1226 ( .A(n_10), .Y(n_1226) );
INVx2_ASAP7_75t_L g406 ( .A(n_11), .Y(n_406) );
OAI22xp5_ASAP7_75t_SL g1040 ( .A1(n_12), .A2(n_278), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_12), .A2(n_278), .B1(n_825), .B2(n_826), .C(n_1056), .Y(n_1055) );
XNOR2x1_ASAP7_75t_L g1019 ( .A(n_13), .B(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_14), .A2(n_125), .B1(n_1429), .B2(n_1431), .Y(n_1428) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_14), .A2(n_169), .B1(n_649), .B2(n_1189), .Y(n_1444) );
INVx1_ASAP7_75t_L g1245 ( .A(n_15), .Y(n_1245) );
OAI222xp33_ASAP7_75t_L g1267 ( .A1(n_15), .A2(n_171), .B1(n_867), .B2(n_1142), .C1(n_1268), .C2(n_1272), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_16), .A2(n_229), .B1(n_782), .B2(n_1122), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_16), .A2(n_141), .B1(n_1133), .B2(n_1135), .Y(n_1132) );
INVx1_ASAP7_75t_L g750 ( .A(n_17), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_18), .A2(n_265), .B1(n_944), .B2(n_1198), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_18), .A2(n_260), .B1(n_588), .B2(n_775), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_19), .A2(n_165), .B1(n_643), .B2(n_799), .Y(n_851) );
OAI211xp5_ASAP7_75t_L g853 ( .A1(n_19), .A2(n_803), .B(n_854), .C(n_858), .Y(n_853) );
OAI22xp33_ASAP7_75t_L g1439 ( .A1(n_20), .A2(n_211), .B1(n_787), .B2(n_788), .Y(n_1439) );
INVx1_ASAP7_75t_L g1446 ( .A(n_20), .Y(n_1446) );
AOI22xp33_ASAP7_75t_SL g1435 ( .A1(n_21), .A2(n_88), .B1(n_925), .B2(n_1125), .Y(n_1435) );
AOI22xp33_ASAP7_75t_SL g1452 ( .A1(n_21), .A2(n_243), .B1(n_1134), .B2(n_1135), .Y(n_1452) );
AOI22xp5_ASAP7_75t_L g1504 ( .A1(n_22), .A2(n_221), .B1(n_1484), .B2(n_1487), .Y(n_1504) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_23), .A2(n_299), .B1(n_643), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_24), .A2(n_90), .B1(n_609), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_24), .A2(n_36), .B1(n_885), .B2(n_886), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g1155 ( .A(n_25), .Y(n_1155) );
INVx1_ASAP7_75t_L g1054 ( .A(n_26), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1465 ( .A(n_27), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_27), .B(n_1463), .Y(n_1478) );
AOI22xp5_ASAP7_75t_L g1493 ( .A1(n_28), .A2(n_194), .B1(n_1484), .B2(n_1487), .Y(n_1493) );
OAI22xp5_ASAP7_75t_SL g693 ( .A1(n_29), .A2(n_283), .B1(n_353), .B2(n_379), .Y(n_693) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_29), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_30), .A2(n_222), .B1(n_777), .B2(n_782), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_30), .A2(n_311), .B1(n_836), .B2(n_839), .C(n_840), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_31), .Y(n_899) );
INVx1_ASAP7_75t_L g974 ( .A(n_32), .Y(n_974) );
OAI211xp5_ASAP7_75t_L g983 ( .A1(n_32), .A2(n_947), .B(n_984), .C(n_990), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_33), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_34), .A2(n_318), .B1(n_636), .B2(n_1198), .Y(n_1299) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_34), .A2(n_298), .B1(n_782), .B2(n_1251), .Y(n_1311) );
AOI22xp5_ASAP7_75t_L g1529 ( .A1(n_35), .A2(n_273), .B1(n_1484), .B2(n_1487), .Y(n_1529) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_36), .A2(n_327), .B1(n_606), .B2(n_840), .C(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_37), .A2(n_53), .B1(n_575), .B2(n_660), .Y(n_1396) );
INVx1_ASAP7_75t_L g1406 ( .A(n_37), .Y(n_1406) );
INVx1_ASAP7_75t_L g771 ( .A(n_38), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_38), .A2(n_247), .B1(n_823), .B2(n_826), .C(n_829), .Y(n_822) );
INVx1_ASAP7_75t_L g1337 ( .A(n_39), .Y(n_1337) );
INVx1_ASAP7_75t_L g1265 ( .A(n_40), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_41), .A2(n_50), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_41), .A2(n_163), .B1(n_782), .B2(n_889), .Y(n_1353) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_42), .A2(n_301), .B1(n_606), .B2(n_706), .C(n_998), .Y(n_997) );
INVxp67_ASAP7_75t_SL g1006 ( .A(n_42), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g1500 ( .A1(n_43), .A2(n_122), .B1(n_1484), .B2(n_1487), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1744 ( .A1(n_43), .A2(n_1745), .B1(n_1748), .B2(n_1799), .Y(n_1744) );
OAI22xp5_ASAP7_75t_L g1750 ( .A1(n_43), .A2(n_1751), .B1(n_1752), .B2(n_1753), .Y(n_1750) );
INVx1_ASAP7_75t_L g1751 ( .A(n_43), .Y(n_1751) );
INVx1_ASAP7_75t_L g980 ( .A(n_44), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_44), .A2(n_213), .B1(n_803), .B2(n_1000), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1387 ( .A1(n_45), .A2(n_336), .B1(n_462), .B2(n_1388), .C(n_1389), .Y(n_1387) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_45), .A2(n_123), .B1(n_696), .B2(n_1101), .C(n_1405), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_46), .A2(n_277), .B1(n_916), .B2(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g950 ( .A(n_46), .Y(n_950) );
INVx1_ASAP7_75t_L g1212 ( .A(n_47), .Y(n_1212) );
OAI21xp5_ASAP7_75t_L g1303 ( .A1(n_48), .A2(n_1025), .B(n_1304), .Y(n_1303) );
AOI22xp5_ASAP7_75t_L g1498 ( .A1(n_49), .A2(n_174), .B1(n_1477), .B2(n_1499), .Y(n_1498) );
AOI22xp33_ASAP7_75t_SL g1346 ( .A1(n_50), .A2(n_176), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
INVx1_ASAP7_75t_L g1211 ( .A(n_51), .Y(n_1211) );
INVx1_ASAP7_75t_L g1264 ( .A(n_52), .Y(n_1264) );
INVx1_ASAP7_75t_L g1401 ( .A(n_53), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g1772 ( .A1(n_54), .A2(n_197), .B1(n_649), .B2(n_709), .Y(n_1772) );
INVx1_ASAP7_75t_L g1797 ( .A(n_54), .Y(n_1797) );
INVxp67_ASAP7_75t_SL g996 ( .A(n_55), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_55), .A2(n_139), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
INVxp67_ASAP7_75t_L g1417 ( .A(n_56), .Y(n_1417) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_57), .Y(n_355) );
INVx1_ASAP7_75t_L g855 ( .A(n_58), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_58), .A2(n_105), .B1(n_753), .B2(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g908 ( .A(n_60), .Y(n_908) );
INVx1_ASAP7_75t_L g1115 ( .A(n_61), .Y(n_1115) );
OAI222xp33_ASAP7_75t_L g1141 ( .A1(n_61), .A2(n_342), .B1(n_866), .B2(n_1142), .C1(n_1143), .C2(n_1148), .Y(n_1141) );
INVx1_ASAP7_75t_L g1053 ( .A(n_62), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1774 ( .A1(n_63), .A2(n_232), .B1(n_808), .B2(n_1134), .Y(n_1774) );
INVx1_ASAP7_75t_L g1791 ( .A(n_63), .Y(n_1791) );
AOI22xp33_ASAP7_75t_L g1608 ( .A1(n_64), .A2(n_245), .B1(n_1477), .B2(n_1495), .Y(n_1608) );
CKINVDCx5p33_ASAP7_75t_R g1140 ( .A(n_65), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1705 ( .A1(n_66), .A2(n_240), .B1(n_434), .B2(n_782), .Y(n_1705) );
AOI221xp5_ASAP7_75t_L g1717 ( .A1(n_66), .A2(n_172), .B1(n_513), .B2(n_606), .C(n_706), .Y(n_1717) );
AOI22xp33_ASAP7_75t_L g1704 ( .A1(n_67), .A2(n_172), .B1(n_782), .B2(n_916), .Y(n_1704) );
AOI22xp33_ASAP7_75t_L g1718 ( .A1(n_67), .A2(n_240), .B1(n_609), .B2(n_636), .Y(n_1718) );
INVx1_ASAP7_75t_L g376 ( .A(n_68), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_69), .A2(n_326), .B1(n_836), .B2(n_860), .C(n_862), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_69), .A2(n_292), .B1(n_889), .B2(n_890), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_70), .A2(n_1284), .B1(n_1285), .B2(n_1314), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_70), .Y(n_1314) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_71), .A2(n_323), .B1(n_630), .B2(n_1324), .C(n_1325), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_71), .A2(n_286), .B1(n_914), .B2(n_1351), .C(n_1352), .Y(n_1350) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_72), .A2(n_177), .B1(n_912), .B2(n_914), .Y(n_911) );
INVxp67_ASAP7_75t_SL g956 ( .A(n_72), .Y(n_956) );
OAI211xp5_ASAP7_75t_SL g1379 ( .A1(n_73), .A2(n_579), .B(n_1362), .C(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1409 ( .A(n_73), .Y(n_1409) );
INVx1_ASAP7_75t_L g1291 ( .A(n_74), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_75), .A2(n_252), .B1(n_451), .B2(n_455), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_75), .A2(n_252), .B1(n_501), .B2(n_503), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g1709 ( .A(n_76), .Y(n_1709) );
INVxp67_ASAP7_75t_SL g1342 ( .A(n_77), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_77), .A2(n_331), .B1(n_1355), .B2(n_1358), .Y(n_1354) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_78), .A2(n_337), .B1(n_775), .B2(n_784), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_78), .A2(n_145), .B1(n_700), .B2(n_810), .C(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g1292 ( .A(n_79), .Y(n_1292) );
OR2x2_ASAP7_75t_L g978 ( .A(n_80), .B(n_796), .Y(n_978) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_81), .A2(n_210), .B1(n_826), .B2(n_992), .C(n_993), .Y(n_991) );
OAI322xp33_ASAP7_75t_L g1004 ( .A1(n_81), .A2(n_437), .A3(n_734), .B1(n_788), .B2(n_1005), .C1(n_1007), .C2(n_1010), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_82), .A2(n_135), .B1(n_1016), .B2(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_83), .A2(n_175), .B1(n_1477), .B2(n_1484), .Y(n_1513) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_84), .A2(n_204), .B1(n_782), .B2(n_916), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_84), .A2(n_97), .B1(n_944), .B2(n_1097), .Y(n_1096) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_85), .A2(n_162), .B1(n_611), .B2(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_85), .Y(n_746) );
INVx1_ASAP7_75t_L g1023 ( .A(n_86), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_87), .A2(n_279), .B1(n_748), .B2(n_1033), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_87), .A2(n_99), .B1(n_700), .B2(n_813), .C(n_940), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1443 ( .A1(n_88), .A2(n_309), .B1(n_606), .B2(n_839), .C(n_989), .Y(n_1443) );
INVx1_ASAP7_75t_L g964 ( .A(n_89), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_90), .A2(n_327), .B1(n_885), .B2(n_886), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_91), .A2(n_293), .B1(n_1487), .B2(n_1495), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_92), .A2(n_271), .B1(n_775), .B2(n_1033), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1187 ( .A1(n_92), .A2(n_266), .B1(n_696), .B2(n_989), .C(n_1095), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1756 ( .A1(n_93), .A2(n_127), .B1(n_951), .B2(n_1722), .C(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1779 ( .A(n_93), .Y(n_1779) );
AOI22xp5_ASAP7_75t_L g1476 ( .A1(n_94), .A2(n_159), .B1(n_1477), .B2(n_1481), .Y(n_1476) );
OAI21xp33_ASAP7_75t_L g1151 ( .A1(n_95), .A2(n_1152), .B(n_1153), .Y(n_1151) );
INVx1_ASAP7_75t_L g1026 ( .A(n_96), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_97), .A2(n_281), .B1(n_782), .B2(n_916), .Y(n_1087) );
INVx1_ASAP7_75t_L g1174 ( .A(n_98), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_98), .A2(n_290), .B1(n_944), .B2(n_1189), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_99), .A2(n_191), .B1(n_914), .B2(n_1015), .Y(n_1039) );
INVx1_ASAP7_75t_L g1759 ( .A(n_100), .Y(n_1759) );
OAI221xp5_ASAP7_75t_SL g1783 ( .A1(n_100), .A2(n_126), .B1(n_436), .B2(n_595), .C(n_732), .Y(n_1783) );
INVx1_ASAP7_75t_L g370 ( .A(n_101), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_102), .A2(n_316), .B1(n_775), .B2(n_1033), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g1259 ( .A(n_102), .Y(n_1259) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_103), .Y(n_1080) );
XNOR2xp5_ASAP7_75t_L g1201 ( .A(n_104), .B(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g857 ( .A(n_105), .Y(n_857) );
OAI211xp5_ASAP7_75t_L g1721 ( .A1(n_106), .A2(n_1722), .B(n_1723), .C(n_1724), .Y(n_1721) );
INVx1_ASAP7_75t_L g1737 ( .A(n_106), .Y(n_1737) );
INVx1_ASAP7_75t_L g994 ( .A(n_107), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1609 ( .A1(n_108), .A2(n_320), .B1(n_1484), .B2(n_1487), .Y(n_1609) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_109), .A2(n_239), .B1(n_611), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_109), .A2(n_256), .B1(n_739), .B2(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g399 ( .A(n_110), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g1216 ( .A1(n_111), .A2(n_696), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1225 ( .A(n_111), .Y(n_1225) );
INVx1_ASAP7_75t_L g675 ( .A(n_112), .Y(n_675) );
INVx1_ASAP7_75t_L g1164 ( .A(n_113), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g865 ( .A1(n_114), .A2(n_268), .B1(n_823), .B2(n_866), .C(n_868), .Y(n_865) );
INVx1_ASAP7_75t_L g894 ( .A(n_114), .Y(n_894) );
INVx1_ASAP7_75t_L g1463 ( .A(n_115), .Y(n_1463) );
AOI221xp5_ASAP7_75t_L g1206 ( .A1(n_116), .A2(n_254), .B1(n_989), .B2(n_1101), .C(n_1207), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_116), .A2(n_181), .B1(n_763), .B2(n_775), .Y(n_1227) );
INVx1_ASAP7_75t_L g1075 ( .A(n_117), .Y(n_1075) );
INVx1_ASAP7_75t_L g1074 ( .A(n_118), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_119), .A2(n_280), .B1(n_925), .B2(n_1015), .C(n_1083), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1094 ( .A1(n_119), .A2(n_236), .B1(n_813), .B2(n_1066), .C(n_1095), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1773 ( .A1(n_120), .A2(n_155), .B1(n_813), .B2(n_998), .C(n_1770), .Y(n_1773) );
INVx1_ASAP7_75t_L g1787 ( .A(n_120), .Y(n_1787) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_121), .A2(n_185), .B1(n_916), .B2(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g954 ( .A(n_121), .Y(n_954) );
INVx1_ASAP7_75t_L g1394 ( .A(n_123), .Y(n_1394) );
OAI222xp33_ASAP7_75t_L g583 ( .A1(n_124), .A2(n_322), .B1(n_584), .B2(n_590), .C1(n_592), .C2(n_596), .Y(n_583) );
INVx1_ASAP7_75t_L g618 ( .A(n_124), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g1451 ( .A1(n_125), .A2(n_706), .B(n_838), .Y(n_1451) );
INVx1_ASAP7_75t_L g1765 ( .A(n_126), .Y(n_1765) );
INVx1_ASAP7_75t_L g1777 ( .A(n_127), .Y(n_1777) );
INVx1_ASAP7_75t_L g564 ( .A(n_128), .Y(n_564) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_129), .A2(n_682), .B(n_684), .C(n_686), .Y(n_681) );
INVxp33_ASAP7_75t_SL g720 ( .A(n_129), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_130), .Y(n_1179) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_131), .A2(n_170), .B1(n_549), .B2(n_1366), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g1368 ( .A(n_131), .Y(n_1368) );
INVx1_ASAP7_75t_L g1297 ( .A(n_132), .Y(n_1297) );
INVx1_ASAP7_75t_L g1763 ( .A(n_133), .Y(n_1763) );
OAI21xp33_ASAP7_75t_L g1781 ( .A1(n_133), .A2(n_722), .B(n_1782), .Y(n_1781) );
AOI22xp33_ASAP7_75t_SL g1528 ( .A1(n_134), .A2(n_215), .B1(n_1477), .B2(n_1495), .Y(n_1528) );
INVx1_ASAP7_75t_L g1146 ( .A(n_135), .Y(n_1146) );
INVx1_ASAP7_75t_L g1170 ( .A(n_136), .Y(n_1170) );
AOI21xp33_ASAP7_75t_L g1196 ( .A1(n_136), .A2(n_696), .B(n_840), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_137), .A2(n_168), .B1(n_643), .B2(n_1025), .Y(n_1165) );
OAI211xp5_ASAP7_75t_L g1185 ( .A1(n_137), .A2(n_1129), .B(n_1186), .C(n_1190), .Y(n_1185) );
INVx1_ASAP7_75t_L g903 ( .A(n_138), .Y(n_903) );
OAI222xp33_ASAP7_75t_L g946 ( .A1(n_138), .A2(n_207), .B1(n_866), .B2(n_947), .C1(n_948), .C2(n_955), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_139), .A2(n_223), .B1(n_606), .B2(n_700), .C(n_989), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_140), .A2(n_260), .B1(n_813), .B2(n_1066), .C(n_1101), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_140), .A2(n_265), .B1(n_763), .B2(n_775), .Y(n_1309) );
AOI22xp33_ASAP7_75t_SL g1120 ( .A1(n_141), .A2(n_233), .B1(n_782), .B2(n_922), .Y(n_1120) );
OAI22xp33_ASAP7_75t_L g1378 ( .A1(n_142), .A2(n_341), .B1(n_549), .B2(n_1366), .Y(n_1378) );
INVxp33_ASAP7_75t_SL g1413 ( .A(n_142), .Y(n_1413) );
AOI22xp5_ASAP7_75t_L g1698 ( .A1(n_143), .A2(n_1699), .B1(n_1738), .B2(n_1739), .Y(n_1698) );
CKINVDCx5p33_ASAP7_75t_R g1738 ( .A(n_143), .Y(n_1738) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_144), .Y(n_1381) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_145), .A2(n_192), .B1(n_740), .B2(n_775), .Y(n_774) );
OA21x2_ASAP7_75t_L g1021 ( .A1(n_146), .A2(n_796), .B(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1385 ( .A(n_147), .Y(n_1385) );
AOI221xp5_ASAP7_75t_L g1399 ( .A1(n_147), .A2(n_248), .B1(n_696), .B2(n_1101), .C(n_1400), .Y(n_1399) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_148), .A2(n_163), .B1(n_1322), .B2(n_1328), .C(n_1329), .Y(n_1327) );
AOI221xp5_ASAP7_75t_L g1349 ( .A1(n_148), .A2(n_323), .B1(n_578), .B2(n_740), .C(n_775), .Y(n_1349) );
AOI221xp5_ASAP7_75t_SL g1769 ( .A1(n_149), .A2(n_306), .B1(n_706), .B2(n_998), .C(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1794 ( .A(n_149), .Y(n_1794) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_150), .A2(n_311), .B1(n_777), .B2(n_779), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_150), .A2(n_222), .B1(n_807), .B2(n_808), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g1767 ( .A(n_151), .Y(n_1767) );
INVx1_ASAP7_75t_L g1287 ( .A(n_152), .Y(n_1287) );
INVx1_ASAP7_75t_L g930 ( .A(n_153), .Y(n_930) );
INVx1_ASAP7_75t_L g1422 ( .A(n_154), .Y(n_1422) );
OAI221xp5_ASAP7_75t_SL g1448 ( .A1(n_154), .A2(n_258), .B1(n_823), .B2(n_866), .C(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1798 ( .A(n_155), .Y(n_1798) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_156), .Y(n_797) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_157), .A2(n_164), .B1(n_476), .B2(n_479), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_157), .A2(n_164), .B1(n_488), .B2(n_494), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g1213 ( .A1(n_158), .A2(n_333), .B1(n_867), .B2(n_1142), .C(n_1214), .Y(n_1213) );
OAI22xp33_ASAP7_75t_L g1232 ( .A1(n_158), .A2(n_333), .B1(n_728), .B2(n_1042), .Y(n_1232) );
INVx1_ASAP7_75t_L g1156 ( .A(n_159), .Y(n_1156) );
INVx1_ASAP7_75t_L g1733 ( .A(n_160), .Y(n_1733) );
INVx1_ASAP7_75t_L g465 ( .A(n_161), .Y(n_465) );
INVx1_ASAP7_75t_L g737 ( .A(n_162), .Y(n_737) );
INVx1_ASAP7_75t_L g386 ( .A(n_166), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_167), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_169), .A2(n_302), .B1(n_1431), .B2(n_1433), .Y(n_1432) );
INVxp67_ASAP7_75t_SL g1336 ( .A(n_170), .Y(n_1336) );
INVx1_ASAP7_75t_L g1244 ( .A(n_171), .Y(n_1244) );
INVx1_ASAP7_75t_L g558 ( .A(n_173), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_173), .A2(n_262), .B1(n_609), .B2(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g1330 ( .A(n_176), .Y(n_1330) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_177), .A2(n_225), .B1(n_862), .B2(n_936), .C(n_939), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_178), .Y(n_687) );
INVx1_ASAP7_75t_L g702 ( .A(n_179), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g1204 ( .A1(n_180), .A2(n_1129), .B(n_1205), .C(n_1210), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_180), .A2(n_325), .B1(n_643), .B2(n_1025), .Y(n_1235) );
AOI22xp33_ASAP7_75t_SL g1218 ( .A1(n_181), .A2(n_305), .B1(n_611), .B2(n_1198), .Y(n_1218) );
INVx1_ASAP7_75t_L g1031 ( .A(n_182), .Y(n_1031) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_182), .A2(n_228), .B1(n_1063), .B2(n_1066), .C(n_1067), .Y(n_1062) );
OAI211xp5_ASAP7_75t_L g1713 ( .A1(n_183), .A2(n_1714), .B(n_1715), .C(n_1720), .Y(n_1713) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_183), .B(n_760), .Y(n_1728) );
XNOR2x2_ASAP7_75t_L g765 ( .A(n_184), .B(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_185), .A2(n_277), .B1(n_807), .B2(n_942), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g1085 ( .A1(n_186), .A2(n_236), .B1(n_914), .B2(n_1015), .C(n_1086), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_186), .A2(n_280), .B1(n_698), .B2(n_944), .Y(n_1099) );
INVx2_ASAP7_75t_L g1480 ( .A(n_187), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_187), .B(n_291), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_187), .B(n_1486), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_188), .A2(n_335), .B1(n_779), .B2(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1271 ( .A(n_188), .Y(n_1271) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_189), .Y(n_1003) );
INVx1_ASAP7_75t_L g1192 ( .A(n_190), .Y(n_1192) );
INVx1_ASAP7_75t_L g1061 ( .A(n_191), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g831 ( .A(n_192), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g1506 ( .A1(n_193), .A2(n_251), .B1(n_1477), .B2(n_1487), .Y(n_1506) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_195), .A2(n_264), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g816 ( .A(n_195), .Y(n_816) );
INVx1_ASAP7_75t_L g1438 ( .A(n_196), .Y(n_1438) );
INVx1_ASAP7_75t_L g1786 ( .A(n_197), .Y(n_1786) );
INVx1_ASAP7_75t_L g652 ( .A(n_198), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g1507 ( .A1(n_199), .A2(n_205), .B1(n_1481), .B2(n_1484), .Y(n_1507) );
INVx1_ASAP7_75t_L g928 ( .A(n_200), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g1706 ( .A1(n_201), .A2(n_289), .B1(n_588), .B2(n_775), .Y(n_1706) );
AOI22xp33_ASAP7_75t_L g1716 ( .A1(n_201), .A2(n_275), .B1(n_636), .B2(n_709), .Y(n_1716) );
AOI22xp33_ASAP7_75t_SL g1175 ( .A1(n_202), .A2(n_266), .B1(n_775), .B2(n_1033), .Y(n_1175) );
AOI22xp33_ASAP7_75t_SL g1197 ( .A1(n_202), .A2(n_271), .B1(n_864), .B2(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1281 ( .A(n_203), .Y(n_1281) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_204), .A2(n_281), .B1(n_840), .B2(n_1066), .C(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1038 ( .A(n_206), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_206), .A2(n_270), .B1(n_636), .B2(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g905 ( .A(n_207), .Y(n_905) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_208), .A2(n_435), .B(n_460), .C(n_464), .Y(n_459) );
INVx1_ASAP7_75t_L g519 ( .A(n_208), .Y(n_519) );
INVx1_ASAP7_75t_L g1118 ( .A(n_209), .Y(n_1118) );
OAI211xp5_ASAP7_75t_L g1128 ( .A1(n_209), .A2(n_1129), .B(n_1130), .C(n_1137), .Y(n_1128) );
INVx1_ASAP7_75t_L g973 ( .A(n_210), .Y(n_973) );
INVx1_ASAP7_75t_L g1447 ( .A(n_211), .Y(n_1447) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_212), .Y(n_561) );
INVx1_ASAP7_75t_L g976 ( .A(n_213), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g1215 ( .A(n_214), .Y(n_1215) );
INVx1_ASAP7_75t_L g1017 ( .A(n_215), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g1725 ( .A(n_216), .Y(n_1725) );
INVx2_ASAP7_75t_L g405 ( .A(n_217), .Y(n_405) );
INVx1_ASAP7_75t_L g444 ( .A(n_217), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_217), .B(n_406), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_218), .Y(n_1138) );
AOI22xp5_ASAP7_75t_L g1483 ( .A1(n_219), .A2(n_332), .B1(n_1484), .B2(n_1487), .Y(n_1483) );
INVx1_ASAP7_75t_L g573 ( .A(n_220), .Y(n_573) );
NAND2xp33_ASAP7_75t_SL g637 ( .A(n_220), .B(n_513), .Y(n_637) );
INVx1_ASAP7_75t_L g1008 ( .A(n_223), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_224), .A2(n_307), .B1(n_424), .B2(n_917), .Y(n_1252) );
INVx1_ASAP7_75t_L g1269 ( .A(n_224), .Y(n_1269) );
AOI22xp33_ASAP7_75t_SL g1249 ( .A1(n_226), .A2(n_250), .B1(n_775), .B2(n_890), .Y(n_1249) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_226), .Y(n_1273) );
INVx1_ASAP7_75t_L g398 ( .A(n_227), .Y(n_398) );
INVx1_ASAP7_75t_L g1037 ( .A(n_228), .Y(n_1037) );
INVx1_ASAP7_75t_L g1145 ( .A(n_229), .Y(n_1145) );
INVx1_ASAP7_75t_L g987 ( .A(n_230), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g1726 ( .A1(n_231), .A2(n_296), .B1(n_1722), .B2(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1736 ( .A(n_231), .Y(n_1736) );
INVx1_ASAP7_75t_L g1795 ( .A(n_232), .Y(n_1795) );
INVx1_ASAP7_75t_L g1149 ( .A(n_233), .Y(n_1149) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_234), .A2(n_575), .B(n_578), .Y(n_574) );
INVx1_ASAP7_75t_L g641 ( .A(n_235), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g1278 ( .A1(n_237), .A2(n_1025), .B(n_1279), .Y(n_1278) );
BUFx3_ASAP7_75t_L g411 ( .A(n_238), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_239), .A2(n_272), .B1(n_740), .B2(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g1092 ( .A(n_241), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_242), .Y(n_1382) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_243), .A2(n_309), .B1(n_923), .B2(n_1125), .Y(n_1427) );
INVx1_ASAP7_75t_L g543 ( .A(n_244), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_244), .B(n_549), .Y(n_548) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_246), .A2(n_696), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g736 ( .A(n_246), .Y(n_736) );
INVx1_ASAP7_75t_L g770 ( .A(n_247), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g1395 ( .A1(n_248), .A2(n_563), .B(n_1352), .Y(n_1395) );
XOR2x2_ASAP7_75t_L g670 ( .A(n_249), .B(n_671), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g1261 ( .A1(n_250), .A2(n_813), .B(n_940), .Y(n_1261) );
BUFx3_ASAP7_75t_L g368 ( .A(n_253), .Y(n_368) );
INVx1_ASAP7_75t_L g497 ( .A(n_253), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_254), .A2(n_305), .B1(n_775), .B2(n_914), .Y(n_1231) );
XNOR2x1_ASAP7_75t_L g1071 ( .A(n_255), .B(n_1072), .Y(n_1071) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_256), .B(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_SL g1425 ( .A(n_257), .Y(n_1425) );
OAI211xp5_ASAP7_75t_SL g1441 ( .A1(n_257), .A2(n_803), .B(n_1442), .C(n_1445), .Y(n_1441) );
INVx1_ASAP7_75t_L g1423 ( .A(n_258), .Y(n_1423) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_259), .Y(n_1386) );
CKINVDCx5p33_ASAP7_75t_R g1758 ( .A(n_261), .Y(n_1758) );
INVx1_ASAP7_75t_L g569 ( .A(n_262), .Y(n_569) );
INVx1_ASAP7_75t_L g1091 ( .A(n_263), .Y(n_1091) );
INVx1_ASAP7_75t_L g819 ( .A(n_264), .Y(n_819) );
INVx1_ASAP7_75t_L g985 ( .A(n_267), .Y(n_985) );
INVx1_ASAP7_75t_L g892 ( .A(n_268), .Y(n_892) );
INVx1_ASAP7_75t_L g1191 ( .A(n_269), .Y(n_1191) );
NAND2xp33_ASAP7_75t_SL g1034 ( .A(n_270), .B(n_917), .Y(n_1034) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_272), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g1369 ( .A(n_274), .Y(n_1369) );
AOI22xp33_ASAP7_75t_SL g1703 ( .A1(n_275), .A2(n_343), .B1(n_775), .B2(n_1033), .Y(n_1703) );
INVx1_ASAP7_75t_L g413 ( .A(n_276), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_276), .Y(n_420) );
INVx1_ASAP7_75t_L g1058 ( .A(n_279), .Y(n_1058) );
INVx1_ASAP7_75t_L g1150 ( .A(n_282), .Y(n_1150) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_283), .A2(n_714), .B(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g1247 ( .A(n_284), .Y(n_1247) );
AOI22xp5_ASAP7_75t_SL g1503 ( .A1(n_285), .A2(n_339), .B1(n_1477), .B2(n_1481), .Y(n_1503) );
INVx1_ASAP7_75t_L g1331 ( .A(n_286), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_287), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_288), .Y(n_1078) );
AOI221xp5_ASAP7_75t_SL g1719 ( .A1(n_289), .A2(n_343), .B1(n_513), .B2(n_813), .C(n_838), .Y(n_1719) );
INVx1_ASAP7_75t_L g1181 ( .A(n_290), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_291), .B(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1486 ( .A(n_291), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_292), .Y(n_873) );
INVx1_ASAP7_75t_L g471 ( .A(n_294), .Y(n_471) );
OAI211xp5_ASAP7_75t_L g509 ( .A1(n_294), .A2(n_360), .B(n_510), .C(n_515), .Y(n_509) );
INVx1_ASAP7_75t_L g1302 ( .A(n_295), .Y(n_1302) );
INVx1_ASAP7_75t_L g1710 ( .A(n_296), .Y(n_1710) );
XNOR2xp5_ASAP7_75t_L g1370 ( .A(n_297), .B(n_1371), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g802 ( .A1(n_299), .A2(n_803), .B(n_805), .C(n_815), .Y(n_802) );
INVx1_ASAP7_75t_L g352 ( .A(n_300), .Y(n_352) );
INVxp67_ASAP7_75t_SL g1012 ( .A(n_301), .Y(n_1012) );
INVx1_ASAP7_75t_L g1450 ( .A(n_302), .Y(n_1450) );
INVx1_ASAP7_75t_L g1301 ( .A(n_303), .Y(n_1301) );
CKINVDCx16_ASAP7_75t_R g587 ( .A(n_304), .Y(n_587) );
INVx1_ASAP7_75t_L g1789 ( .A(n_306), .Y(n_1789) );
AOI22xp5_ASAP7_75t_L g1262 ( .A1(n_307), .A2(n_335), .B1(n_698), .B2(n_944), .Y(n_1262) );
OAI21xp33_ASAP7_75t_L g926 ( .A1(n_308), .A2(n_799), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1373 ( .A(n_310), .Y(n_1373) );
OAI21xp5_ASAP7_75t_SL g1103 ( .A1(n_312), .A2(n_1025), .B(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1392 ( .A(n_313), .Y(n_1392) );
INVx1_ASAP7_75t_L g385 ( .A(n_314), .Y(n_385) );
INVx1_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
INVxp67_ASAP7_75t_SL g1276 ( .A(n_316), .Y(n_1276) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_317), .Y(n_869) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_317), .A2(n_326), .B1(n_739), .B2(n_883), .Y(n_882) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_319), .Y(n_357) );
INVx1_ASAP7_75t_L g1230 ( .A(n_321), .Y(n_1230) );
NOR2xp33_ASAP7_75t_R g625 ( .A(n_322), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g532 ( .A(n_324), .Y(n_532) );
INVxp67_ASAP7_75t_SL g1340 ( .A(n_328), .Y(n_1340) );
OAI221xp5_ASAP7_75t_L g1364 ( .A1(n_328), .A2(n_330), .B1(n_579), .B2(n_592), .C(n_596), .Y(n_1364) );
INVx1_ASAP7_75t_L g1234 ( .A(n_329), .Y(n_1234) );
OAI221xp5_ASAP7_75t_L g1326 ( .A1(n_330), .A2(n_331), .B1(n_615), .B2(n_620), .C(n_638), .Y(n_1326) );
INVx2_ASAP7_75t_L g366 ( .A(n_334), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_334), .Y(n_394) );
INVx1_ASAP7_75t_L g443 ( .A(n_334), .Y(n_443) );
INVx1_ASAP7_75t_L g1402 ( .A(n_336), .Y(n_1402) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_337), .Y(n_834) );
OAI22xp33_ASAP7_75t_SL g1183 ( .A1(n_338), .A2(n_340), .B1(n_728), .B2(n_1042), .Y(n_1183) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_338), .A2(n_340), .B1(n_823), .B2(n_867), .C(n_1194), .Y(n_1193) );
XNOR2xp5_ASAP7_75t_L g1161 ( .A(n_339), .B(n_1162), .Y(n_1161) );
INVxp67_ASAP7_75t_SL g1376 ( .A(n_341), .Y(n_1376) );
INVx1_ASAP7_75t_L g1114 ( .A(n_342), .Y(n_1114) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_1458), .B(n_1469), .Y(n_344) );
XNOR2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_663), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_530), .B1(n_661), .B2(n_662), .Y(n_346) );
INVx1_ASAP7_75t_L g661 ( .A(n_347), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_449), .C(n_486), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_400), .Y(n_349) );
OAI33xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_363), .A3(n_369), .B1(n_384), .B2(n_387), .B3(n_397), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_358), .B2(n_359), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_352), .A2(n_385), .B1(n_423), .B2(n_428), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_353), .A2(n_377), .B1(n_398), .B2(n_399), .Y(n_397) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g634 ( .A(n_354), .Y(n_634) );
BUFx2_ASAP7_75t_L g953 ( .A(n_354), .Y(n_953) );
BUFx3_ASAP7_75t_L g1270 ( .A(n_354), .Y(n_1270) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_355), .B(n_357), .Y(n_362) );
OR2x2_ASAP7_75t_L g375 ( .A(n_355), .B(n_357), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_355), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g499 ( .A(n_355), .Y(n_499) );
AND2x2_ASAP7_75t_L g514 ( .A(n_355), .B(n_357), .Y(n_514) );
BUFx2_ASAP7_75t_L g518 ( .A(n_355), .Y(n_518) );
INVx1_ASAP7_75t_L g542 ( .A(n_355), .Y(n_542) );
AND2x2_ASAP7_75t_L g612 ( .A(n_355), .B(n_383), .Y(n_612) );
AND2x2_ASAP7_75t_L g541 ( .A(n_356), .B(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_356), .Y(n_691) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g383 ( .A(n_357), .Y(n_383) );
AND2x2_ASAP7_75t_L g498 ( .A(n_357), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g524 ( .A(n_357), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_358), .A2(n_386), .B1(n_433), .B2(n_435), .Y(n_432) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_360), .A2(n_371), .B1(n_385), .B2(n_386), .Y(n_384) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x6_ASAP7_75t_L g638 ( .A(n_361), .B(n_639), .Y(n_638) );
INVx4_ASAP7_75t_L g685 ( .A(n_361), .Y(n_685) );
BUFx4f_ASAP7_75t_L g949 ( .A(n_361), .Y(n_949) );
BUFx4f_ASAP7_75t_L g1260 ( .A(n_361), .Y(n_1260) );
BUFx4f_ASAP7_75t_L g1727 ( .A(n_361), .Y(n_1727) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g627 ( .A(n_362), .Y(n_627) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_364), .B(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g1329 ( .A1(n_364), .A2(n_949), .B1(n_1270), .B2(n_1330), .C(n_1331), .Y(n_1329) );
HB1xp67_ASAP7_75t_L g1403 ( .A(n_364), .Y(n_1403) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g658 ( .A(n_365), .Y(n_658) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_365), .B(n_578), .Y(n_1083) );
OR2x6_ASAP7_75t_L g1255 ( .A(n_365), .B(n_578), .Y(n_1255) );
BUFx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g600 ( .A(n_366), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_366), .B(n_617), .Y(n_622) );
AND2x4_ASAP7_75t_L g395 ( .A(n_368), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g493 ( .A(n_368), .Y(n_493) );
BUFx2_ASAP7_75t_L g508 ( .A(n_368), .Y(n_508) );
AND2x4_ASAP7_75t_L g522 ( .A(n_368), .B(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_376), .B2(n_377), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_370), .A2(n_398), .B1(n_408), .B2(n_414), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_371), .A2(n_869), .B1(n_870), .B2(n_873), .C(n_874), .Y(n_868) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g830 ( .A(n_373), .Y(n_830) );
BUFx3_ASAP7_75t_L g1057 ( .A(n_373), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_373), .A2(n_1277), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
OAI22x1_ASAP7_75t_SL g1405 ( .A1(n_373), .A2(n_1277), .B1(n_1386), .B2(n_1406), .Y(n_1405) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g491 ( .A(n_374), .Y(n_491) );
BUFx4f_ASAP7_75t_L g683 ( .A(n_374), .Y(n_683) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_376), .A2(n_399), .B1(n_446), .B2(n_448), .Y(n_445) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_SL g833 ( .A(n_380), .Y(n_833) );
INVx2_ASAP7_75t_L g872 ( .A(n_380), .Y(n_872) );
BUFx6f_ASAP7_75t_L g961 ( .A(n_380), .Y(n_961) );
INVx1_ASAP7_75t_L g1060 ( .A(n_380), .Y(n_1060) );
INVx2_ASAP7_75t_L g1277 ( .A(n_380), .Y(n_1277) );
INVx8_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g507 ( .A(n_381), .B(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g995 ( .A(n_381), .Y(n_995) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_395), .Y(n_389) );
AND2x4_ASAP7_75t_L g1407 ( .A(n_390), .B(n_395), .Y(n_1407) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g403 ( .A(n_392), .B(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_392), .Y(n_485) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_392), .B(n_395), .Y(n_631) );
OR2x2_ASAP7_75t_L g718 ( .A(n_392), .B(n_552), .Y(n_718) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g529 ( .A(n_393), .Y(n_529) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_395), .B(n_695), .C(n_697), .D(n_699), .Y(n_694) );
INVx4_ASAP7_75t_L g813 ( .A(n_395), .Y(n_813) );
INVx1_ASAP7_75t_SL g862 ( .A(n_395), .Y(n_862) );
INVx4_ASAP7_75t_L g989 ( .A(n_395), .Y(n_989) );
INVx1_ASAP7_75t_L g527 ( .A(n_396), .Y(n_527) );
AND2x4_ASAP7_75t_L g707 ( .A(n_396), .B(n_493), .Y(n_707) );
OAI33xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_407), .A3(n_422), .B1(n_432), .B2(n_437), .B3(n_445), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_SL g1168 ( .A1(n_402), .A2(n_1169), .B1(n_1176), .B2(n_1177), .Y(n_1168) );
OAI33xp33_ASAP7_75t_L g1784 ( .A1(n_402), .A2(n_1083), .A3(n_1785), .B1(n_1788), .B2(n_1792), .B3(n_1796), .Y(n_1784) );
BUFx4f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_L g734 ( .A(n_403), .Y(n_734) );
BUFx4f_ASAP7_75t_L g1029 ( .A(n_403), .Y(n_1029) );
BUFx8_ASAP7_75t_L g1222 ( .A(n_403), .Y(n_1222) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_404), .Y(n_1352) );
NAND2xp33_ASAP7_75t_SL g404 ( .A(n_405), .B(n_406), .Y(n_404) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_405), .Y(n_483) );
AND2x2_ASAP7_75t_L g565 ( .A(n_405), .B(n_469), .Y(n_565) );
INVx1_ASAP7_75t_L g582 ( .A(n_405), .Y(n_582) );
AND3x4_ASAP7_75t_L g773 ( .A(n_405), .B(n_469), .C(n_600), .Y(n_773) );
INVx3_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
BUFx3_ASAP7_75t_L g469 ( .A(n_406), .Y(n_469) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_409), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g1785 ( .A1(n_409), .A2(n_416), .B1(n_1786), .B2(n_1787), .Y(n_1785) );
OAI22xp33_ASAP7_75t_L g1796 ( .A1(n_409), .A2(n_436), .B1(n_1797), .B2(n_1798), .Y(n_1796) );
BUFx4f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x4_ASAP7_75t_L g453 ( .A(n_410), .B(n_454), .Y(n_453) );
OR2x4_ASAP7_75t_L g478 ( .A(n_410), .B(n_441), .Y(n_478) );
INVx2_ASAP7_75t_L g755 ( .A(n_410), .Y(n_755) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_411), .Y(n_421) );
INVx2_ASAP7_75t_L g427 ( .A(n_411), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_411), .B(n_420), .Y(n_431) );
AND2x4_ASAP7_75t_L g462 ( .A(n_411), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g577 ( .A(n_412), .Y(n_577) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g426 ( .A(n_413), .Y(n_426) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g572 ( .A(n_417), .Y(n_572) );
OR2x2_ASAP7_75t_L g725 ( .A(n_417), .B(n_718), .Y(n_725) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g436 ( .A(n_418), .Y(n_436) );
BUFx2_ASAP7_75t_L g560 ( .A(n_418), .Y(n_560) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
BUFx2_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g463 ( .A(n_420), .Y(n_463) );
BUFx2_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
INVx2_ASAP7_75t_L g595 ( .A(n_421), .Y(n_595) );
AND2x4_ASAP7_75t_L g660 ( .A(n_421), .B(n_599), .Y(n_660) );
INVx1_ASAP7_75t_L g885 ( .A(n_423), .Y(n_885) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_424), .Y(n_434) );
AND2x4_ASAP7_75t_L g480 ( .A(n_424), .B(n_454), .Y(n_480) );
INVx2_ASAP7_75t_L g778 ( .A(n_424), .Y(n_778) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_424), .Y(n_916) );
INVx2_ASAP7_75t_L g1178 ( .A(n_424), .Y(n_1178) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g553 ( .A(n_425), .Y(n_553) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_425), .Y(n_563) );
BUFx8_ASAP7_75t_L g791 ( .A(n_425), .Y(n_791) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AND2x4_ASAP7_75t_L g576 ( .A(n_427), .B(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_428), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g448 ( .A(n_429), .Y(n_448) );
INVx3_ASAP7_75t_L g557 ( .A(n_429), .Y(n_557) );
CKINVDCx8_ASAP7_75t_R g1180 ( .A(n_429), .Y(n_1180) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g723 ( .A(n_430), .Y(n_723) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g458 ( .A(n_431), .Y(n_458) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI33xp33_ASAP7_75t_L g881 ( .A1(n_438), .A2(n_773), .A3(n_882), .B1(n_884), .B2(n_887), .B3(n_888), .Y(n_881) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g785 ( .A(n_439), .Y(n_785) );
BUFx2_ASAP7_75t_L g920 ( .A(n_439), .Y(n_920) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_439), .Y(n_1126) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g742 ( .A(n_440), .Y(n_742) );
NAND3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .C(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g454 ( .A(n_441), .Y(n_454) );
OR2x6_ASAP7_75t_L g457 ( .A(n_441), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g461 ( .A(n_441), .B(n_462), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_441), .B(n_444), .Y(n_578) );
AND2x4_ASAP7_75t_L g581 ( .A(n_441), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_443), .B(n_540), .Y(n_628) );
INVx1_ASAP7_75t_L g655 ( .A(n_443), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g1007 ( .A1(n_446), .A2(n_994), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g735 ( .A1(n_448), .A2(n_567), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_448), .A2(n_778), .B1(n_985), .B2(n_1006), .Y(n_1005) );
OAI31xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_459), .A3(n_475), .B(n_481), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g1013 ( .A(n_458), .Y(n_1013) );
INVx1_ASAP7_75t_L g1173 ( .A(n_458), .Y(n_1173) );
CKINVDCx8_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g589 ( .A(n_462), .Y(n_589) );
BUFx3_ASAP7_75t_L g740 ( .A(n_462), .Y(n_740) );
BUFx2_ASAP7_75t_L g763 ( .A(n_462), .Y(n_763) );
BUFx2_ASAP7_75t_L g784 ( .A(n_462), .Y(n_784) );
BUFx2_ASAP7_75t_L g883 ( .A(n_462), .Y(n_883) );
BUFx2_ASAP7_75t_L g925 ( .A(n_462), .Y(n_925) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_462), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_462), .B(n_1357), .Y(n_1359) );
INVx1_ASAP7_75t_L g599 ( .A(n_463), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_471), .B2(n_472), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_465), .A2(n_516), .B1(n_519), .B2(n_520), .Y(n_515) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
AND2x4_ASAP7_75t_L g473 ( .A(n_468), .B(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI31xp33_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_500), .A3(n_509), .B(n_525), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_489), .B(n_1468), .Y(n_1467) );
AND2x4_ASAP7_75t_SL g1746 ( .A(n_489), .B(n_1747), .Y(n_1746) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
OR2x6_ASAP7_75t_L g502 ( .A(n_491), .B(n_496), .Y(n_502) );
INVxp67_ASAP7_75t_L g1275 ( .A(n_491), .Y(n_1275) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g512 ( .A(n_493), .Y(n_512) );
INVx3_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
INVx2_ASAP7_75t_L g607 ( .A(n_498), .Y(n_607) );
BUFx3_ASAP7_75t_L g696 ( .A(n_498), .Y(n_696) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g517 ( .A(n_508), .B(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
AND2x4_ASAP7_75t_SL g677 ( .A(n_513), .B(n_540), .Y(n_677) );
BUFx3_ASAP7_75t_L g700 ( .A(n_513), .Y(n_700) );
AND2x6_ASAP7_75t_L g814 ( .A(n_513), .B(n_617), .Y(n_814) );
BUFx3_ASAP7_75t_L g839 ( .A(n_513), .Y(n_839) );
INVx1_ASAP7_75t_L g861 ( .A(n_513), .Y(n_861) );
BUFx3_ASAP7_75t_L g998 ( .A(n_513), .Y(n_998) );
BUFx6f_ASAP7_75t_L g1095 ( .A(n_513), .Y(n_1095) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_513), .Y(n_1101) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g938 ( .A(n_514), .Y(n_938) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g624 ( .A(n_518), .Y(n_624) );
BUFx2_ASAP7_75t_L g688 ( .A(n_518), .Y(n_688) );
INVx1_ASAP7_75t_L g828 ( .A(n_518), .Y(n_828) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_523), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g1468 ( .A(n_527), .Y(n_1468) );
NOR2xp33_ASAP7_75t_L g1747 ( .A(n_527), .B(n_1460), .Y(n_1747) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g538 ( .A(n_529), .Y(n_538) );
OR2x2_ASAP7_75t_L g615 ( .A(n_529), .B(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_L g645 ( .A(n_529), .Y(n_645) );
OR2x2_ASAP7_75t_L g800 ( .A(n_529), .B(n_616), .Y(n_800) );
INVx1_ASAP7_75t_L g662 ( .A(n_530), .Y(n_662) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
XNOR2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_601), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_547), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B1(n_543), .B2(n_544), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_536), .A2(n_585), .B1(n_587), .B2(n_588), .Y(n_584) );
INVx3_ASAP7_75t_L g752 ( .A(n_537), .Y(n_752) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_537), .Y(n_1372) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x4_ASAP7_75t_L g544 ( .A(n_538), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g818 ( .A(n_539), .Y(n_818) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_539), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_539), .A2(n_821), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AND2x2_ASAP7_75t_L g545 ( .A(n_540), .B(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g692 ( .A(n_540), .Y(n_692) );
AND2x4_ASAP7_75t_L g804 ( .A(n_540), .B(n_611), .Y(n_804) );
AND2x4_ASAP7_75t_L g821 ( .A(n_540), .B(n_546), .Y(n_821) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_540), .B(n_649), .Y(n_1047) );
INVx3_ASAP7_75t_L g610 ( .A(n_541), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_541), .B(n_617), .Y(n_656) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_541), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_544), .B(n_1368), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_544), .B(n_1376), .Y(n_1375) );
INVx2_ASAP7_75t_L g1732 ( .A(n_544), .Y(n_1732) );
INVx2_ASAP7_75t_L g812 ( .A(n_546), .Y(n_812) );
BUFx6f_ASAP7_75t_L g940 ( .A(n_546), .Y(n_940) );
INVx1_ASAP7_75t_L g1208 ( .A(n_546), .Y(n_1208) );
OAI31xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_554), .A3(n_583), .B(n_600), .Y(n_547) );
OR2x6_ASAP7_75t_SL g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_551), .Y(n_591) );
AND2x4_ASAP7_75t_L g659 ( .A(n_551), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g1357 ( .A(n_552), .Y(n_1357) );
INVx3_ASAP7_75t_L g716 ( .A(n_553), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_553), .A2(n_1170), .B1(n_1171), .B2(n_1174), .C(n_1175), .Y(n_1169) );
INVx1_ASAP7_75t_L g1347 ( .A(n_553), .Y(n_1347) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_553), .Y(n_1430) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_559), .B1(n_566), .B2(n_570), .C(n_579), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_562), .B2(n_564), .C(n_565), .Y(n_559) );
OR2x6_ASAP7_75t_L g579 ( .A(n_560), .B(n_580), .Y(n_579) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_561), .A2(n_633), .B(n_635), .C(n_637), .Y(n_632) );
INVx2_ASAP7_75t_L g1351 ( .A(n_562), .Y(n_1351) );
OAI221xp5_ASAP7_75t_L g1384 ( .A1(n_562), .A2(n_745), .B1(n_1385), .B2(n_1386), .C(n_1387), .Y(n_1384) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_SL g567 ( .A(n_563), .Y(n_567) );
INVx5_ASAP7_75t_L g744 ( .A(n_563), .Y(n_744) );
OAI211xp5_ASAP7_75t_L g1030 ( .A1(n_567), .A2(n_1031), .B(n_1032), .C(n_1034), .Y(n_1030) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_573), .B(n_574), .Y(n_570) );
OAI211xp5_ASAP7_75t_L g1393 ( .A1(n_571), .A2(n_1394), .B(n_1395), .C(n_1396), .Y(n_1393) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g1009 ( .A(n_572), .Y(n_1009) );
BUFx2_ASAP7_75t_L g889 ( .A(n_575), .Y(n_889) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx8_ASAP7_75t_L g586 ( .A(n_576), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_576), .B(n_581), .Y(n_644) );
BUFx3_ASAP7_75t_L g739 ( .A(n_576), .Y(n_739) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_576), .Y(n_748) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_576), .B(n_1357), .Y(n_1356) );
INVx3_ASAP7_75t_L g1390 ( .A(n_578), .Y(n_1390) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x6_ASAP7_75t_L g593 ( .A(n_581), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g597 ( .A(n_581), .B(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g729 ( .A(n_581), .B(n_655), .Y(n_729) );
AND2x4_ASAP7_75t_L g929 ( .A(n_585), .B(n_790), .Y(n_929) );
AND2x4_ASAP7_75t_L g1105 ( .A(n_585), .B(n_790), .Y(n_1105) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx8_ASAP7_75t_L g775 ( .A(n_586), .Y(n_775) );
INVx3_ASAP7_75t_L g922 ( .A(n_586), .Y(n_922) );
INVx2_ASAP7_75t_L g1015 ( .A(n_586), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_586), .Y(n_1388) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_587), .A2(n_614), .B1(n_618), .B2(n_619), .Y(n_613) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g890 ( .A(n_589), .Y(n_890) );
INVx2_ASAP7_75t_L g914 ( .A(n_589), .Y(n_914) );
INVx1_ASAP7_75t_L g1016 ( .A(n_589), .Y(n_1016) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_593), .A2(n_597), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
NAND2x1_ASAP7_75t_L g728 ( .A(n_594), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g893 ( .A(n_594), .B(n_729), .Y(n_893) );
AND2x2_ASAP7_75t_L g904 ( .A(n_594), .B(n_729), .Y(n_904) );
AND2x4_ASAP7_75t_SL g1079 ( .A(n_594), .B(n_729), .Y(n_1079) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g732 ( .A(n_598), .Y(n_732) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g712 ( .A(n_600), .Y(n_712) );
INVx2_ASAP7_75t_SL g841 ( .A(n_600), .Y(n_841) );
OAI31xp33_ASAP7_75t_SL g1377 ( .A1(n_600), .A2(n_1378), .A3(n_1379), .B(n_1383), .Y(n_1377) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_640), .C(n_651), .Y(n_601) );
NOR3xp33_ASAP7_75t_SL g602 ( .A(n_603), .B(n_625), .C(n_629), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_608), .B(n_613), .Y(n_603) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g838 ( .A(n_607), .Y(n_838) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g698 ( .A(n_610), .Y(n_698) );
INVx2_ASAP7_75t_L g807 ( .A(n_610), .Y(n_807) );
INVx2_ASAP7_75t_L g1097 ( .A(n_610), .Y(n_1097) );
INVx2_ASAP7_75t_SL g1198 ( .A(n_610), .Y(n_1198) );
BUFx2_ASAP7_75t_L g808 ( .A(n_611), .Y(n_808) );
INVx1_ASAP7_75t_L g1136 ( .A(n_611), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx3_ASAP7_75t_L g636 ( .A(n_612), .Y(n_636) );
INVx2_ASAP7_75t_L g650 ( .A(n_612), .Y(n_650) );
BUFx3_ASAP7_75t_L g944 ( .A(n_612), .Y(n_944) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g1766 ( .A(n_616), .Y(n_1766) );
INVx1_ASAP7_75t_L g680 ( .A(n_617), .Y(n_680) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_617), .B(n_688), .Y(n_1102) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g1410 ( .A(n_620), .Y(n_1410) );
NAND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g639 ( .A(n_621), .Y(n_639) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx2_ASAP7_75t_SL g704 ( .A(n_627), .Y(n_704) );
BUFx2_ASAP7_75t_SL g1144 ( .A(n_627), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_627), .B(n_628), .Y(n_1339) );
INVx1_ASAP7_75t_L g648 ( .A(n_628), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_638), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_638), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
OR2x6_ASAP7_75t_L g760 ( .A(n_644), .B(n_645), .Y(n_760) );
INVx2_ASAP7_75t_L g1363 ( .A(n_644), .Y(n_1363) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g1332 ( .A1(n_647), .A2(n_1333), .B1(n_1336), .B2(n_1337), .C1(n_1338), .C2(n_1340), .Y(n_1332) );
AOI222xp33_ASAP7_75t_L g1408 ( .A1(n_647), .A2(n_1381), .B1(n_1392), .B2(n_1409), .C1(n_1410), .C2(n_1411), .Y(n_1408) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g864 ( .A(n_650), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
AND2x4_ASAP7_75t_L g796 ( .A(n_654), .B(n_722), .Y(n_796) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g1334 ( .A(n_655), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_656), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g876 ( .A(n_658), .Y(n_876) );
BUFx2_ASAP7_75t_L g963 ( .A(n_658), .Y(n_963) );
AOI21xp5_ASAP7_75t_SL g1754 ( .A1(n_658), .A2(n_1755), .B(n_1768), .Y(n_1754) );
INVx3_ASAP7_75t_L g1366 ( .A(n_659), .Y(n_1366) );
INVx5_ASAP7_75t_L g780 ( .A(n_660), .Y(n_780) );
BUFx12f_ASAP7_75t_L g782 ( .A(n_660), .Y(n_782) );
BUFx3_ASAP7_75t_L g886 ( .A(n_660), .Y(n_886) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_660), .Y(n_1348) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_1453), .C(n_1456), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_1107), .C(n_1415), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g1456 ( .A(n_665), .B(n_1454), .C(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g1453 ( .A1(n_666), .A2(n_1107), .B1(n_1108), .B2(n_1415), .C(n_1454), .Y(n_1453) );
XNOR2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_966), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_843), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_764), .B1(n_765), .B2(n_842), .Y(n_669) );
INVx2_ASAP7_75t_L g842 ( .A(n_670), .Y(n_842) );
AND5x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_726), .C(n_749), .D(n_757), .E(n_761), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_710), .B(n_713), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_674), .B(n_678), .C(n_694), .D(n_701), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AOI221x1_ASAP7_75t_L g726 ( .A1(n_675), .A2(n_687), .B1(n_727), .B2(n_730), .C(n_733), .Y(n_726) );
AOI222xp33_ASAP7_75t_L g1098 ( .A1(n_676), .A2(n_1078), .B1(n_1080), .B2(n_1099), .C1(n_1100), .C2(n_1102), .Y(n_1098) );
AOI222xp33_ASAP7_75t_L g1290 ( .A1(n_676), .A2(n_1102), .B1(n_1291), .B2(n_1292), .C1(n_1293), .C2(n_1295), .Y(n_1290) );
BUFx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g825 ( .A(n_677), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B1(n_692), .B2(n_693), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g1720 ( .A1(n_679), .A2(n_692), .B1(n_1721), .B2(n_1726), .Y(n_1720) );
A2O1A1Ixp33_ASAP7_75t_L g1761 ( .A1(n_679), .A2(n_700), .B(n_1762), .C(n_1763), .Y(n_1761) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2x1_ASAP7_75t_L g827 ( .A(n_680), .B(n_828), .Y(n_827) );
INVx4_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx6f_ASAP7_75t_L g958 ( .A(n_683), .Y(n_958) );
INVx3_ASAP7_75t_L g1722 ( .A(n_683), .Y(n_1722) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_684), .A2(n_1147), .B1(n_1269), .B2(n_1270), .C(n_1271), .Y(n_1268) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g1195 ( .A(n_685), .Y(n_1195) );
INVx2_ASAP7_75t_L g1723 ( .A(n_685), .Y(n_1723) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g1724 ( .A1(n_688), .A2(n_690), .B1(n_1709), .B2(n_1725), .Y(n_1724) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_689), .A2(n_720), .B1(n_721), .B2(n_724), .Y(n_719) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g1755 ( .A1(n_692), .A2(n_1756), .B(n_1760), .Y(n_1755) );
AOI22xp33_ASAP7_75t_L g1757 ( .A1(n_700), .A2(n_944), .B1(n_1758), .B2(n_1759), .Y(n_1757) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_705), .C(n_708), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_702), .A2(n_744), .B1(n_745), .B2(n_746), .C(n_747), .Y(n_743) );
OAI211xp5_ASAP7_75t_L g1214 ( .A1(n_703), .A2(n_1215), .B(n_1216), .C(n_1218), .Y(n_1214) );
OAI211xp5_ASAP7_75t_L g1449 ( .A1(n_703), .A2(n_1450), .B(n_1451), .C(n_1452), .Y(n_1449) );
INVx5_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g840 ( .A(n_707), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_707), .A2(n_949), .B1(n_950), .B2(n_951), .C(n_954), .Y(n_948) );
INVx2_ASAP7_75t_L g1067 ( .A(n_707), .Y(n_1067) );
INVx1_ASAP7_75t_L g1217 ( .A(n_707), .Y(n_1217) );
INVx3_ASAP7_75t_L g1051 ( .A(n_709), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g1134 ( .A(n_709), .Y(n_1134) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g1344 ( .A1(n_711), .A2(n_1345), .B(n_1360), .C(n_1367), .Y(n_1344) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_712), .Y(n_1219) );
AOI21x1_ASAP7_75t_L g1712 ( .A1(n_712), .A2(n_1713), .B(n_1728), .Y(n_1712) );
NAND2x1_ASAP7_75t_L g1731 ( .A(n_714), .B(n_1732), .Y(n_1731) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_715), .A2(n_1091), .B1(n_1092), .B2(n_1105), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_715), .A2(n_1105), .B1(n_1264), .B2(n_1265), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_715), .A2(n_929), .B1(n_1301), .B2(n_1302), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1778 ( .A1(n_715), .A2(n_724), .B1(n_1767), .B2(n_1779), .Y(n_1778) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx2_ASAP7_75t_L g1036 ( .A(n_716), .Y(n_1036) );
INVx2_ASAP7_75t_L g1793 ( .A(n_716), .Y(n_1793) );
INVxp67_ASAP7_75t_L g756 ( .A(n_717), .Y(n_756) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g722 ( .A(n_718), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g790 ( .A(n_718), .Y(n_790) );
AOI222xp33_ASAP7_75t_L g1735 ( .A1(n_721), .A2(n_724), .B1(n_1105), .B2(n_1725), .C1(n_1736), .C2(n_1737), .Y(n_1735) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
BUFx3_ASAP7_75t_L g745 ( .A(n_723), .Y(n_745) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g799 ( .A(n_725), .B(n_800), .Y(n_799) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_725), .B(n_800), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_727), .A2(n_730), .B1(n_770), .B2(n_771), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_727), .A2(n_1114), .B1(n_1115), .B2(n_1116), .Y(n_1113) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g730 ( .A(n_729), .B(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g762 ( .A(n_729), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_SL g1043 ( .A(n_729), .B(n_731), .Y(n_1043) );
A2O1A1Ixp33_ASAP7_75t_L g1782 ( .A1(n_729), .A2(n_775), .B(n_1758), .C(n_1783), .Y(n_1782) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_730), .A2(n_892), .B1(n_893), .B2(n_894), .Y(n_891) );
AO22x1_ASAP7_75t_L g902 ( .A1(n_730), .A2(n_903), .B1(n_904), .B2(n_905), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_730), .A2(n_904), .B1(n_973), .B2(n_974), .Y(n_972) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_730), .Y(n_1116) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_730), .A2(n_893), .B1(n_1422), .B2(n_1423), .Y(n_1421) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_735), .B1(n_741), .B2(n_743), .Y(n_733) );
INVx2_ASAP7_75t_SL g913 ( .A(n_739), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_741), .A2(n_1029), .B1(n_1030), .B2(n_1035), .Y(n_1028) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g1176 ( .A(n_742), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1228 ( .A(n_742), .Y(n_1228) );
AOI33xp33_ASAP7_75t_L g1426 ( .A1(n_742), .A2(n_910), .A3(n_1427), .B1(n_1428), .B2(n_1432), .B3(n_1435), .Y(n_1426) );
BUFx3_ASAP7_75t_L g1011 ( .A(n_744), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1788 ( .A1(n_744), .A2(n_1789), .B1(n_1790), .B2(n_1791), .Y(n_1788) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g1343 ( .A(n_752), .Y(n_1343) );
OR2x6_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
OR2x2_ASAP7_75t_L g787 ( .A(n_754), .B(n_756), .Y(n_787) );
INVx2_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_759), .B(n_908), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_759), .B(n_1118), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_759), .B(n_1247), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_759), .B(n_1425), .Y(n_1424) );
INVx5_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx3_ASAP7_75t_L g977 ( .A(n_760), .Y(n_977) );
AND4x1_ASAP7_75t_L g877 ( .A(n_761), .B(n_878), .C(n_881), .D(n_891), .Y(n_877) );
NAND5xp2_ASAP7_75t_L g971 ( .A(n_761), .B(n_972), .C(n_975), .D(n_978), .E(n_979), .Y(n_971) );
NAND3xp33_ASAP7_75t_SL g1076 ( .A(n_761), .B(n_1077), .C(n_1081), .Y(n_1076) );
AND4x1_ASAP7_75t_L g1112 ( .A(n_761), .B(n_1113), .C(n_1117), .D(n_1119), .Y(n_1112) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx3_ASAP7_75t_L g793 ( .A(n_762), .Y(n_793) );
NOR3xp33_ASAP7_75t_SL g1027 ( .A(n_762), .B(n_1028), .C(n_1040), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1167 ( .A(n_762), .Y(n_1167) );
NOR3xp33_ASAP7_75t_L g1220 ( .A(n_762), .B(n_1221), .C(n_1232), .Y(n_1220) );
AOI211xp5_ASAP7_75t_L g1305 ( .A1(n_762), .A2(n_977), .B(n_1297), .C(n_1306), .Y(n_1305) );
AOI221xp5_ASAP7_75t_L g1708 ( .A1(n_762), .A2(n_1043), .B1(n_1079), .B2(n_1709), .C(n_1710), .Y(n_1708) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_794), .C(n_801), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_786), .C(n_792), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .Y(n_768) );
AOI33xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .A3(n_776), .B1(n_781), .B2(n_783), .B3(n_785), .Y(n_772) );
BUFx3_ASAP7_75t_L g910 ( .A(n_773), .Y(n_910) );
INVx1_ASAP7_75t_L g1086 ( .A(n_773), .Y(n_1086) );
AOI33xp33_ASAP7_75t_L g1248 ( .A1(n_773), .A2(n_1249), .A3(n_1250), .B1(n_1252), .B2(n_1253), .B3(n_1254), .Y(n_1248) );
AOI33xp33_ASAP7_75t_L g1308 ( .A1(n_773), .A2(n_1309), .A3(n_1310), .B1(n_1311), .B2(n_1312), .B3(n_1313), .Y(n_1308) );
AOI33xp33_ASAP7_75t_L g1702 ( .A1(n_773), .A2(n_1703), .A3(n_1704), .B1(n_1705), .B2(n_1706), .B3(n_1707), .Y(n_1702) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_775), .Y(n_1125) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g917 ( .A(n_780), .Y(n_917) );
INVx1_ASAP7_75t_L g1431 ( .A(n_780), .Y(n_1431) );
BUFx2_ASAP7_75t_L g919 ( .A(n_782), .Y(n_919) );
INVxp67_ASAP7_75t_L g1070 ( .A(n_788), .Y(n_1070) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g880 ( .A(n_789), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_789), .A2(n_928), .B1(n_929), .B2(n_930), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_789), .A2(n_929), .B1(n_1138), .B2(n_1140), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_789), .A2(n_929), .B1(n_1191), .B2(n_1192), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_789), .A2(n_929), .B1(n_1211), .B2(n_1212), .Y(n_1236) );
AND2x4_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx2_ASAP7_75t_SL g1224 ( .A(n_791), .Y(n_1224) );
INVx3_ASAP7_75t_L g1434 ( .A(n_791), .Y(n_1434) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g906 ( .A(n_793), .B(n_907), .Y(n_906) );
AND4x1_ASAP7_75t_L g1242 ( .A(n_793), .B(n_1243), .C(n_1246), .D(n_1248), .Y(n_1242) );
NAND4xp25_ASAP7_75t_SL g1420 ( .A(n_793), .B(n_1421), .C(n_1424), .D(n_1426), .Y(n_1420) );
AOI21xp33_ASAP7_75t_SL g794 ( .A1(n_795), .A2(n_797), .B(n_798), .Y(n_794) );
AOI21xp33_ASAP7_75t_L g849 ( .A1(n_795), .A2(n_850), .B(n_851), .Y(n_849) );
AOI211x1_ASAP7_75t_L g898 ( .A1(n_795), .A2(n_899), .B(n_900), .C(n_926), .Y(n_898) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_795), .A2(n_977), .B1(n_1074), .B2(n_1075), .C(n_1076), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_795), .B(n_1155), .Y(n_1154) );
AOI21xp5_ASAP7_75t_L g1163 ( .A1(n_795), .A2(n_1164), .B(n_1165), .Y(n_1163) );
AOI21xp5_ASAP7_75t_L g1233 ( .A1(n_795), .A2(n_1234), .B(n_1235), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_795), .B(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_795), .B(n_1287), .Y(n_1286) );
AOI211x1_ASAP7_75t_L g1418 ( .A1(n_795), .A2(n_1419), .B(n_1420), .C(n_1436), .Y(n_1418) );
INVx8_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g1002 ( .A(n_799), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_799), .Y(n_1152) );
INVx2_ASAP7_75t_SL g1411 ( .A(n_800), .Y(n_1411) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_822), .B(n_841), .Y(n_801) );
INVx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_R g945 ( .A(n_804), .B(n_908), .Y(n_945) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_804), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_804), .B(n_1247), .Y(n_1266) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_809), .B(n_814), .Y(n_805) );
BUFx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g1066 ( .A(n_812), .Y(n_1066) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_814), .A2(n_859), .B(n_863), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g934 ( .A1(n_814), .A2(n_935), .B(n_941), .Y(n_934) );
INVx1_ASAP7_75t_L g990 ( .A(n_814), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_814), .A2(n_1026), .B1(n_1047), .B2(n_1048), .C(n_1049), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_814), .A2(n_1047), .B1(n_1074), .B2(n_1094), .C(n_1096), .Y(n_1093) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_814), .A2(n_1131), .B(n_1132), .Y(n_1130) );
AOI21xp5_ASAP7_75t_L g1186 ( .A1(n_814), .A2(n_1187), .B(n_1188), .Y(n_1186) );
AOI21xp5_ASAP7_75t_L g1205 ( .A1(n_814), .A2(n_1206), .B(n_1209), .Y(n_1205) );
AOI221xp5_ASAP7_75t_L g1296 ( .A1(n_814), .A2(n_1047), .B1(n_1297), .B2(n_1298), .C(n_1299), .Y(n_1296) );
AOI21xp5_ASAP7_75t_L g1442 ( .A1(n_814), .A2(n_1443), .B(n_1444), .Y(n_1442) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_817), .A2(n_821), .B1(n_928), .B2(n_930), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_817), .A2(n_1138), .B1(n_1139), .B2(n_1140), .Y(n_1137) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_820), .A2(n_855), .B1(n_856), .B2(n_857), .Y(n_854) );
INVxp67_ASAP7_75t_SL g992 ( .A(n_820), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_820), .A2(n_856), .B1(n_1446), .B2(n_1447), .Y(n_1445) );
BUFx6f_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_821), .A2(n_856), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_821), .A2(n_856), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_821), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_821), .A2(n_856), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
AOI22xp5_ASAP7_75t_L g1263 ( .A1(n_821), .A2(n_856), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_821), .A2(n_856), .B1(n_1301), .B2(n_1302), .Y(n_1300) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g947 ( .A(n_824), .Y(n_947) );
INVx2_ASAP7_75t_L g1142 ( .A(n_824), .Y(n_1142) );
INVx4_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g867 ( .A(n_827), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_832), .B2(n_834), .C(n_835), .Y(n_829) );
OAI221xp5_ASAP7_75t_L g984 ( .A1(n_830), .A2(n_985), .B1(n_986), .B2(n_987), .C(n_988), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_830), .A2(n_994), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_830), .A2(n_870), .B1(n_1149), .B2(n_1150), .Y(n_1148) );
INVx1_ASAP7_75t_L g1322 ( .A(n_830), .Y(n_1322) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_833), .Y(n_986) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g1771 ( .A(n_838), .Y(n_1771) );
INVx1_ASAP7_75t_L g1147 ( .A(n_840), .Y(n_1147) );
O2A1O1Ixp5_ASAP7_75t_L g1127 ( .A1(n_841), .A2(n_1128), .B(n_1141), .C(n_1151), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_896), .B2(n_965), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AO21x2_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B(n_895), .Y(n_846) );
NAND3xp33_ASAP7_75t_SL g848 ( .A(n_849), .B(n_852), .C(n_877), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_865), .B(n_876), .Y(n_852) );
INVx1_ASAP7_75t_L g1000 ( .A(n_856), .Y(n_1000) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g875 ( .A(n_861), .Y(n_875) );
BUFx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g1321 ( .A(n_871), .Y(n_1321) );
BUFx6f_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OAI31xp33_ASAP7_75t_L g982 ( .A1(n_876), .A2(n_983), .A3(n_991), .B(n_999), .Y(n_982) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1041 ( .A(n_893), .Y(n_1041) );
INVx2_ASAP7_75t_L g965 ( .A(n_896), .Y(n_965) );
XOR2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_964), .Y(n_896) );
NAND2xp5_ASAP7_75t_SL g897 ( .A(n_898), .B(n_931), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_901), .B(n_909), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_906), .Y(n_901) );
AOI33xp33_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_911), .A3(n_915), .B1(n_918), .B2(n_920), .B3(n_921), .Y(n_909) );
AOI33xp33_ASAP7_75t_L g1119 ( .A1(n_910), .A2(n_1120), .A3(n_1121), .B1(n_1123), .B2(n_1124), .B3(n_1126), .Y(n_1119) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_929), .B(n_980), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_929), .A2(n_1053), .B1(n_1054), .B2(n_1070), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1776 ( .A(n_929), .B(n_1777), .Y(n_1776) );
OAI21xp5_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_946), .B(n_962), .Y(n_931) );
NAND3xp33_ASAP7_75t_SL g932 ( .A(n_933), .B(n_934), .C(n_945), .Y(n_932) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1294 ( .A(n_937), .Y(n_1294) );
BUFx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g1065 ( .A(n_938), .Y(n_1065) );
BUFx3_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_SL g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_SL g943 ( .A(n_944), .Y(n_943) );
INVxp67_ASAP7_75t_SL g1325 ( .A(n_949), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_951), .A2(n_1144), .B1(n_1145), .B2(n_1146), .C(n_1147), .Y(n_1143) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx4_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_957), .B1(n_959), .B2(n_960), .Y(n_955) );
INVx2_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx5_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g1088 ( .A1(n_962), .A2(n_1089), .B(n_1103), .Y(n_1088) );
OAI21xp5_ASAP7_75t_L g1184 ( .A1(n_962), .A2(n_1185), .B(n_1193), .Y(n_1184) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g1068 ( .A(n_963), .Y(n_1068) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B1(n_1018), .B2(n_1106), .Y(n_967) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
XNOR2x1_ASAP7_75t_L g969 ( .A(n_970), .B(n_1017), .Y(n_969) );
NOR2x1_ASAP7_75t_L g970 ( .A(n_971), .B(n_981), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_977), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_977), .A2(n_1023), .B1(n_1024), .B2(n_1026), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_1001), .Y(n_981) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_987), .A2(n_1011), .B1(n_1012), .B2(n_1013), .C(n_1014), .Y(n_1010) );
NAND4xp25_ASAP7_75t_L g1257 ( .A(n_990), .B(n_1258), .C(n_1263), .D(n_1266), .Y(n_1257) );
INVx1_ASAP7_75t_L g1328 ( .A(n_995), .Y(n_1328) );
AOI21xp5_ASAP7_75t_SL g1001 ( .A1(n_1002), .A2(n_1003), .B(n_1004), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g1437 ( .A1(n_1002), .A2(n_1438), .B(n_1439), .Y(n_1437) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1011), .Y(n_1122) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_1013), .A2(n_1036), .B1(n_1037), .B2(n_1038), .C(n_1039), .Y(n_1035) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1018), .Y(n_1106) );
XNOR2x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1071), .Y(n_1018) );
NAND4xp75_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1027), .C(n_1044), .D(n_1069), .Y(n_1020) );
INVx1_ASAP7_75t_SL g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_1043), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1243 ( .A1(n_1043), .A2(n_1079), .B1(n_1244), .B2(n_1245), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_1043), .A2(n_1079), .B1(n_1291), .B2(n_1292), .Y(n_1307) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1055), .B(n_1068), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1052), .Y(n_1045) );
INVx2_ASAP7_75t_L g1714 ( .A(n_1047), .Y(n_1714) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_1051), .Y(n_1189) );
INVx2_ASAP7_75t_L g1762 ( .A(n_1051), .Y(n_1762) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1059), .B2(n_1061), .C(n_1062), .Y(n_1056) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
AOI21xp5_ASAP7_75t_L g1288 ( .A1(n_1068), .A2(n_1289), .B(n_1303), .Y(n_1288) );
OAI21xp33_ASAP7_75t_L g1440 ( .A1(n_1068), .A2(n_1441), .B(n_1448), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1088), .Y(n_1072) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1084), .B1(n_1085), .B2(n_1087), .Y(n_1081) );
NAND3xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1093), .C(n_1098), .Y(n_1089) );
AOI22xp33_ASAP7_75t_SL g1764 ( .A1(n_1102), .A2(n_1765), .B1(n_1766), .B2(n_1767), .Y(n_1764) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1107), .Y(n_1457) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
OA22x2_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1110), .B1(n_1157), .B2(n_1158), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
XOR2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1156), .Y(n_1110) );
NAND3x1_ASAP7_75t_SL g1111 ( .A(n_1112), .B(n_1127), .C(n_1154), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
XNOR2x1_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1238), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
AO22x2_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1200), .B1(n_1201), .B2(n_1237), .Y(n_1160) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1161), .Y(n_1237) );
AND4x1_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1166), .C(n_1184), .D(n_1199), .Y(n_1162) );
NOR3xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1168), .C(n_1183), .Y(n_1166) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_1171), .A2(n_1224), .B1(n_1225), .B2(n_1226), .C(n_1227), .Y(n_1223) );
INVx3_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
BUFx2_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1173), .Y(n_1790) );
OAI221xp5_ASAP7_75t_L g1177 ( .A1(n_1178), .A2(n_1179), .B1(n_1180), .B2(n_1181), .C(n_1182), .Y(n_1177) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1178), .Y(n_1251) );
OAI211xp5_ASAP7_75t_L g1194 ( .A1(n_1179), .A2(n_1195), .B(n_1196), .C(n_1197), .Y(n_1194) );
OAI221xp5_ASAP7_75t_L g1229 ( .A1(n_1180), .A2(n_1215), .B1(n_1224), .B2(n_1230), .C(n_1231), .Y(n_1229) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AND4x1_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1220), .C(n_1233), .D(n_1236), .Y(n_1202) );
OAI21xp5_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1213), .B(n_1219), .Y(n_1203) );
INVx2_ASAP7_75t_SL g1207 ( .A(n_1208), .Y(n_1207) );
O2A1O1Ixp5_ASAP7_75t_SL g1256 ( .A1(n_1219), .A2(n_1257), .B(n_1267), .C(n_1278), .Y(n_1256) );
OAI22xp5_ASAP7_75t_SL g1221 ( .A1(n_1222), .A2(n_1223), .B1(n_1228), .B2(n_1229), .Y(n_1221) );
XOR2xp5_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1315), .Y(n_1238) );
XNOR2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1283), .Y(n_1239) );
XOR2xp5_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1282), .Y(n_1240) );
NAND3xp33_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1256), .C(n_1280), .Y(n_1241) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_SL g1313 ( .A(n_1255), .Y(n_1313) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1255), .Y(n_1707) );
OAI211xp5_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1260), .B(n_1261), .C(n_1262), .Y(n_1258) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1270), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1274), .B1(n_1276), .B2(n_1277), .Y(n_1272) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
NAND3xp33_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1288), .C(n_1305), .Y(n_1285) );
NAND3xp33_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1296), .C(n_1300), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
XNOR2x1_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1370), .Y(n_1315) );
XNOR2x1_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1369), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1344), .Y(n_1317) );
NAND3xp33_ASAP7_75t_SL g1318 ( .A(n_1319), .B(n_1332), .C(n_1341), .Y(n_1318) );
AOI211xp5_ASAP7_75t_SL g1319 ( .A1(n_1320), .A2(n_1323), .B(n_1326), .C(n_1327), .Y(n_1319) );
AOI21xp33_ASAP7_75t_SL g1412 ( .A1(n_1333), .A2(n_1413), .B(n_1414), .Y(n_1412) );
AND2x4_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1335), .Y(n_1333) );
AOI211xp5_ASAP7_75t_L g1360 ( .A1(n_1337), .A2(n_1361), .B(n_1364), .C(n_1365), .Y(n_1360) );
AOI222xp33_ASAP7_75t_L g1398 ( .A1(n_1338), .A2(n_1382), .B1(n_1399), .B2(n_1403), .C1(n_1404), .C2(n_1407), .Y(n_1398) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
AOI221xp5_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1349), .B1(n_1350), .B2(n_1353), .C(n_1354), .Y(n_1345) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1391 ( .A1(n_1356), .A2(n_1359), .B1(n_1373), .B2(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
AOI211x1_ASAP7_75t_L g1371 ( .A1(n_1372), .A2(n_1373), .B(n_1374), .C(n_1397), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1377), .Y(n_1374) );
NAND3xp33_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1391), .C(n_1393), .Y(n_1383) );
INVx3_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NAND3xp33_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1408), .C(n_1412), .Y(n_1397) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1416), .Y(n_1455) );
XNOR2x2_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1440), .Y(n_1436) );
INVx1_ASAP7_75t_SL g1454 ( .A(n_1455), .Y(n_1454) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1466), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1464), .Y(n_1461) );
NOR2xp33_ASAP7_75t_L g1743 ( .A(n_1462), .B(n_1465), .Y(n_1743) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1462), .Y(n_1802) );
HB1xp67_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
NOR2xp33_ASAP7_75t_L g1804 ( .A(n_1465), .B(n_1802), .Y(n_1804) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1695), .B1(n_1698), .B2(n_1740), .C(n_1744), .Y(n_1469) );
NOR5xp2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1610), .C(n_1672), .D(n_1678), .E(n_1689), .Y(n_1470) );
AOI31xp33_ASAP7_75t_L g1471 ( .A1(n_1472), .A2(n_1554), .A3(n_1584), .B(n_1604), .Y(n_1471) );
AOI211xp5_ASAP7_75t_SL g1472 ( .A1(n_1473), .A2(n_1489), .B(n_1508), .C(n_1522), .Y(n_1472) );
A2O1A1Ixp33_ASAP7_75t_L g1611 ( .A1(n_1473), .A2(n_1612), .B(n_1614), .C(n_1626), .Y(n_1611) );
CKINVDCx6p67_ASAP7_75t_R g1473 ( .A(n_1474), .Y(n_1473) );
CKINVDCx6p67_ASAP7_75t_R g1474 ( .A(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1475), .B(n_1550), .Y(n_1552) );
INVx2_ASAP7_75t_L g1562 ( .A(n_1475), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1621 ( .A(n_1475), .B(n_1622), .Y(n_1621) );
OAI22xp5_ASAP7_75t_L g1632 ( .A1(n_1475), .A2(n_1633), .B1(n_1635), .B2(n_1637), .Y(n_1632) );
AND2x4_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1483), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1476), .B(n_1483), .Y(n_1514) );
AND2x6_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1479), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1478), .B(n_1482), .Y(n_1481) );
AND2x4_ASAP7_75t_L g1484 ( .A(n_1478), .B(n_1485), .Y(n_1484) );
AND2x6_ASAP7_75t_L g1487 ( .A(n_1478), .B(n_1488), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1478), .B(n_1482), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1478), .B(n_1482), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1480), .B(n_1486), .Y(n_1485) );
INVx2_ASAP7_75t_L g1697 ( .A(n_1487), .Y(n_1697) );
HB1xp67_ASAP7_75t_L g1801 ( .A(n_1488), .Y(n_1801) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1496), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1491), .B(n_1537), .Y(n_1536) );
NAND2xp5_ASAP7_75t_SL g1558 ( .A(n_1491), .B(n_1559), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1491), .B(n_1638), .Y(n_1637) );
INVx2_ASAP7_75t_L g1641 ( .A(n_1491), .Y(n_1641) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx3_ASAP7_75t_L g1516 ( .A(n_1492), .Y(n_1516) );
NOR2xp33_ASAP7_75t_L g1534 ( .A(n_1492), .B(n_1497), .Y(n_1534) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1492), .B(n_1567), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1492), .B(n_1497), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1492), .B(n_1531), .Y(n_1593) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1492), .B(n_1580), .Y(n_1623) );
NOR2xp33_ASAP7_75t_L g1631 ( .A(n_1492), .B(n_1542), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1494), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1496), .B(n_1526), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1501), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g1557 ( .A(n_1497), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1497), .B(n_1569), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1497), .B(n_1520), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1658 ( .A(n_1497), .B(n_1533), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_1497), .B(n_1594), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1500), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1498), .B(n_1500), .Y(n_1518) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1501), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1501), .B(n_1589), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1501), .B(n_1557), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1505), .Y(n_1501) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1502), .Y(n_1521) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1502), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1504), .Y(n_1502) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1505), .Y(n_1520) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1505), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1505), .B(n_1521), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1560 ( .A(n_1505), .B(n_1521), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1507), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1515), .Y(n_1508) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
OR2x2_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1514), .Y(n_1510) );
INVx3_ASAP7_75t_L g1531 ( .A(n_1511), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1511), .B(n_1548), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1511), .B(n_1562), .Y(n_1561) );
OR2x2_ASAP7_75t_L g1564 ( .A(n_1511), .B(n_1549), .Y(n_1564) );
NOR2xp33_ASAP7_75t_L g1572 ( .A(n_1511), .B(n_1525), .Y(n_1572) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1511), .B(n_1514), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1511), .B(n_1525), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1511), .B(n_1576), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1636 ( .A(n_1511), .B(n_1580), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1511), .B(n_1626), .Y(n_1644) );
INVx3_ASAP7_75t_L g1688 ( .A(n_1511), .Y(n_1688) );
AND2x4_ASAP7_75t_SL g1511 ( .A(n_1512), .B(n_1513), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1514), .B(n_1531), .Y(n_1530) );
OR2x2_ASAP7_75t_L g1538 ( .A(n_1514), .B(n_1527), .Y(n_1538) );
OR2x2_ASAP7_75t_L g1549 ( .A(n_1514), .B(n_1550), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1514), .B(n_1527), .Y(n_1576) );
NOR2xp33_ASAP7_75t_L g1659 ( .A(n_1514), .B(n_1607), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1517), .Y(n_1515) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1516), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1516), .B(n_1546), .Y(n_1613) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1516), .B(n_1560), .Y(n_1616) );
O2A1O1Ixp33_ASAP7_75t_L g1618 ( .A1(n_1516), .A2(n_1576), .B(n_1619), .C(n_1620), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1516), .B(n_1550), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1516), .B(n_1652), .Y(n_1651) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1516), .B(n_1658), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1660 ( .A(n_1516), .B(n_1661), .Y(n_1660) );
NAND3xp33_ASAP7_75t_L g1664 ( .A(n_1516), .B(n_1626), .C(n_1665), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1516), .B(n_1548), .Y(n_1681) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1517), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1519), .Y(n_1517) );
AOI32xp33_ASAP7_75t_L g1535 ( .A1(n_1518), .A2(n_1536), .A3(n_1539), .B1(n_1543), .B2(n_1547), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1544 ( .A(n_1518), .B(n_1545), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1518), .B(n_1583), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1518), .B(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1519), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1519), .B(n_1557), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1519), .B(n_1534), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1519), .B(n_1603), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1521), .Y(n_1519) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1521), .Y(n_1569) );
OAI211xp5_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1532), .B(n_1535), .C(n_1551), .Y(n_1522) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1530), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1525), .B(n_1588), .Y(n_1634) );
O2A1O1Ixp33_ASAP7_75t_L g1682 ( .A1(n_1525), .A2(n_1613), .B(n_1619), .C(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1525), .Y(n_1685) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1526), .B(n_1588), .Y(n_1587) );
AOI322xp5_ASAP7_75t_L g1656 ( .A1(n_1526), .A2(n_1572), .A3(n_1598), .B1(n_1644), .B2(n_1657), .C1(n_1659), .C2(n_1660), .Y(n_1656) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1527), .Y(n_1550) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1527), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1529), .Y(n_1527) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1530), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1655 ( .A(n_1531), .B(n_1537), .Y(n_1655) );
OR2x2_ASAP7_75t_L g1667 ( .A(n_1531), .B(n_1538), .Y(n_1667) );
AOI32xp33_ASAP7_75t_L g1691 ( .A1(n_1531), .A2(n_1536), .A3(n_1625), .B1(n_1626), .B2(n_1692), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1534), .Y(n_1532) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1533), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1534), .B(n_1546), .Y(n_1553) );
AOI311xp33_ASAP7_75t_L g1639 ( .A1(n_1537), .A2(n_1640), .A3(n_1641), .B(n_1642), .C(n_1653), .Y(n_1639) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
OAI321xp33_ASAP7_75t_L g1590 ( .A1(n_1538), .A2(n_1591), .A3(n_1592), .B1(n_1594), .B2(n_1595), .C(n_1597), .Y(n_1590) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1542), .Y(n_1540) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
OR2x2_ASAP7_75t_L g1694 ( .A(n_1545), .B(n_1557), .Y(n_1694) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1546), .B(n_1575), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1546), .B(n_1589), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1548), .B(n_1575), .Y(n_1671) );
INVx2_ASAP7_75t_SL g1548 ( .A(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1553), .Y(n_1551) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1552), .Y(n_1591) );
AOI221xp5_ASAP7_75t_L g1554 ( .A1(n_1555), .A2(n_1561), .B1(n_1563), .B2(n_1565), .C(n_1570), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
OR2x2_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1557), .B(n_1594), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1557), .B(n_1616), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1557), .B(n_1569), .Y(n_1652) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1559), .B(n_1589), .Y(n_1654) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1561), .Y(n_1617) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVxp67_ASAP7_75t_SL g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
A2O1A1Ixp33_ASAP7_75t_L g1570 ( .A1(n_1571), .A2(n_1573), .B(n_1577), .C(n_1578), .Y(n_1570) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1576), .Y(n_1574) );
CKINVDCx14_ASAP7_75t_R g1690 ( .A(n_1576), .Y(n_1690) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1577), .B(n_1638), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1581), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1673 ( .A(n_1579), .B(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1582), .B(n_1630), .Y(n_1629) );
AOI211xp5_ASAP7_75t_L g1584 ( .A1(n_1585), .A2(n_1587), .B(n_1590), .C(n_1601), .Y(n_1584) );
NAND3xp33_ASAP7_75t_L g1649 ( .A(n_1585), .B(n_1606), .C(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
A2O1A1Ixp33_ASAP7_75t_L g1642 ( .A1(n_1586), .A2(n_1643), .B(n_1645), .C(n_1649), .Y(n_1642) );
NOR2xp33_ASAP7_75t_L g1620 ( .A(n_1591), .B(n_1595), .Y(n_1620) );
OAI221xp5_ASAP7_75t_SL g1653 ( .A1(n_1591), .A2(n_1595), .B1(n_1654), .B2(n_1655), .C(n_1656), .Y(n_1653) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1594), .Y(n_1665) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
OAI21xp5_ASAP7_75t_L g1597 ( .A1(n_1598), .A2(n_1599), .B(n_1600), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1599), .B(n_1685), .Y(n_1684) );
AOI221xp5_ASAP7_75t_L g1627 ( .A1(n_1600), .A2(n_1603), .B1(n_1628), .B2(n_1629), .C(n_1632), .Y(n_1627) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1600), .Y(n_1693) );
INVxp67_ASAP7_75t_SL g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1606), .B(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1607), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
NAND4xp25_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1627), .C(n_1639), .D(n_1662), .Y(n_1610) );
CKINVDCx14_ASAP7_75t_R g1675 ( .A(n_1612), .Y(n_1675) );
OAI211xp5_ASAP7_75t_SL g1614 ( .A1(n_1615), .A2(n_1617), .B(n_1618), .C(n_1621), .Y(n_1614) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1619), .Y(n_1638) );
O2A1O1Ixp33_ASAP7_75t_L g1662 ( .A1(n_1619), .A2(n_1663), .B(n_1666), .C(n_1668), .Y(n_1662) );
NOR2xp33_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1637), .Y(n_1674) );
O2A1O1Ixp33_ASAP7_75t_L g1668 ( .A1(n_1643), .A2(n_1654), .B(n_1669), .C(n_1670), .Y(n_1668) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1647), .Y(n_1645) );
O2A1O1Ixp33_ASAP7_75t_L g1678 ( .A1(n_1646), .A2(n_1679), .B(n_1682), .C(n_1686), .Y(n_1678) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
INVxp67_ASAP7_75t_SL g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
A2O1A1Ixp33_ASAP7_75t_L g1689 ( .A1(n_1667), .A2(n_1675), .B(n_1690), .C(n_1691), .Y(n_1689) );
INVxp67_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
AOI31xp33_ASAP7_75t_L g1672 ( .A1(n_1673), .A2(n_1675), .A3(n_1676), .B(n_1677), .Y(n_1672) );
INVxp67_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
NOR2xp33_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1694), .Y(n_1692) );
CKINVDCx20_ASAP7_75t_R g1695 ( .A(n_1696), .Y(n_1695) );
CKINVDCx20_ASAP7_75t_R g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1699), .Y(n_1739) );
NOR4xp25_ASAP7_75t_L g1699 ( .A(n_1700), .B(n_1711), .C(n_1729), .D(n_1734), .Y(n_1699) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1708), .Y(n_1701) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
AOI22xp5_ASAP7_75t_L g1715 ( .A1(n_1716), .A2(n_1717), .B1(n_1718), .B2(n_1719), .Y(n_1715) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1731), .B(n_1733), .Y(n_1730) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
CKINVDCx5p33_ASAP7_75t_R g1740 ( .A(n_1741), .Y(n_1740) );
BUFx3_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
BUFx3_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
BUFx4f_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
HB1xp67_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
INVx2_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
OR2x2_ASAP7_75t_L g1753 ( .A(n_1754), .B(n_1775), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1761), .B(n_1764), .Y(n_1760) );
AOI22xp5_ASAP7_75t_L g1768 ( .A1(n_1769), .A2(n_1772), .B1(n_1773), .B2(n_1774), .Y(n_1768) );
INVx2_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
NAND3xp33_ASAP7_75t_SL g1775 ( .A(n_1776), .B(n_1778), .C(n_1780), .Y(n_1775) );
NOR2xp33_ASAP7_75t_SL g1780 ( .A(n_1781), .B(n_1784), .Y(n_1780) );
OAI22xp5_ASAP7_75t_L g1792 ( .A1(n_1790), .A2(n_1793), .B1(n_1794), .B2(n_1795), .Y(n_1792) );
HB1xp67_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
OAI21xp5_ASAP7_75t_L g1800 ( .A1(n_1801), .A2(n_1802), .B(n_1803), .Y(n_1800) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
endmodule