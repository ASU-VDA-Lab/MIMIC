module real_jpeg_29780_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_57;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_58;
wire n_52;
wire n_31;
wire n_9;
wire n_10;
wire n_49;
wire n_63;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_61;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_56;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_28),
.B(n_34),
.Y(n_33)
);

A2O1A1O1Ixp25_ASAP7_75t_L g51 ( 
.A1(n_1),
.A2(n_52),
.B(n_54),
.C(n_55),
.D(n_58),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_52),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_14),
.B1(n_18),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_3),
.A2(n_31),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_4),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_5),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_13)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_5),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_5),
.B(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_6),
.A2(n_14),
.B1(n_18),
.B2(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_41),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_32),
.B(n_40),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_20),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_11),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_19),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_13),
.A2(n_52),
.B(n_56),
.C(n_57),
.Y(n_55)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g60 ( 
.A1(n_17),
.A2(n_18),
.A3(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_23),
.B(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_62),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);


endmodule