module fake_jpeg_2946_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_5),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_46),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_49),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_50),
.B(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_84),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_56),
.B(n_76),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx9p33_ASAP7_75t_R g131 ( 
.A(n_62),
.Y(n_131)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_33),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_82),
.Y(n_105)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_66),
.Y(n_151)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_69),
.Y(n_102)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_35),
.Y(n_77)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_80),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_29),
.B(n_1),
.C(n_3),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_85),
.B(n_39),
.Y(n_136)
);

NAND2x1_ASAP7_75t_SL g86 ( 
.A(n_15),
.B(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_87),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_91),
.Y(n_112)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_90),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_95),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_98),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_12),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_3),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_1),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_15),
.B1(n_40),
.B2(n_38),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_101),
.A2(n_111),
.B1(n_142),
.B2(n_149),
.Y(n_188)
);

OA22x2_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_40),
.B1(n_41),
.B2(n_24),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_103),
.A2(n_143),
.B1(n_7),
.B2(n_9),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_45),
.A2(n_41),
.B1(n_18),
.B2(n_19),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_9),
.B1(n_12),
.B2(n_143),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_15),
.B1(n_38),
.B2(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_116),
.B(n_130),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_39),
.B1(n_36),
.B2(n_32),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_152),
.B1(n_71),
.B2(n_88),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_50),
.B(n_32),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_136),
.A2(n_144),
.B(n_145),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_142)
);

OA22x2_ASAP7_75t_SL g143 ( 
.A1(n_56),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_53),
.B(n_18),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_54),
.B(n_19),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_96),
.A2(n_98),
.B1(n_87),
.B2(n_93),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_79),
.A2(n_16),
.B1(n_4),
.B2(n_6),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_16),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_92),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_157),
.B(n_161),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_158),
.A2(n_201),
.B1(n_109),
.B2(n_108),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_178),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_84),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_170),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_83),
.B1(n_80),
.B2(n_47),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_162),
.A2(n_174),
.B1(n_177),
.B2(n_111),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_68),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_64),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_52),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_117),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_166),
.A2(n_172),
.B1(n_180),
.B2(n_185),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_3),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_173),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_103),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_12),
.B(n_9),
.C(n_10),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_176),
.B(n_194),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_115),
.A2(n_124),
.B1(n_142),
.B2(n_152),
.Y(n_180)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_101),
.B(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_190),
.Y(n_220)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_189),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_107),
.A2(n_118),
.B1(n_122),
.B2(n_149),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_156),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_138),
.B1(n_135),
.B2(n_114),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_197),
.B1(n_167),
.B2(n_181),
.Y(n_213)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_100),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_100),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_195),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_114),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_202),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_140),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_148),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_150),
.A2(n_132),
.B1(n_139),
.B2(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_216),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_235),
.B1(n_207),
.B2(n_206),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_102),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_230),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_186),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_228),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_151),
.B(n_139),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_191),
.B(n_108),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_186),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_102),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_132),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_166),
.A2(n_135),
.B1(n_138),
.B2(n_126),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_235),
.A2(n_187),
.B1(n_208),
.B2(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_252),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_171),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_211),
.B(n_219),
.Y(n_270)
);

OR2x2_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_173),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_257),
.B(n_261),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_160),
.C(n_159),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_247),
.C(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_170),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_173),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_175),
.C(n_190),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_188),
.B1(n_199),
.B2(n_194),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_260),
.B(n_212),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_256),
.B1(n_206),
.B2(n_235),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_222),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_168),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_177),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_208),
.A2(n_188),
.B1(n_185),
.B2(n_176),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_258),
.B1(n_248),
.B2(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_188),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_188),
.B1(n_198),
.B2(n_191),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_263),
.A2(n_265),
.B1(n_266),
.B2(n_225),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_232),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_264),
.B(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_211),
.B1(n_221),
.B2(n_231),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_277),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_227),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_238),
.B(n_250),
.C(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_217),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_279),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_262),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_281),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_245),
.B(n_219),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_282),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_260),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_287),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_227),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_243),
.C(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_243),
.B(n_259),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_246),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_224),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_286),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_295),
.C(n_296),
.Y(n_312)
);

AO22x1_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_238),
.B1(n_251),
.B2(n_248),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_304),
.Y(n_328)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_252),
.C(n_258),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_242),
.C(n_207),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_298),
.B(n_284),
.Y(n_331)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_255),
.B(n_221),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_265),
.B(n_272),
.Y(n_316)
);

AOI22x1_ASAP7_75t_L g304 ( 
.A1(n_267),
.A2(n_255),
.B1(n_254),
.B2(n_256),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_244),
.Y(n_305)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_308),
.B1(n_297),
.B2(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_301),
.B(n_302),
.Y(n_311)
);

NAND2x1_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_293),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_283),
.B1(n_279),
.B2(n_281),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_288),
.B1(n_234),
.B2(n_214),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_295),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_318),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_316),
.B(n_319),
.Y(n_344)
);

A2O1A1O1Ixp25_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_278),
.B(n_270),
.C(n_274),
.D(n_285),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_317),
.B(n_292),
.C(n_330),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_264),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_274),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_272),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_307),
.A2(n_287),
.B1(n_241),
.B2(n_275),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_290),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_241),
.Y(n_329)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_315),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_291),
.A2(n_209),
.B1(n_230),
.B2(n_213),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_303),
.B1(n_291),
.B2(n_304),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_318),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_289),
.C(n_294),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_340),
.C(n_342),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_338),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_298),
.C(n_300),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_303),
.C(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_351),
.B1(n_320),
.B2(n_325),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_292),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_349),
.Y(n_356)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_321),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_363),
.B1(n_343),
.B2(n_347),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_339),
.A2(n_320),
.B1(n_328),
.B2(n_332),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_353),
.B(n_361),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_334),
.B(n_316),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_359),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_337),
.A2(n_328),
.B1(n_311),
.B2(n_313),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_328),
.C(n_327),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_365),
.C(n_341),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_343),
.B1(n_344),
.B2(n_336),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_327),
.C(n_317),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_370),
.C(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_342),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_363),
.A2(n_349),
.B(n_345),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_374),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_358),
.B(n_355),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_373),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_352),
.A2(n_338),
.B1(n_335),
.B2(n_351),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_223),
.C(n_215),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_375),
.B(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_223),
.C(n_215),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_366),
.C(n_222),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_370),
.C(n_375),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_382),
.C(n_226),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_360),
.C(n_356),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_364),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_356),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_386),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_376),
.B(n_222),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_378),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_229),
.A3(n_222),
.B1(n_236),
.B2(n_202),
.C1(n_134),
.C2(n_216),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_388),
.B(n_391),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_216),
.B1(n_214),
.B2(n_236),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_392),
.Y(n_397)
);

AOI322xp5_ASAP7_75t_L g391 ( 
.A1(n_383),
.A2(n_229),
.A3(n_236),
.B1(n_216),
.B2(n_196),
.C1(n_148),
.C2(n_195),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_226),
.C(n_189),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_394),
.B(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_396),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_389),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_216),
.C(n_169),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_399),
.B(n_400),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_393),
.A2(n_183),
.B1(n_184),
.B2(n_126),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_395),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_397),
.A2(n_192),
.B(n_203),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_399),
.B(n_148),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_406),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_407),
.A2(n_402),
.B(n_403),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_401),
.Y(n_409)
);


endmodule