module fake_jpeg_19800_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_0),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_81),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_49),
.B1(n_70),
.B2(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_92),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_63),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_52),
.B(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_110),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_63),
.B1(n_47),
.B2(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_123),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_1),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_117),
.B1(n_69),
.B2(n_8),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_121),
.B(n_124),
.Y(n_128)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_65),
.B1(n_74),
.B2(n_72),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_1),
.CI(n_2),
.CON(n_119),
.SN(n_119)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_4),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_76),
.B1(n_62),
.B2(n_61),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_67),
.B1(n_64),
.B2(n_51),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_2),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_3),
.C(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_135),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_6),
.B(n_10),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_5),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_137),
.A2(n_124),
.B1(n_117),
.B2(n_13),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_138),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_126),
.B(n_133),
.C(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_15),
.Y(n_148)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.C(n_148),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_142),
.B(n_143),
.C(n_140),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_133),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_144),
.B(n_129),
.C(n_21),
.D(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_19),
.B(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_23),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_25),
.B(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_27),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_28),
.Y(n_160)
);


endmodule