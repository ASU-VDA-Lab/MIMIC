module fake_jpeg_2626_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_46),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

BUFx12f_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_50),
.B1(n_55),
.B2(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_47),
.B1(n_55),
.B2(n_50),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_46),
.B1(n_42),
.B2(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_47),
.B1(n_42),
.B2(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_72),
.Y(n_76)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_70),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_88),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_86),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_98),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_97),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_73),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_5),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_19),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_2),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_118),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_22),
.A3(n_23),
.B1(n_26),
.B2(n_29),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_13),
.B(n_14),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_121),
.B(n_100),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_94),
.C(n_20),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_100),
.B(n_101),
.C(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_115),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.C(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_16),
.C(n_21),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_120),
.B1(n_33),
.B2(n_36),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_134),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_131),
.A2(n_40),
.B1(n_126),
.B2(n_130),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_145),
.B(n_125),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_137),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_128),
.Y(n_154)
);

XNOR2x2_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_141),
.Y(n_155)
);


endmodule