module real_aes_5899_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_1100, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_1101, n_1102, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_1100;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_1101;
input n_1102;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_792;
wire n_673;
wire n_386;
wire n_1067;
wire n_518;
wire n_635;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_994;
wire n_495;
wire n_892;
wire n_1072;
wire n_370;
wire n_1078;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_316;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_307;
wire n_500;
wire n_1076;
wire n_463;
wire n_601;
wire n_396;
wire n_661;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_0), .A2(n_570), .B(n_573), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_1), .A2(n_156), .B1(n_426), .B2(n_427), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_2), .A2(n_109), .B1(n_463), .B2(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g593 ( .A(n_3), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_4), .A2(n_7), .B1(n_532), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g674 ( .A(n_5), .Y(n_674) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_6), .Y(n_785) );
AND2x4_ASAP7_75t_L g797 ( .A(n_6), .B(n_798), .Y(n_797) );
AND2x4_ASAP7_75t_L g806 ( .A(n_6), .B(n_289), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_8), .A2(n_155), .B1(n_809), .B2(n_823), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_9), .A2(n_247), .B1(n_413), .B2(n_422), .Y(n_703) );
INVx1_ASAP7_75t_L g712 ( .A(n_10), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_11), .A2(n_192), .B1(n_365), .B2(n_510), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_12), .A2(n_264), .B1(n_420), .B2(n_426), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_13), .A2(n_175), .B1(n_342), .B2(n_346), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_14), .A2(n_117), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_15), .A2(n_152), .B1(n_530), .B2(n_627), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_16), .A2(n_100), .B1(n_1082), .B2(n_1084), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_17), .A2(n_34), .B1(n_422), .B2(n_423), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g1092 ( .A1(n_18), .A2(n_249), .B1(n_468), .B2(n_565), .Y(n_1092) );
INVx1_ASAP7_75t_L g771 ( .A(n_19), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_20), .A2(n_135), .B1(n_308), .B2(n_468), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_21), .Y(n_807) );
INVxp33_ASAP7_75t_SL g833 ( .A(n_22), .Y(n_833) );
AO22x2_ASAP7_75t_L g858 ( .A1(n_23), .A2(n_82), .B1(n_809), .B2(n_823), .Y(n_858) );
AO22x1_ASAP7_75t_L g859 ( .A1(n_24), .A2(n_296), .B1(n_838), .B2(n_844), .Y(n_859) );
INVx1_ASAP7_75t_L g378 ( .A(n_25), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_26), .A2(n_102), .B1(n_413), .B2(n_434), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_27), .A2(n_278), .B1(n_498), .B2(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_28), .B(n_1077), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_29), .A2(n_97), .B1(n_560), .B2(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_30), .A2(n_101), .B1(n_351), .B2(n_358), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_31), .A2(n_173), .B1(n_453), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g753 ( .A(n_32), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_33), .A2(n_1068), .B1(n_1069), .B2(n_1093), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_33), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_35), .A2(n_259), .B1(n_413), .B2(n_414), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_36), .B(n_501), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_37), .A2(n_122), .B1(n_405), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_38), .A2(n_87), .B1(n_455), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_39), .A2(n_292), .B1(n_308), .B2(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g1037 ( .A(n_40), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_41), .A2(n_191), .B1(n_501), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_42), .A2(n_286), .B1(n_466), .B2(n_559), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_43), .A2(n_186), .B1(n_331), .B2(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g630 ( .A(n_44), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_45), .A2(n_98), .B1(n_532), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_46), .A2(n_294), .B1(n_405), .B2(n_651), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_47), .A2(n_148), .B1(n_805), .B2(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g328 ( .A(n_48), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_48), .B(n_223), .Y(n_385) );
INVxp67_ASAP7_75t_L g404 ( .A(n_48), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_49), .A2(n_52), .B1(n_447), .B2(n_710), .C(n_711), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_50), .A2(n_244), .B1(n_504), .B2(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g638 ( .A(n_51), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_53), .A2(n_174), .B1(n_414), .B2(n_423), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_54), .A2(n_237), .B1(n_799), .B2(n_809), .Y(n_812) );
INVx1_ASAP7_75t_L g1024 ( .A(n_54), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_54), .A2(n_1067), .B1(n_1094), .B2(n_1096), .Y(n_1066) );
INVx1_ASAP7_75t_L g596 ( .A(n_55), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_56), .A2(n_149), .B1(n_838), .B2(n_840), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_57), .A2(n_60), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g1090 ( .A1(n_58), .A2(n_234), .B1(n_346), .B2(n_461), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_59), .A2(n_236), .B1(n_466), .B2(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_61), .B(n_313), .Y(n_323) );
INVx1_ASAP7_75t_L g646 ( .A(n_62), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_63), .A2(n_196), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_64), .A2(n_131), .B1(n_455), .B2(n_456), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g548 ( .A1(n_65), .A2(n_390), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g586 ( .A(n_66), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_67), .A2(n_140), .B1(n_535), .B2(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g1027 ( .A(n_68), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_69), .A2(n_268), .B1(n_431), .B2(n_481), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_70), .A2(n_255), .B1(n_823), .B2(n_851), .Y(n_850) );
INVx1_ASAP7_75t_SL g1034 ( .A(n_71), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_72), .A2(n_180), .B1(n_358), .B2(n_466), .Y(n_724) );
INVx2_ASAP7_75t_L g783 ( .A(n_73), .Y(n_783) );
INVxp33_ASAP7_75t_SL g810 ( .A(n_74), .Y(n_810) );
INVx1_ASAP7_75t_L g796 ( .A(n_75), .Y(n_796) );
AND2x4_ASAP7_75t_L g802 ( .A(n_75), .B(n_783), .Y(n_802) );
INVx1_ASAP7_75t_SL g839 ( .A(n_75), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_76), .A2(n_210), .B1(n_542), .B2(n_547), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_77), .A2(n_115), .B1(n_809), .B2(n_823), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_78), .A2(n_218), .B1(n_308), .B2(n_331), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_79), .A2(n_144), .B1(n_416), .B2(n_417), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_80), .A2(n_280), .B1(n_510), .B2(n_539), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_81), .A2(n_170), .B1(n_464), .B2(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g1030 ( .A(n_83), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_84), .A2(n_93), .B1(n_1044), .B2(n_1046), .Y(n_1043) );
INVx1_ASAP7_75t_L g591 ( .A(n_85), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_86), .A2(n_253), .B1(n_363), .B2(n_365), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g1072 ( .A1(n_88), .A2(n_1073), .B(n_1074), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_89), .A2(n_228), .B1(n_346), .B2(n_461), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_90), .A2(n_128), .B1(n_623), .B2(n_624), .Y(n_622) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_91), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_92), .A2(n_142), .B1(n_331), .B2(n_463), .Y(n_725) );
INVx1_ASAP7_75t_L g579 ( .A(n_94), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_95), .B(n_429), .Y(n_428) );
XOR2x2_ASAP7_75t_L g489 ( .A(n_96), .B(n_490), .Y(n_489) );
AO22x2_ASAP7_75t_L g626 ( .A1(n_99), .A2(n_198), .B1(n_627), .B2(n_628), .Y(n_626) );
XOR2x2_ASAP7_75t_L g616 ( .A(n_103), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_104), .A2(n_182), .B1(n_396), .B2(n_481), .Y(n_1039) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_105), .A2(n_205), .B1(n_390), .B2(n_392), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_106), .A2(n_230), .B1(n_416), .B2(n_417), .Y(n_704) );
INVx1_ASAP7_75t_L g314 ( .A(n_107), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_107), .B(n_221), .Y(n_401) );
AOI33xp33_ASAP7_75t_R g512 ( .A1(n_108), .A2(n_254), .A3(n_310), .B1(n_334), .B2(n_513), .B3(n_1100), .Y(n_512) );
INVx1_ASAP7_75t_L g588 ( .A(n_110), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_111), .A2(n_258), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_112), .A2(n_251), .B1(n_683), .B2(n_684), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_113), .A2(n_211), .B1(n_351), .B2(n_530), .Y(n_745) );
AOI21xp5_ASAP7_75t_SL g372 ( .A1(n_114), .A2(n_373), .B(n_377), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_116), .A2(n_265), .B1(n_351), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_118), .A2(n_125), .B1(n_426), .B2(n_432), .Y(n_697) );
XNOR2x2_ASAP7_75t_L g439 ( .A(n_119), .B(n_440), .Y(n_439) );
XOR2xp5_ASAP7_75t_L g517 ( .A(n_119), .B(n_440), .Y(n_517) );
INVx1_ASAP7_75t_L g693 ( .A(n_120), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_121), .Y(n_407) );
AO221x2_ASAP7_75t_L g791 ( .A1(n_121), .A2(n_129), .B1(n_792), .B2(n_799), .C(n_803), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_123), .A2(n_282), .B1(n_365), .B2(n_463), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_124), .A2(n_226), .B1(n_419), .B2(n_420), .Y(n_702) );
INVx1_ASAP7_75t_L g526 ( .A(n_126), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_126), .A2(n_293), .B1(n_794), .B2(n_823), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_127), .A2(n_233), .B1(n_510), .B2(n_539), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_130), .A2(n_257), .B1(n_468), .B2(n_679), .Y(n_1042) );
AOI21xp33_ASAP7_75t_L g751 ( .A1(n_132), .A2(n_431), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g436 ( .A(n_133), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_134), .A2(n_434), .B(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_136), .A2(n_284), .B1(n_419), .B2(n_420), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_137), .A2(n_166), .B1(n_346), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_138), .A2(n_158), .B1(n_537), .B2(n_565), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_139), .A2(n_176), .B1(n_434), .B2(n_479), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_141), .A2(n_225), .B1(n_396), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_143), .A2(n_208), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_145), .A2(n_209), .B1(n_422), .B2(n_423), .Y(n_421) );
AO22x1_ASAP7_75t_L g717 ( .A1(n_146), .A2(n_147), .B1(n_461), .B2(n_565), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g773 ( .A(n_150), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_151), .A2(n_172), .B1(n_416), .B2(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_153), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_154), .A2(n_161), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_157), .A2(n_177), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_159), .A2(n_276), .B1(n_358), .B2(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g640 ( .A(n_160), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_162), .A2(n_227), .B1(n_838), .B2(n_840), .Y(n_837) );
INVx1_ASAP7_75t_L g574 ( .A(n_163), .Y(n_574) );
INVx1_ASAP7_75t_L g635 ( .A(n_164), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_165), .A2(n_241), .B1(n_405), .B2(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_167), .A2(n_189), .B1(n_606), .B2(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g707 ( .A(n_168), .Y(n_707) );
OAI222xp33_ASAP7_75t_L g718 ( .A1(n_168), .A2(n_719), .B1(n_724), .B2(n_725), .C1(n_1101), .C2(n_1102), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_168), .B(n_725), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_169), .A2(n_274), .B1(n_414), .B2(n_419), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_171), .A2(n_256), .B1(n_679), .B2(n_681), .Y(n_678) );
XOR2xp5_ASAP7_75t_L g472 ( .A(n_178), .B(n_473), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g516 ( .A(n_178), .B(n_473), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_179), .A2(n_291), .B1(n_342), .B2(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g1026 ( .A(n_181), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_183), .A2(n_217), .B1(n_363), .B2(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_184), .B(n_456), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_185), .A2(n_267), .B1(n_453), .B2(n_501), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_187), .A2(n_195), .B1(n_723), .B2(n_1080), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_188), .A2(n_235), .B1(n_479), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_190), .A2(n_199), .B1(n_432), .B2(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_193), .A2(n_447), .B(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_194), .A2(n_239), .B1(n_346), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_197), .A2(n_215), .B1(n_794), .B2(n_805), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_200), .A2(n_224), .B1(n_405), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_201), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g1075 ( .A(n_202), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_203), .B(n_499), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_204), .A2(n_295), .B1(n_468), .B2(n_565), .Y(n_564) );
OA22x2_ASAP7_75t_L g318 ( .A1(n_206), .A2(n_223), .B1(n_313), .B2(n_317), .Y(n_318) );
INVx1_ASAP7_75t_L g338 ( .A(n_206), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_207), .A2(n_281), .B1(n_429), .B2(n_499), .Y(n_698) );
AO22x2_ASAP7_75t_L g580 ( .A1(n_212), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_212), .Y(n_581) );
INVx1_ASAP7_75t_L g828 ( .A(n_213), .Y(n_828) );
NAND2xp33_ASAP7_75t_L g764 ( .A(n_214), .B(n_369), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_216), .A2(n_273), .B1(n_365), .B2(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_219), .A2(n_266), .B1(n_392), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_220), .A2(n_238), .B1(n_794), .B2(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g330 ( .A(n_221), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_221), .B(n_336), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_222), .A2(n_250), .B1(n_431), .B2(n_432), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g339 ( .A1(n_223), .A2(n_243), .B(n_340), .Y(n_339) );
XNOR2x1_ASAP7_75t_L g409 ( .A(n_227), .B(n_410), .Y(n_409) );
XNOR2x2_ASAP7_75t_SL g437 ( .A(n_227), .B(n_410), .Y(n_437) );
INVx1_ASAP7_75t_L g661 ( .A(n_229), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_231), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g738 ( .A(n_232), .Y(n_738) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_240), .Y(n_1058) );
INVx1_ASAP7_75t_SL g829 ( .A(n_242), .Y(n_829) );
INVx1_ASAP7_75t_L g316 ( .A(n_243), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_243), .B(n_279), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_245), .A2(n_270), .B1(n_510), .B2(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_246), .B(n_431), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_248), .Y(n_1055) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_252), .A2(n_670), .B(n_673), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_260), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_261), .A2(n_275), .B1(n_351), .B2(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_262), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_263), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g550 ( .A(n_269), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_271), .A2(n_285), .B1(n_447), .B2(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g1051 ( .A(n_272), .Y(n_1051) );
AOI22x1_ASAP7_75t_L g395 ( .A1(n_277), .A2(n_288), .B1(n_396), .B2(n_405), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_279), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g643 ( .A(n_283), .Y(n_643) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_287), .Y(n_1052) );
INVx1_ASAP7_75t_L g798 ( .A(n_289), .Y(n_798) );
INVx1_ASAP7_75t_L g644 ( .A(n_290), .Y(n_644) );
AOI31xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_774), .A3(n_777), .B(n_786), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_518), .B(n_655), .C(n_657), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_300), .B(n_519), .Y(n_656) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_300), .A2(n_656), .B(n_775), .C(n_776), .Y(n_774) );
XNOR2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_438), .Y(n_300) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_408), .B2(n_437), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
XNOR2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_407), .Y(n_304) );
NOR3xp33_ASAP7_75t_SL g305 ( .A(n_306), .B(n_349), .C(n_367), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_341), .Y(n_306) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_308), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx8_ASAP7_75t_L g565 ( .A(n_309), .Y(n_565) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_319), .Y(n_309) );
AND2x4_ASAP7_75t_L g343 ( .A(n_310), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g371 ( .A(n_310), .B(n_360), .Y(n_371) );
AND2x2_ASAP7_75t_L g406 ( .A(n_310), .B(n_356), .Y(n_406) );
AND2x4_ASAP7_75t_L g413 ( .A(n_310), .B(n_319), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_310), .B(n_348), .Y(n_414) );
AND2x4_ASAP7_75t_L g426 ( .A(n_310), .B(n_356), .Y(n_426) );
AND2x2_ASAP7_75t_L g431 ( .A(n_310), .B(n_360), .Y(n_431) );
AND2x2_ASAP7_75t_L g536 ( .A(n_310), .B(n_319), .Y(n_536) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_318), .Y(n_310) );
INVx1_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g317 ( .A(n_313), .Y(n_317) );
INVx3_ASAP7_75t_L g322 ( .A(n_313), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g329 ( .A(n_313), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_314), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g403 ( .A1(n_316), .A2(n_340), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g355 ( .A(n_318), .Y(n_355) );
AND2x2_ASAP7_75t_L g376 ( .A(n_318), .B(n_354), .Y(n_376) );
AND2x2_ASAP7_75t_L g402 ( .A(n_318), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g333 ( .A(n_319), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g364 ( .A(n_319), .B(n_353), .Y(n_364) );
AND2x4_ASAP7_75t_L g419 ( .A(n_319), .B(n_353), .Y(n_419) );
AND2x4_ASAP7_75t_L g422 ( .A(n_319), .B(n_334), .Y(n_422) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_319), .Y(n_513) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
OR2x2_ASAP7_75t_L g345 ( .A(n_320), .B(n_325), .Y(n_345) );
AND2x4_ASAP7_75t_L g356 ( .A(n_320), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
AND2x2_ASAP7_75t_L g399 ( .A(n_320), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_322), .B(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g336 ( .A(n_322), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_323), .B(n_335), .C(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g357 ( .A(n_326), .Y(n_357) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx4_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx4_ASAP7_75t_L g468 ( .A(n_332), .Y(n_468) );
INVx4_ASAP7_75t_L g537 ( .A(n_332), .Y(n_537) );
INVx2_ASAP7_75t_SL g744 ( .A(n_332), .Y(n_744) );
INVx2_ASAP7_75t_L g762 ( .A(n_332), .Y(n_762) );
INVx8_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g347 ( .A(n_334), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g394 ( .A(n_334), .B(n_360), .Y(n_394) );
AND2x4_ASAP7_75t_L g423 ( .A(n_334), .B(n_348), .Y(n_423) );
AND2x4_ASAP7_75t_L g432 ( .A(n_334), .B(n_360), .Y(n_432) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
BUFx12f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_343), .Y(n_461) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_343), .Y(n_506) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_343), .Y(n_532) );
BUFx3_ASAP7_75t_L g683 ( .A(n_343), .Y(n_683) );
AND2x4_ASAP7_75t_L g420 ( .A(n_344), .B(n_353), .Y(n_420) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g348 ( .A(n_345), .Y(n_348) );
BUFx3_ASAP7_75t_L g624 ( .A(n_346), .Y(n_624) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx6_ASAP7_75t_L g505 ( .A(n_347), .Y(n_505) );
AND2x4_ASAP7_75t_L g366 ( .A(n_348), .B(n_353), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_362), .Y(n_349) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_351), .Y(n_1057) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_352), .Y(n_466) );
INVx3_ASAP7_75t_L g610 ( .A(n_352), .Y(n_610) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_353), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g416 ( .A(n_353), .B(n_356), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_353), .B(n_360), .Y(n_417) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
AND2x4_ASAP7_75t_L g375 ( .A(n_356), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g434 ( .A(n_356), .B(n_376), .Y(n_434) );
AND2x4_ASAP7_75t_L g360 ( .A(n_357), .B(n_361), .Y(n_360) );
BUFx5_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx3_ASAP7_75t_L g508 ( .A(n_359), .Y(n_508) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_359), .Y(n_530) );
INVx1_ASAP7_75t_L g561 ( .A(n_359), .Y(n_561) );
AND2x4_ASAP7_75t_L g391 ( .A(n_360), .B(n_376), .Y(n_391) );
AND2x2_ASAP7_75t_L g429 ( .A(n_360), .B(n_376), .Y(n_429) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_364), .Y(n_463) );
BUFx12f_ASAP7_75t_L g510 ( .A(n_364), .Y(n_510) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_366), .Y(n_464) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_366), .Y(n_511) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_366), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g367 ( .A(n_368), .B(n_372), .C(n_389), .D(n_395), .Y(n_367) );
INVx3_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g544 ( .A(n_370), .Y(n_544) );
INVx2_ASAP7_75t_L g572 ( .A(n_370), .Y(n_572) );
INVx2_ASAP7_75t_L g672 ( .A(n_370), .Y(n_672) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g445 ( .A(n_371), .Y(n_445) );
BUFx3_ASAP7_75t_L g598 ( .A(n_371), .Y(n_598) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_375), .Y(n_447) );
BUFx3_ASAP7_75t_L g493 ( .A(n_375), .Y(n_493) );
BUFx3_ASAP7_75t_L g547 ( .A(n_375), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_379), .B(n_753), .Y(n_752) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_380), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g481 ( .A(n_380), .Y(n_481) );
INVx2_ASAP7_75t_L g499 ( .A(n_380), .Y(n_499) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_380), .Y(n_601) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g458 ( .A(n_381), .Y(n_458) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_387), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_383), .B(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_384), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx8_ASAP7_75t_SL g452 ( .A(n_391), .Y(n_452) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_391), .Y(n_476) );
BUFx3_ASAP7_75t_L g501 ( .A(n_391), .Y(n_501) );
INVx2_ASAP7_75t_L g578 ( .A(n_391), .Y(n_578) );
INVx2_ASAP7_75t_L g1033 ( .A(n_391), .Y(n_1033) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g453 ( .A(n_393), .Y(n_453) );
INVx2_ASAP7_75t_L g494 ( .A(n_393), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_393), .A2(n_592), .B1(n_643), .B2(n_644), .Y(n_642) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_394), .Y(n_542) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_394), .Y(n_723) );
INVx4_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g455 ( .A(n_397), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_397), .A2(n_574), .B(n_575), .Y(n_573) );
INVx2_ASAP7_75t_L g768 ( .A(n_397), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g1074 ( .A1(n_397), .A2(n_1075), .B(n_1076), .Y(n_1074) );
INVx5_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g496 ( .A(n_398), .Y(n_496) );
BUFx4f_ASAP7_75t_L g651 ( .A(n_398), .Y(n_651) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
AND2x4_ASAP7_75t_L g427 ( .A(n_399), .B(n_402), .Y(n_427) );
AND2x2_ASAP7_75t_L g479 ( .A(n_399), .B(n_402), .Y(n_479) );
INVx3_ASAP7_75t_L g589 ( .A(n_405), .Y(n_589) );
BUFx3_ASAP7_75t_L g668 ( .A(n_405), .Y(n_668) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
BUFx3_ASAP7_75t_L g721 ( .A(n_406), .Y(n_721) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_424), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .C(n_418), .D(n_421), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .C(n_430), .D(n_433), .Y(n_424) );
BUFx3_ASAP7_75t_L g522 ( .A(n_437), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_469), .B1(n_470), .B2(n_517), .Y(n_438) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_459), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .C(n_451), .D(n_454), .Y(n_441) );
INVx1_ASAP7_75t_L g1038 ( .A(n_443), .Y(n_1038) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g498 ( .A(n_445), .Y(n_498) );
INVx4_ASAP7_75t_L g639 ( .A(n_447), .Y(n_639) );
INVx1_ASAP7_75t_L g1028 ( .A(n_448), .Y(n_1028) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g568 ( .A(n_449), .Y(n_568) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_449), .Y(n_641) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g1086 ( .A(n_450), .Y(n_1086) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_457), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g652 ( .A(n_457), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_457), .B(n_712), .Y(n_711) );
INVx4_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g1078 ( .A(n_458), .Y(n_1078) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .C(n_465), .D(n_467), .Y(n_459) );
BUFx3_ASAP7_75t_L g634 ( .A(n_464), .Y(n_634) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AO22x1_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_487), .B1(n_488), .B2(n_514), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .C(n_478), .D(n_480), .Y(n_474) );
INVx2_ASAP7_75t_L g592 ( .A(n_476), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .C(n_485), .D(n_486), .Y(n_482) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .C(n_497), .D(n_500), .Y(n_491) );
INVx1_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
BUFx2_ASAP7_75t_L g667 ( .A(n_493), .Y(n_667) );
BUFx3_ASAP7_75t_L g1073 ( .A(n_498), .Y(n_1073) );
INVx3_ASAP7_75t_L g772 ( .A(n_499), .Y(n_772) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .C(n_509), .D(n_512), .Y(n_502) );
INVx5_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g612 ( .A(n_505), .Y(n_612) );
INVx2_ASAP7_75t_L g685 ( .A(n_505), .Y(n_685) );
INVx1_ASAP7_75t_L g716 ( .A(n_505), .Y(n_716) );
INVx2_ASAP7_75t_L g742 ( .A(n_505), .Y(n_742) );
BUFx3_ASAP7_75t_L g623 ( .A(n_506), .Y(n_623) );
BUFx2_ASAP7_75t_L g688 ( .A(n_508), .Y(n_688) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_510), .Y(n_632) );
INVx1_ASAP7_75t_L g680 ( .A(n_510), .Y(n_680) );
BUFx12f_ASAP7_75t_L g1089 ( .A(n_510), .Y(n_1089) );
INVx1_ASAP7_75t_L g1045 ( .A(n_511), .Y(n_1045) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g775 ( .A(n_518), .Y(n_775) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AO22x1_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_553), .B2(n_654), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_551), .B2(n_552), .Y(n_521) );
INVx2_ASAP7_75t_L g551 ( .A(n_522), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_523), .Y(n_552) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
XNOR2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
NOR4xp75_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .C(n_540), .D(n_545), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
BUFx2_ASAP7_75t_SL g628 ( .A(n_530), .Y(n_628) );
INVx1_ASAP7_75t_L g1059 ( .A(n_530), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_536), .Y(n_606) );
BUFx2_ASAP7_75t_L g621 ( .A(n_537), .Y(n_621) );
BUFx3_ASAP7_75t_L g681 ( .A(n_539), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx3_ASAP7_75t_L g594 ( .A(n_542), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_548), .Y(n_545) );
INVx2_ASAP7_75t_L g1083 ( .A(n_547), .Y(n_1083) );
INVx2_ASAP7_75t_L g654 ( .A(n_553), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_615), .B1(n_616), .B2(n_653), .Y(n_553) );
INVx1_ASAP7_75t_L g653 ( .A(n_554), .Y(n_653) );
AO22x2_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_580), .B1(n_613), .B2(n_614), .Y(n_554) );
INVx1_ASAP7_75t_L g613 ( .A(n_555), .Y(n_613) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_579), .Y(n_555) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_566), .Y(n_556) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .C(n_563), .D(n_564), .Y(n_557) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .C(n_576), .Y(n_566) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g1080 ( .A(n_578), .Y(n_1080) );
INVx2_ASAP7_75t_L g614 ( .A(n_580), .Y(n_614) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_602), .Y(n_583) );
NOR3xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_590), .C(n_595), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g665 ( .A(n_592), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_599), .Y(n_595) );
INVx2_ASAP7_75t_L g710 ( .A(n_597), .Y(n_710) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g649 ( .A(n_598), .Y(n_649) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g627 ( .A(n_610), .Y(n_627) );
INVx1_ASAP7_75t_L g687 ( .A(n_610), .Y(n_687) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_625), .C(n_636), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
OAI22x1_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_631), .B1(n_633), .B2(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR3xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_642), .C(n_645), .Y(n_636) );
OAI22xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_639), .A2(n_1026), .B1(n_1027), .B2(n_1028), .Y(n_1025) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_SL g675 ( .A(n_651), .Y(n_675) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g776 ( .A(n_657), .Y(n_776) );
XNOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_734), .Y(n_657) );
AO22x2_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_690), .B2(n_733), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
XNOR2x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_677), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_666), .C(n_669), .Y(n_663) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_676), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_682), .C(n_686), .D(n_689), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g1053 ( .A(n_683), .Y(n_1053) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g733 ( .A(n_690), .Y(n_733) );
XNOR2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_705), .Y(n_690) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
XNOR2x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
OR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .C(n_698), .D(n_699), .Y(n_695) );
NAND4xp25_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .C(n_703), .D(n_704), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_706), .B(n_726), .Y(n_705) );
AOI21x1_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B(n_718), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_713), .Y(n_708) );
BUFx2_ASAP7_75t_L g727 ( .A(n_709), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g731 ( .A(n_715), .B(n_724), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_717), .Y(n_732) );
INVx1_ASAP7_75t_L g730 ( .A(n_719), .Y(n_730) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx4_ASAP7_75t_L g1035 ( .A(n_723), .Y(n_1035) );
NAND4xp75_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .C(n_731), .D(n_732), .Y(n_726) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
XOR2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_754), .Y(n_735) );
XNOR2x1_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_740), .B(n_747), .Y(n_739) );
NAND4xp25_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .C(n_745), .D(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g1047 ( .A(n_742), .Y(n_1047) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .C(n_750), .D(n_751), .Y(n_747) );
XNOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_773), .Y(n_754) );
NAND4xp75_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .C(n_763), .D(n_766), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
BUFx10_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .C(n_785), .Y(n_780) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_781), .B(n_1064), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_781), .B(n_1065), .Y(n_1095) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OA21x2_ASAP7_75t_L g1097 ( .A1(n_782), .A2(n_839), .B(n_1098), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g795 ( .A(n_783), .B(n_796), .Y(n_795) );
AND3x4_ASAP7_75t_L g838 ( .A(n_783), .B(n_797), .C(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g1064 ( .A(n_784), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_785), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_1019), .B1(n_1020), .B2(n_1062), .C(n_1066), .Y(n_786) );
NOR3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_941), .C(n_981), .Y(n_787) );
OAI211xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_814), .B(n_881), .C(n_915), .Y(n_788) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_811), .Y(n_790) );
INVx2_ASAP7_75t_L g886 ( .A(n_791), .Y(n_886) );
HB1xp67_ASAP7_75t_SL g887 ( .A(n_791), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_791), .B(n_890), .Y(n_934) );
AOI31xp33_ASAP7_75t_L g941 ( .A1(n_791), .A2(n_942), .A3(n_947), .B(n_974), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_791), .B(n_868), .Y(n_1008) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_793), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
AND2x4_ASAP7_75t_L g805 ( .A(n_795), .B(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g840 ( .A(n_795), .B(n_806), .Y(n_840) );
AND2x2_ASAP7_75t_L g844 ( .A(n_795), .B(n_806), .Y(n_844) );
AND2x4_ASAP7_75t_L g801 ( .A(n_797), .B(n_802), .Y(n_801) );
AND2x4_ASAP7_75t_L g823 ( .A(n_797), .B(n_802), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_797), .B(n_802), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g1098 ( .A(n_797), .Y(n_1098) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
AND2x4_ASAP7_75t_L g809 ( .A(n_802), .B(n_806), .Y(n_809) );
AND2x2_ASAP7_75t_L g821 ( .A(n_802), .B(n_806), .Y(n_821) );
AND2x2_ASAP7_75t_L g851 ( .A(n_802), .B(n_806), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B1(n_808), .B2(n_810), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_804), .A2(n_808), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g891 ( .A(n_811), .Y(n_891) );
OR2x2_ASAP7_75t_L g914 ( .A(n_811), .B(n_856), .Y(n_914) );
AND2x2_ASAP7_75t_L g956 ( .A(n_811), .B(n_931), .Y(n_956) );
OR2x2_ASAP7_75t_L g986 ( .A(n_811), .B(n_987), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_846), .B1(n_853), .B2(n_860), .C(n_861), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_824), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_817), .B(n_835), .Y(n_860) );
AND2x2_ASAP7_75t_L g879 ( .A(n_817), .B(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g895 ( .A(n_817), .B(n_835), .Y(n_895) );
AND2x2_ASAP7_75t_L g908 ( .A(n_817), .B(n_885), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_817), .B(n_842), .Y(n_965) );
NOR3xp33_ASAP7_75t_L g1017 ( .A(n_817), .B(n_918), .C(n_994), .Y(n_1017) );
INVx3_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx3_ASAP7_75t_L g864 ( .A(n_819), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_819), .B(n_854), .Y(n_877) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_819), .B(n_842), .Y(n_1014) );
AND2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_834), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g867 ( .A(n_825), .B(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_825), .B(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_825), .B(n_890), .Y(n_898) );
INVx1_ASAP7_75t_L g909 ( .A(n_825), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_825), .B(n_929), .Y(n_963) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g854 ( .A(n_826), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_826), .B(n_849), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_826), .B(n_864), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_826), .B(n_857), .Y(n_951) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_826), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_826), .B(n_849), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_826), .B(n_848), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_826), .B(n_892), .Y(n_1015) );
OR2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_830), .Y(n_826) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_832), .Y(n_1019) );
INVx1_ASAP7_75t_L g875 ( .A(n_834), .Y(n_875) );
OAI221xp5_ASAP7_75t_SL g888 ( .A1(n_834), .A2(n_889), .B1(n_893), .B2(n_894), .C(n_896), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_834), .B(n_905), .Y(n_990) );
OR2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_842), .Y(n_834) );
AND2x2_ASAP7_75t_L g880 ( .A(n_835), .B(n_842), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_835), .B(n_864), .Y(n_930) );
OR2x2_ASAP7_75t_L g973 ( .A(n_835), .B(n_864), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_835), .B(n_998), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
OR2x2_ASAP7_75t_L g863 ( .A(n_836), .B(n_842), .Y(n_863) );
AND2x2_ASAP7_75t_L g885 ( .A(n_836), .B(n_842), .Y(n_885) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_841), .Y(n_836) );
AOI322xp5_ASAP7_75t_L g896 ( .A1(n_842), .A2(n_869), .A3(n_890), .B1(n_897), .B2(n_899), .C1(n_900), .C2(n_903), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_842), .B(n_864), .Y(n_919) );
INVx1_ASAP7_75t_L g924 ( .A(n_842), .Y(n_924) );
AND2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g899 ( .A(n_847), .Y(n_899) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g866 ( .A(n_848), .B(n_857), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
OR2x2_ASAP7_75t_L g856 ( .A(n_849), .B(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g870 ( .A(n_849), .Y(n_870) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_849), .Y(n_872) );
AND2x2_ASAP7_75t_L g892 ( .A(n_849), .B(n_857), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_849), .B(n_921), .Y(n_920) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_849), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_849), .B(n_854), .Y(n_971) );
AND2x4_ASAP7_75t_L g849 ( .A(n_850), .B(n_852), .Y(n_849) );
AND2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
INVx1_ASAP7_75t_SL g918 ( .A(n_854), .Y(n_918) );
AND2x2_ASAP7_75t_L g946 ( .A(n_854), .B(n_880), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_855), .A2(n_907), .B1(n_911), .B2(n_914), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_855), .A2(n_943), .B(n_944), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_855), .B(n_879), .Y(n_966) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
CKINVDCx6p67_ASAP7_75t_R g869 ( .A(n_857), .Y(n_869) );
AOI321xp33_ASAP7_75t_L g881 ( .A1(n_857), .A2(n_882), .A3(n_886), .B1(n_887), .B2(n_888), .C(n_906), .Y(n_881) );
OR2x2_ASAP7_75t_L g921 ( .A(n_857), .B(n_891), .Y(n_921) );
INVx1_ASAP7_75t_L g932 ( .A(n_857), .Y(n_932) );
OR2x6_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_864), .B1(n_865), .B2(n_867), .C(n_871), .Y(n_861) );
INVx1_ASAP7_75t_L g959 ( .A(n_862), .Y(n_959) );
OR2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_863), .B(n_877), .Y(n_926) );
INVx1_ASAP7_75t_L g938 ( .A(n_863), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_863), .B(n_989), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_863), .B(n_901), .Y(n_1018) );
AND2x2_ASAP7_75t_L g884 ( .A(n_864), .B(n_885), .Y(n_884) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_864), .Y(n_913) );
AND2x2_ASAP7_75t_L g937 ( .A(n_864), .B(n_938), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_864), .B(n_946), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_864), .B(n_875), .Y(n_976) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_866), .B(n_890), .Y(n_893) );
AOI32xp33_ASAP7_75t_L g1016 ( .A1(n_866), .A2(n_897), .A3(n_972), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_868), .B(n_918), .Y(n_923) );
INVx1_ASAP7_75t_L g927 ( .A(n_868), .Y(n_927) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_869), .B(n_891), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_870), .B(n_945), .Y(n_944) );
AND2x2_ASAP7_75t_L g992 ( .A(n_870), .B(n_891), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_878), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
AND2x2_ASAP7_75t_L g983 ( .A(n_879), .B(n_970), .Y(n_983) );
AND2x2_ASAP7_75t_L g903 ( .A(n_880), .B(n_904), .Y(n_903) );
AND2x2_ASAP7_75t_L g912 ( .A(n_880), .B(n_913), .Y(n_912) );
AOI211xp5_ASAP7_75t_L g947 ( .A1(n_880), .A2(n_948), .B(n_949), .C(n_960), .Y(n_947) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g1009 ( .A(n_884), .Y(n_1009) );
INVx1_ASAP7_75t_L g901 ( .A(n_885), .Y(n_901) );
AND2x2_ASAP7_75t_L g943 ( .A(n_885), .B(n_904), .Y(n_943) );
INVx1_ASAP7_75t_L g910 ( .A(n_886), .Y(n_910) );
INVxp67_ASAP7_75t_L g1002 ( .A(n_887), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .Y(n_889) );
INVx5_ASAP7_75t_L g940 ( .A(n_890), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_890), .B(n_958), .Y(n_980) );
NOR3xp33_ASAP7_75t_L g1000 ( .A(n_890), .B(n_901), .C(n_1001), .Y(n_1000) );
INVx3_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AND2x2_ASAP7_75t_L g995 ( .A(n_891), .B(n_931), .Y(n_995) );
INVx2_ASAP7_75t_L g987 ( .A(n_892), .Y(n_987) );
INVx1_ASAP7_75t_L g948 ( .A(n_893), .Y(n_948) );
CKINVDCx16_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
A2O1A1Ixp33_ASAP7_75t_SL g982 ( .A1(n_899), .A2(n_931), .B(n_975), .C(n_983), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g939 ( .A(n_902), .Y(n_939) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_903), .B(n_958), .Y(n_1012) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .C(n_910), .Y(n_907) );
INVx1_ASAP7_75t_L g954 ( .A(n_908), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_909), .B(n_959), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_911), .B(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_920), .B1(n_922), .B2(n_933), .C(n_935), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_918), .B(n_929), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g960 ( .A1(n_921), .A2(n_961), .B(n_966), .C(n_967), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_921), .A2(n_928), .B1(n_986), .B2(n_1011), .Y(n_1010) );
OAI222xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_924), .B1(n_925), .B2(n_927), .C1(n_928), .C2(n_931), .Y(n_922) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_931), .B(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g936 ( .A(n_937), .B(n_939), .C(n_940), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_952), .B1(n_955), .B2(n_957), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_954), .A2(n_994), .B1(n_996), .B2(n_997), .C(n_999), .Y(n_993) );
A2O1A1Ixp33_ASAP7_75t_L g1013 ( .A1(n_954), .A2(n_1014), .B(n_1015), .C(n_1016), .Y(n_1013) );
A2O1A1Ixp33_ASAP7_75t_L g1004 ( .A1(n_955), .A2(n_980), .B(n_1005), .C(n_1006), .Y(n_1004) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_958), .B(n_965), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g961 ( .A(n_962), .B(n_964), .Y(n_961) );
INVxp33_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVxp67_ASAP7_75t_SL g967 ( .A(n_968), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_972), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
OAI21xp33_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_977), .B(n_979), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
A2O1A1Ixp33_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_984), .B(n_1002), .C(n_1003), .Y(n_981) );
AOI221xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_988), .B1(n_990), .B2(n_991), .C(n_993), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g1005 ( .A(n_990), .Y(n_1005) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
NOR3xp33_ASAP7_75t_SL g1003 ( .A(n_1004), .B(n_1010), .C(n_1013), .Y(n_1003) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NOR2xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
INVxp67_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
AO22x2_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1023), .B1(n_1040), .B2(n_1060), .Y(n_1021) );
NOR4xp25_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1025), .C(n_1029), .D(n_1036), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_1024), .Y(n_1023) );
NOR3xp33_ASAP7_75t_SL g1061 ( .A(n_1025), .B(n_1029), .C(n_1036), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1031), .B1(n_1034), .B2(n_1035), .Y(n_1029) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_1033), .Y(n_1032) );
OAI21xp33_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1038), .B(n_1039), .Y(n_1036) );
NAND2xp5_ASAP7_75t_SL g1060 ( .A(n_1040), .B(n_1061), .Y(n_1060) );
NOR3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1048), .C(n_1054), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1051), .B1(n_1052), .B2(n_1053), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
OAI22x1_ASAP7_75t_SL g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1058), .B2(n_1059), .Y(n_1054) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1069), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1087), .Y(n_1070) );
NAND3xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1079), .C(n_1081), .Y(n_1071) );
INVx4_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NAND4xp25_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1090), .C(n_1091), .D(n_1092), .Y(n_1087) );
BUFx2_ASAP7_75t_SL g1094 ( .A(n_1095), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
endmodule