module fake_jpeg_10120_n_19 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_19;

wire n_13;
wire n_14;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

AOI22xp33_ASAP7_75t_L g11 ( 
.A1(n_6),
.A2(n_3),
.B1(n_9),
.B2(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_10),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_0),
.B(n_1),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_7),
.A2(n_4),
.B1(n_2),
.B2(n_8),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

AOI21x1_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_16),
.B(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_4),
.B1(n_11),
.B2(n_14),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_12),
.C(n_13),
.Y(n_19)
);


endmodule