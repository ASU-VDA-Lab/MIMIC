module fake_jpeg_2628_n_231 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_231);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.Y(n_98)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_81),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_79),
.B1(n_59),
.B2(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_78),
.B1(n_62),
.B2(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_78),
.B1(n_62),
.B2(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_71),
.B1(n_69),
.B2(n_75),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_71),
.B1(n_69),
.B2(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_69),
.B1(n_85),
.B2(n_75),
.Y(n_110)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_84),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_85),
.B1(n_82),
.B2(n_57),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_132),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_137),
.Y(n_159)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_4),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_72),
.A3(n_63),
.B1(n_70),
.B2(n_56),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_64),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_83),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

CKINVDCx9p33_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_142),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_53),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_117),
.B1(n_109),
.B2(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_143),
.A2(n_161),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_103),
.B1(n_109),
.B2(n_101),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_64),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_128),
.B(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_52),
.C(n_49),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_153),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_48),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_3),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_46),
.B1(n_45),
.B2(n_41),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_130),
.B1(n_122),
.B2(n_128),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_7),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_6),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_27),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_39),
.C(n_38),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_29),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_122),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_168),
.C(n_152),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_153),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_174),
.B(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_123),
.B(n_37),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_178),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_172),
.B(n_177),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_123),
.B(n_34),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_155),
.B(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_165),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_190),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_192),
.C(n_179),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_185),
.B(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_195),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_28),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_24),
.C(n_10),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_196),
.B1(n_176),
.B2(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_9),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_202),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_206),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_167),
.B(n_169),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_14),
.B(n_15),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_190),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_173),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_176),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_213),
.C(n_218),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_16),
.C(n_17),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_202),
.B1(n_207),
.B2(n_200),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_216),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_217),
.A3(n_218),
.B1(n_200),
.B2(n_213),
.C(n_21),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_224),
.B(n_219),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_221),
.C(n_19),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_18),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_20),
.C(n_22),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_20),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_22),
.Y(n_231)
);


endmodule