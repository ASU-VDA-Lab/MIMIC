module fake_ariane_556_n_492 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_492);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_492;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_139;
wire n_391;
wire n_349;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_401;
wire n_485;
wire n_267;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_247;
wire n_369;
wire n_240;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_478;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_163;
wire n_141;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_468;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_252;
wire n_215;
wire n_161;
wire n_454;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;

INVx2_ASAP7_75t_SL g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_18),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_44),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_20),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_13),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_67),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_81),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_51),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_38),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

BUFx2_ASAP7_75t_SL g163 ( 
.A(n_91),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_27),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_47),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_15),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_6),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_43),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_35),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_48),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_71),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_21),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_22),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_90),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_33),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_50),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_64),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_87),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_39),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_108),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_25),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_74),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_36),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_23),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_84),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_94),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_63),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_4),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_9),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_143),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_150),
.B(n_205),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_139),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_137),
.B(n_158),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

CKINVDCx8_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_147),
.B(n_0),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_148),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_168),
.B(n_1),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_152),
.B(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_156),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_161),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_162),
.B(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_166),
.A2(n_186),
.B1(n_204),
.B2(n_187),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_172),
.B(n_5),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_150),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_205),
.Y(n_251)
);

AO22x2_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_187),
.B1(n_134),
.B2(n_190),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_151),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_173),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_174),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_175),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_177),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_151),
.Y(n_267)
);

INVx3_ASAP7_75t_R g268 ( 
.A(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_179),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_217),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_181),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_182),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_185),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_192),
.B1(n_188),
.B2(n_209),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_239),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_260),
.B(n_235),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_244),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_247),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_235),
.B(n_238),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_248),
.B1(n_242),
.B2(n_238),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_215),
.B1(n_197),
.B2(n_199),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_142),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_282),
.B(n_138),
.Y(n_301)
);

AND2x4_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_201),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_259),
.B(n_146),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_203),
.B(n_208),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_206),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_149),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_157),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_272),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_252),
.A2(n_265),
.B1(n_271),
.B2(n_281),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_212),
.B1(n_169),
.B2(n_178),
.Y(n_318)
);

NAND2x1p5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_159),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_154),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_151),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_210),
.C(n_207),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_164),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_254),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

BUFx4f_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_263),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

NAND2x1p5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_312),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_308),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_184),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

NAND2x1p5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_263),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_278),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_268),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_327),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_278),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_298),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

NAND2x1p5_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_257),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_294),
.A2(n_191),
.B1(n_176),
.B2(n_184),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_180),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_291),
.A2(n_140),
.B(n_196),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_303),
.A2(n_202),
.B1(n_198),
.B2(n_189),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_306),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_258),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_287),
.B(n_276),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

A2O1A1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_304),
.A2(n_194),
.B(n_184),
.C(n_9),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_343),
.A2(n_295),
.B1(n_301),
.B2(n_300),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

NAND2x1_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_350),
.Y(n_374)
);

AND2x6_ASAP7_75t_SL g375 ( 
.A(n_357),
.B(n_324),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_347),
.A2(n_346),
.B(n_360),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_366),
.B(n_358),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

NAND2x1p5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_328),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_332),
.A2(n_310),
.B(n_319),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_318),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_339),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_323),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_344),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_355),
.A2(n_322),
.B(n_194),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_369),
.B(n_336),
.C(n_337),
.Y(n_390)
);

BUFx2_ASAP7_75t_SL g391 ( 
.A(n_330),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_355),
.A2(n_194),
.B(n_7),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_322),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_354),
.A2(n_352),
.B(n_363),
.Y(n_394)
);

AO21x2_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_322),
.B(n_11),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_362),
.A2(n_78),
.B(n_12),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_79),
.B(n_16),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_365),
.A2(n_340),
.B(n_359),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_373),
.A2(n_338),
.B1(n_345),
.B2(n_330),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_348),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_371),
.A2(n_343),
.B1(n_367),
.B2(n_361),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_390),
.A2(n_353),
.B(n_351),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_378),
.A2(n_397),
.B(n_396),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_343),
.B1(n_385),
.B2(n_370),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_385),
.A2(n_343),
.B1(n_367),
.B2(n_364),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_380),
.A2(n_353),
.B(n_351),
.C(n_8),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_391),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_19),
.B(n_24),
.C(n_26),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_384),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_383),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_387),
.B1(n_376),
.B2(n_388),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

OA211x2_ASAP7_75t_L g417 ( 
.A1(n_374),
.A2(n_34),
.B(n_40),
.C(n_41),
.Y(n_417)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_42),
.B(n_45),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_383),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_419)
);

OR2x2_ASAP7_75t_SL g420 ( 
.A(n_403),
.B(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_399),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_399),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_399),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_387),
.B1(n_392),
.B2(n_393),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_405),
.B(n_392),
.Y(n_429)
);

OAI221xp5_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_382),
.B1(n_375),
.B2(n_398),
.C(n_395),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_398),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_382),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_R g437 ( 
.A(n_435),
.B(n_394),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_395),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_422),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_413),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_433),
.B(n_408),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_389),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_418),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_428),
.A2(n_419),
.B1(n_417),
.B2(n_56),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_417),
.C(n_54),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_434),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_427),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_429),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_440),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_439),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_429),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

AOI211x1_ASAP7_75t_L g460 ( 
.A1(n_447),
.A2(n_420),
.B(n_429),
.C(n_62),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_426),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_452),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_426),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_60),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_65),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_438),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_69),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_456),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_449),
.C(n_451),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_448),
.Y(n_472)
);

OAI21xp33_ASAP7_75t_L g473 ( 
.A1(n_455),
.A2(n_444),
.B(n_437),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_444),
.Y(n_474)
);

AOI322xp5_ASAP7_75t_L g475 ( 
.A1(n_473),
.A2(n_454),
.A3(n_465),
.B1(n_462),
.B2(n_467),
.C1(n_453),
.C2(n_466),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_471),
.A2(n_472),
.B(n_464),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_476),
.A2(n_469),
.B(n_459),
.C(n_470),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_474),
.Y(n_479)
);

AOI21xp33_ASAP7_75t_L g480 ( 
.A1(n_478),
.A2(n_461),
.B(n_463),
.Y(n_480)
);

AOI211xp5_ASAP7_75t_L g481 ( 
.A1(n_479),
.A2(n_461),
.B(n_475),
.C(n_72),
.Y(n_481)
);

NAND4xp25_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_73),
.C(n_76),
.D(n_80),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_480),
.B(n_82),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_95),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_97),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_484),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_486),
.B(n_485),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_99),
.B(n_100),
.Y(n_488)
);

XNOR2x1_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_112),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_117),
.B(n_119),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_120),
.Y(n_491)
);

AOI221x1_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_123),
.B1(n_126),
.B2(n_129),
.C(n_130),
.Y(n_492)
);


endmodule