module fake_jpeg_31240_n_370 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_370);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_370;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_66),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_61),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_8),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_75),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_21),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_42),
.B1(n_20),
.B2(n_36),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_34),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_17),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_45),
.B1(n_59),
.B2(n_65),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_77),
.B(n_102),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_87),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_84),
.A2(n_111),
.B(n_117),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_36),
.B1(n_23),
.B2(n_38),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_107),
.B1(n_112),
.B2(n_118),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_18),
.B1(n_38),
.B2(n_42),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_98),
.B1(n_100),
.B2(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_120),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_44),
.A2(n_23),
.B1(n_36),
.B2(n_18),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_38),
.B1(n_18),
.B2(n_42),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_63),
.A2(n_42),
.B1(n_39),
.B2(n_20),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_58),
.B1(n_70),
.B2(n_55),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_41),
.B1(n_40),
.B2(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_41),
.B1(n_31),
.B2(n_29),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_35),
.B1(n_27),
.B2(n_29),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_31),
.B1(n_28),
.B2(n_22),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_49),
.A2(n_28),
.B(n_1),
.C(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_66),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_51),
.A2(n_56),
.B1(n_68),
.B2(n_64),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_50),
.B(n_0),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_72),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_46),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_10),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_127),
.B(n_143),
.Y(n_192)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_77),
.B1(n_96),
.B2(n_110),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_136),
.Y(n_171)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_108),
.B1(n_93),
.B2(n_114),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_106),
.B1(n_77),
.B2(n_119),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_79),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_151),
.Y(n_172)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_140),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_142),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_9),
.B(n_15),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_57),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_144),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_146),
.Y(n_200)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_72),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_82),
.B(n_0),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_9),
.Y(n_151)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_158),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_157),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_1),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_94),
.B(n_5),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_10),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_10),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_11),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_1),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_77),
.C(n_89),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_166),
.B(n_188),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_169),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_96),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_175),
.A2(n_186),
.B(n_138),
.C(n_133),
.D(n_152),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_110),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_80),
.Y(n_182)
);

BUFx24_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_81),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_119),
.C(n_81),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_81),
.C(n_109),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_163),
.C(n_164),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_109),
.B(n_3),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_3),
.B(n_4),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_2),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_124),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_11),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_125),
.B1(n_129),
.B2(n_137),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_222),
.B1(n_179),
.B2(n_186),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_158),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_209),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_214),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_145),
.B(n_134),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_212),
.A2(n_167),
.B(n_202),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_219),
.B(n_223),
.Y(n_252)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_146),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_176),
.A2(n_125),
.B1(n_137),
.B2(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_229),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_235),
.B(n_179),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_135),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_154),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_153),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_234),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g236 ( 
.A1(n_191),
.A2(n_155),
.B(n_142),
.C(n_15),
.D(n_141),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_182),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_192),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_177),
.B1(n_185),
.B2(n_198),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_217),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_173),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_262),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_196),
.B(n_229),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_175),
.B(n_189),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_223),
.B(n_212),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_207),
.A2(n_169),
.B1(n_168),
.B2(n_167),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_264),
.B1(n_228),
.B2(n_236),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_188),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_207),
.A2(n_222),
.B1(n_206),
.B2(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_168),
.C(n_196),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_219),
.C(n_207),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_266),
.A2(n_273),
.B(n_287),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_237),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_275),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_218),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_269),
.C(n_271),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_219),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_257),
.B1(n_238),
.B2(n_245),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_204),
.C(n_215),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_247),
.C(n_253),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_168),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

BUFx12f_ASAP7_75t_SL g279 ( 
.A(n_259),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_284),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_288),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_286),
.A2(n_251),
.B1(n_258),
.B2(n_249),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_238),
.A2(n_260),
.B(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_242),
.B(n_205),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_297),
.B1(n_300),
.B2(n_295),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_286),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_226),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_257),
.B1(n_261),
.B2(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_261),
.B1(n_263),
.B2(n_250),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.C(n_274),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_255),
.C(n_250),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_317),
.B1(n_318),
.B2(n_306),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_320),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_266),
.B(n_273),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_311),
.A2(n_291),
.B(n_307),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_294),
.B1(n_300),
.B2(n_296),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_278),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_316),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_280),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_269),
.B1(n_268),
.B2(n_276),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_285),
.B1(n_277),
.B2(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_255),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_270),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_323),
.B1(n_298),
.B2(n_217),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_232),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_324),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_326),
.A2(n_318),
.B1(n_312),
.B2(n_298),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_333),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_303),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_324),
.C(n_317),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_294),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_335),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_303),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_337),
.A2(n_309),
.B(n_308),
.Y(n_339)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_216),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_333),
.C(n_335),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_344),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_343),
.A2(n_347),
.B1(n_336),
.B2(n_256),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_323),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_270),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_213),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_329),
.A2(n_256),
.B1(n_177),
.B2(n_234),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_342),
.A2(n_327),
.B(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_351),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_345),
.A2(n_332),
.B1(n_331),
.B2(n_233),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_353),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_224),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g359 ( 
.A1(n_354),
.A2(n_347),
.B(n_184),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_SL g357 ( 
.A(n_355),
.B(n_356),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_338),
.A2(n_199),
.B(n_185),
.Y(n_356)
);

AOI21x1_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_339),
.B(n_345),
.Y(n_358)
);

AOI322xp5_ASAP7_75t_L g363 ( 
.A1(n_358),
.A2(n_348),
.A3(n_352),
.B1(n_350),
.B2(n_340),
.C1(n_341),
.C2(n_174),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_195),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_363),
.A2(n_364),
.B(n_365),
.Y(n_366)
);

OAI221xp5_ASAP7_75t_L g364 ( 
.A1(n_361),
.A2(n_357),
.B1(n_362),
.B2(n_360),
.C(n_174),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_365),
.A2(n_198),
.B(n_194),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_366),
.B(n_194),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_369),
.B(n_128),
.Y(n_370)
);


endmodule